netcdf DISF_NaF {
dimensions:
	NQVALUES = 10 ;
	NTIMES = 2000 ;
	NOCTANS = 8 ;
	OCTANNAME = 8 ;
	NFREQUENCIES = 2000 ;
variables:
	double q(NQVALUES) ;
		q:units = "nm^-1" ;
	double time(NTIMES) ;
		time:units = "ps" ;
	char octan(NOCTANS, OCTANNAME) ;
		octan:units = "unitless" ;
	int qvectors_statistics(NQVALUES, NOCTANS) ;
	double Fqt-Na(NQVALUES, NTIMES) ;
		Fqt-Na:units = "unitless" ;
	double Fqt-total(NQVALUES, NTIMES) ;
		Fqt-total:units = "unitless" ;
	double Fqt-F(NQVALUES, NTIMES) ;
		Fqt-F:units = "unitless" ;
	double frequency(NFREQUENCIES) ;
		frequency:units = "THz" ;
	double angular_frequency(NFREQUENCIES) ;
		angular_frequency:units = "rad ps-1" ;
	double time_resolution(NFREQUENCIES) ;
		time_resolution:units = "unitless" ;
	double frequency_resolution(NFREQUENCIES) ;
		frequency_resolution:units = "unitless" ;
	double Sqw-Na(NQVALUES, NFREQUENCIES) ;
		Sqw-Na:units = "unitless" ;
	double Sqw-total(NQVALUES, NFREQUENCIES) ;
		Sqw-total:units = "unitless" ;
	double Sqw-F(NQVALUES, NFREQUENCIES) ;
		Sqw-F:units = "unitless" ;

// global attributes:
		:title = "DynamicIncoherentStructureFactor_serial" ;
		:jobinfo = "##########################################################################################\n",
			"Job information for DynamicIncoherentStructureFactor_serial analysis.\n",
			"##########################################################################################\n",
			"\n",
			"Job launched on: Tue Jan  8 16:59:52 2013\n",
			"\n",
			"General informations\n",
			"--------------------\n",
			"User: sm37\n",
			"OS: Linux-2.6.32-279.11.1.el6.x86_64\n",
			"Processor: x86_64\n",
			"nMOLDYN version: 3.0.8\n",
			"Estimate run: no\n",
			"\n",
			"Parameters\n",
			"----------\n",
			"subset = all\n",
			"timeinfo = 1:2000:1\n",
			"trajectory = /home/sm37/Projects/NaF-MD/NVT-300K/NPT-1300K/30ps/NaF.nc\n",
			"qvectorsdirection = no\n",
			"pyroserver = monoprocessor\n",
			"qshellvalues = 0.0:100.0:10.0\n",
			"weights = incoherent\n",
			"deuteration = no\n",
			"qshellwidth = 10.0\n",
			"output = /home/sm37/Projects/NaF-MD/NVT-300K/NPT-1300K/30ps/DISF_NaF.nc\n",
			"qvectorsgenerator = 3D isotropic\n",
			"resolution = 10.0\n",
			"qvectorspershell = 50\n",
			"\n",
			"Job status\n",
			"----------\n",
			"\n",
			"Output file written on: Tue Jan  8 17:00:20 2013\n",
			"\n",
			"" ;
data:

 q = 10, 20, 30, 40, 50, 60, 70, 80, 90, 100 ;

 time = 0, 0.0020000000949949026, 0.0040000001899898052, 
    0.0060000002849847078, 0.0080000003799796104, 0.010000000474974513, 
    0.012000000569969416, 0.014000000664964318, 0.016000000759959221, 
    0.018000000854954123, 0.020000000949949026, 0.022000001044943929, 
    0.024000001139938831, 0.026000001234933734, 0.028000001329928637, 
    0.030000001424923539, 0.032000001519918442, 0.034000001614913344, 
    0.036000001709908247, 0.03800000180490315, 0.040000001899898052, 
    0.042000001994892955, 0.044000002089887857, 0.04600000218488276, 
    0.048000002279877663, 0.050000002374872565, 0.052000002469867468, 
    0.05400000256486237, 0.056000002659857273, 0.058000002754852176, 
    0.060000002849847078, 0.062000002944841981, 0.064000003039836884, 
    0.066000003134831786, 0.068000003229826689, 0.070000003324821591, 
    0.072000003419816494, 0.074000003514811397, 0.076000003609806299, 
    0.078000003704801202, 0.080000003799796104, 0.082000003894791007, 
    0.08400000398978591, 0.086000004084780812, 0.088000004179775715, 
    0.090000004274770617, 0.09200000436976552, 0.094000004464760423, 
    0.096000004559755325, 0.098000004654750228, 0.10000000474974513, 
    0.10200000484474003, 0.10400000493973494, 0.10600000503472984, 
    0.10800000512972474, 0.11000000522471964, 0.11200000531971455, 
    0.11400000541470945, 0.11600000550970435, 0.11800000560469925, 
    0.12000000569969416, 0.12200000579468906, 0.12400000588968396, 
    0.12600000598467886, 0.12800000607967377, 0.13000000617466867, 
    0.13200000626966357, 0.13400000636465847, 0.13600000645965338, 
    0.13800000655464828, 0.14000000664964318, 0.14200000674463809, 
    0.14400000683963299, 0.14600000693462789, 0.14800000702962279, 
    0.1500000071246177, 0.1520000072196126, 0.1540000073146075, 
    0.1560000074096024, 0.15800000750459731, 0.16000000759959221, 
    0.16200000769458711, 0.16400000778958201, 0.16600000788457692, 
    0.16800000797957182, 0.17000000807456672, 0.17200000816956162, 
    0.17400000826455653, 0.17600000835955143, 0.17800000845454633, 
    0.18000000854954123, 0.18200000864453614, 0.18400000873953104, 
    0.18600000883452594, 0.18800000892952085, 0.19000000902451575, 
    0.19200000911951065, 0.19400000921450555, 0.19600000930950046, 
    0.19800000940449536, 0.20000000949949026, 0.20200000959448516, 
    0.20400000968948007, 0.20600000978447497, 0.20800000987946987, 
    0.21000000997446477, 0.21200001006945968, 0.21400001016445458, 
    0.21600001025944948, 0.21800001035444438, 0.22000001044943929, 
    0.22200001054443419, 0.22400001063942909, 0.226000010734424, 
    0.2280000108294189, 0.2300000109244138, 0.2320000110194087, 
    0.23400001111440361, 0.23600001120939851, 0.23800001130439341, 
    0.24000001139938831, 0.24200001149438322, 0.24400001158937812, 
    0.24600001168437302, 0.24800001177936792, 0.25000001187436283, 
    0.25200001196935773, 0.25400001206435263, 0.25600001215934753, 
    0.25800001225434244, 0.26000001234933734, 0.26200001244433224, 
    0.26400001253932714, 0.26600001263432205, 0.26800001272931695, 
    0.27000001282431185, 0.27200001291930676, 0.27400001301430166, 
    0.27600001310929656, 0.27800001320429146, 0.28000001329928637, 
    0.28200001339428127, 0.28400001348927617, 0.28600001358427107, 
    0.28800001367926598, 0.29000001377426088, 0.29200001386925578, 
    0.29400001396425068, 0.29600001405924559, 0.29800001415424049, 
    0.30000001424923539, 0.30200001434423029, 0.3040000144392252, 
    0.3060000145342201, 0.308000014629215, 0.3100000147242099, 
    0.31200001481920481, 0.31400001491419971, 0.31600001500919461, 
    0.31800001510418952, 0.32000001519918442, 0.32200001529417932, 
    0.32400001538917422, 0.32600001548416913, 0.32800001557916403, 
    0.33000001567415893, 0.33200001576915383, 0.33400001586414874, 
    0.33600001595914364, 0.33800001605413854, 0.34000001614913344, 
    0.34200001624412835, 0.34400001633912325, 0.34600001643411815, 
    0.34800001652911305, 0.35000001662410796, 0.35200001671910286, 
    0.35400001681409776, 0.35600001690909266, 0.35800001700408757, 
    0.36000001709908247, 0.36200001719407737, 0.36400001728907228, 
    0.36600001738406718, 0.36800001747906208, 0.37000001757405698, 
    0.37200001766905189, 0.37400001776404679, 0.37600001785904169, 
    0.37800001795403659, 0.3800000180490315, 0.3820000181440264, 
    0.3840000182390213, 0.3860000183340162, 0.38800001842901111, 
    0.39000001852400601, 0.39200001861900091, 0.39400001871399581, 
    0.39600001880899072, 0.39800001890398562, 0.40000001899898052, 
    0.40200001909397542, 0.40400001918897033, 0.40600001928396523, 
    0.40800001937896013, 0.41000001947395504, 0.41200001956894994, 
    0.41400001966394484, 0.41600001975893974, 0.41800001985393465, 
    0.42000001994892955, 0.42200002004392445, 0.42400002013891935, 
    0.42600002023391426, 0.42800002032890916, 0.43000002042390406, 
    0.43200002051889896, 0.43400002061389387, 0.43600002070888877, 
    0.43800002080388367, 0.44000002089887857, 0.44200002099387348, 
    0.44400002108886838, 0.44600002118386328, 0.44800002127885818, 
    0.45000002137385309, 0.45200002146884799, 0.45400002156384289, 
    0.4560000216588378, 0.4580000217538327, 0.4600000218488276, 
    0.4620000219438225, 0.46400002203881741, 0.46600002213381231, 
    0.46800002222880721, 0.47000002232380211, 0.47200002241879702, 
    0.47400002251379192, 0.47600002260878682, 0.47800002270378172, 
    0.48000002279877663, 0.48200002289377153, 0.48400002298876643, 
    0.48600002308376133, 0.48800002317875624, 0.49000002327375114, 
    0.49200002336874604, 0.49400002346374094, 0.49600002355873585, 
    0.49800002365373075, 0.50000002374872565, 0.50200002384372056, 
    0.50400002393871546, 0.50600002403371036, 0.50800002412870526, 
    0.51000002422370017, 0.51200002431869507, 0.51400002441368997, 
    0.51600002450868487, 0.51800002460367978, 0.52000002469867468, 
    0.52200002479366958, 0.52400002488866448, 0.52600002498365939, 
    0.52800002507865429, 0.53000002517364919, 0.53200002526864409, 
    0.534000025363639, 0.5360000254586339, 0.5380000255536288, 
    0.5400000256486237, 0.54200002574361861, 0.54400002583861351, 
    0.54600002593360841, 0.54800002602860332, 0.55000002612359822, 
    0.55200002621859312, 0.55400002631358802, 0.55600002640858293, 
    0.55800002650357783, 0.56000002659857273, 0.56200002669356763, 
    0.56400002678856254, 0.56600002688355744, 0.56800002697855234, 
    0.57000002707354724, 0.57200002716854215, 0.57400002726353705, 
    0.57600002735853195, 0.57800002745352685, 0.58000002754852176, 
    0.58200002764351666, 0.58400002773851156, 0.58600002783350646, 
    0.58800002792850137, 0.59000002802349627, 0.59200002811849117, 
    0.59400002821348608, 0.59600002830848098, 0.59800002840347588, 
    0.60000002849847078, 0.60200002859346569, 0.60400002868846059, 
    0.60600002878345549, 0.60800002887845039, 0.6100000289734453, 
    0.6120000290684402, 0.6140000291634351, 0.61600002925843, 
    0.61800002935342491, 0.62000002944841981, 0.62200002954341471, 
    0.62400002963840961, 0.62600002973340452, 0.62800002982839942, 
    0.63000002992339432, 0.63200003001838923, 0.63400003011338413, 
    0.63600003020837903, 0.63800003030337393, 0.64000003039836884, 
    0.64200003049336374, 0.64400003058835864, 0.64600003068335354, 
    0.64800003077834845, 0.65000003087334335, 0.65200003096833825, 
    0.65400003106333315, 0.65600003115832806, 0.65800003125332296, 
    0.66000003134831786, 0.66200003144331276, 0.66400003153830767, 
    0.66600003163330257, 0.66800003172829747, 0.67000003182329237, 
    0.67200003191828728, 0.67400003201328218, 0.67600003210827708, 
    0.67800003220327199, 0.68000003229826689, 0.68200003239326179, 
    0.68400003248825669, 0.6860000325832516, 0.6880000326782465, 
    0.6900000327732414, 0.6920000328682363, 0.69400003296323121, 
    0.69600003305822611, 0.69800003315322101, 0.70000003324821591, 
    0.70200003334321082, 0.70400003343820572, 0.70600003353320062, 
    0.70800003362819552, 0.71000003372319043, 0.71200003381818533, 
    0.71400003391318023, 0.71600003400817513, 0.71800003410317004, 
    0.72000003419816494, 0.72200003429315984, 0.72400003438815475, 
    0.72600003448314965, 0.72800003457814455, 0.73000003467313945, 
    0.73200003476813436, 0.73400003486312926, 0.73600003495812416, 
    0.73800003505311906, 0.74000003514811397, 0.74200003524310887, 
    0.74400003533810377, 0.74600003543309867, 0.74800003552809358, 
    0.75000003562308848, 0.75200003571808338, 0.75400003581307828, 
    0.75600003590807319, 0.75800003600306809, 0.76000003609806299, 
    0.76200003619305789, 0.7640000362880528, 0.7660000363830477, 
    0.7680000364780426, 0.77000003657303751, 0.77200003666803241, 
    0.77400003676302731, 0.77600003685802221, 0.77800003695301712, 
    0.78000003704801202, 0.78200003714300692, 0.78400003723800182, 
    0.78600003733299673, 0.78800003742799163, 0.79000003752298653, 
    0.79200003761798143, 0.79400003771297634, 0.79600003780797124, 
    0.79800003790296614, 0.80000003799796104, 0.80200003809295595, 
    0.80400003818795085, 0.80600003828294575, 0.80800003837794065, 
    0.81000003847293556, 0.81200003856793046, 0.81400003866292536, 
    0.81600003875792027, 0.81800003885291517, 0.82000003894791007, 
    0.82200003904290497, 0.82400003913789988, 0.82600003923289478, 
    0.82800003932788968, 0.83000003942288458, 0.83200003951787949, 
    0.83400003961287439, 0.83600003970786929, 0.83800003980286419, 
    0.8400000398978591, 0.842000039992854, 0.8440000400878489, 
    0.8460000401828438, 0.84800004027783871, 0.85000004037283361, 
    0.85200004046782851, 0.85400004056282341, 0.85600004065781832, 
    0.85800004075281322, 0.86000004084780812, 0.86200004094280303, 
    0.86400004103779793, 0.86600004113279283, 0.86800004122778773, 
    0.87000004132278264, 0.87200004141777754, 0.87400004151277244, 
    0.87600004160776734, 0.87800004170276225, 0.88000004179775715, 
    0.88200004189275205, 0.88400004198774695, 0.88600004208274186, 
    0.88800004217773676, 0.89000004227273166, 0.89200004236772656, 
    0.89400004246272147, 0.89600004255771637, 0.89800004265271127, 
    0.90000004274770617, 0.90200004284270108, 0.90400004293769598, 
    0.90600004303269088, 0.90800004312768579, 0.91000004322268069, 
    0.91200004331767559, 0.91400004341267049, 0.9160000435076654, 
    0.9180000436026603, 0.9200000436976552, 0.9220000437926501, 
    0.92400004388764501, 0.92600004398263991, 0.92800004407763481, 
    0.93000004417262971, 0.93200004426762462, 0.93400004436261952, 
    0.93600004445761442, 0.93800004455260932, 0.94000004464760423, 
    0.94200004474259913, 0.94400004483759403, 0.94600004493258893, 
    0.94800004502758384, 0.95000004512257874, 0.95200004521757364, 
    0.95400004531256855, 0.95600004540756345, 0.95800004550255835, 
    0.96000004559755325, 0.96200004569254816, 0.96400004578754306, 
    0.96600004588253796, 0.96800004597753286, 0.97000004607252777, 
    0.97200004616752267, 0.97400004626251757, 0.97600004635751247, 
    0.97800004645250738, 0.98000004654750228, 0.98200004664249718, 
    0.98400004673749208, 0.98600004683248699, 0.98800004692748189, 
    0.99000004702247679, 0.99200004711747169, 0.9940000472124666, 
    0.9960000473074615, 0.9980000474024564, 1.0000000474974513, 
    1.0020000475924462, 1.0040000476874411, 1.006000047782436, 
    1.0080000478774309, 1.0100000479724258, 1.0120000480674207, 
    1.0140000481624156, 1.0160000482574105, 1.0180000483524054, 
    1.0200000484474003, 1.0220000485423952, 1.0240000486373901, 
    1.026000048732385, 1.0280000488273799, 1.0300000489223748, 
    1.0320000490173697, 1.0340000491123646, 1.0360000492073596, 
    1.0380000493023545, 1.0400000493973494, 1.0420000494923443, 
    1.0440000495873392, 1.0460000496823341, 1.048000049777329, 
    1.0500000498723239, 1.0520000499673188, 1.0540000500623137, 
    1.0560000501573086, 1.0580000502523035, 1.0600000503472984, 
    1.0620000504422933, 1.0640000505372882, 1.0660000506322831, 
    1.068000050727278, 1.0700000508222729, 1.0720000509172678, 
    1.0740000510122627, 1.0760000511072576, 1.0780000512022525, 
    1.0800000512972474, 1.0820000513922423, 1.0840000514872372, 
    1.0860000515822321, 1.088000051677227, 1.0900000517722219, 
    1.0920000518672168, 1.0940000519622117, 1.0960000520572066, 
    1.0980000521522015, 1.1000000522471964, 1.1020000523421913, 
    1.1040000524371862, 1.1060000525321811, 1.108000052627176, 
    1.1100000527221709, 1.1120000528171659, 1.1140000529121608, 
    1.1160000530071557, 1.1180000531021506, 1.1200000531971455, 
    1.1220000532921404, 1.1240000533871353, 1.1260000534821302, 
    1.1280000535771251, 1.13000005367212, 1.1320000537671149, 
    1.1340000538621098, 1.1360000539571047, 1.1380000540520996, 
    1.1400000541470945, 1.1420000542420894, 1.1440000543370843, 
    1.1460000544320792, 1.1480000545270741, 1.150000054622069, 
    1.1520000547170639, 1.1540000548120588, 1.1560000549070537, 
    1.1580000550020486, 1.1600000550970435, 1.1620000551920384, 
    1.1640000552870333, 1.1660000553820282, 1.1680000554770231, 
    1.170000055572018, 1.1720000556670129, 1.1740000557620078, 
    1.1760000558570027, 1.1780000559519976, 1.1800000560469925, 
    1.1820000561419874, 1.1840000562369823, 1.1860000563319772, 
    1.1880000564269722, 1.1900000565219671, 1.192000056616962, 
    1.1940000567119569, 1.1960000568069518, 1.1980000569019467, 
    1.2000000569969416, 1.2020000570919365, 1.2040000571869314, 
    1.2060000572819263, 1.2080000573769212, 1.2100000574719161, 
    1.212000057566911, 1.2140000576619059, 1.2160000577569008, 
    1.2180000578518957, 1.2200000579468906, 1.2220000580418855, 
    1.2240000581368804, 1.2260000582318753, 1.2280000583268702, 
    1.2300000584218651, 1.23200005851686, 1.2340000586118549, 
    1.2360000587068498, 1.2380000588018447, 1.2400000588968396, 
    1.2420000589918345, 1.2440000590868294, 1.2460000591818243, 
    1.2480000592768192, 1.2500000593718141, 1.252000059466809, 
    1.2540000595618039, 1.2560000596567988, 1.2580000597517937, 
    1.2600000598467886, 1.2620000599417835, 1.2640000600367785, 
    1.2660000601317734, 1.2680000602267683, 1.2700000603217632, 
    1.2720000604167581, 1.274000060511753, 1.2760000606067479, 
    1.2780000607017428, 1.2800000607967377, 1.2820000608917326, 
    1.2840000609867275, 1.2860000610817224, 1.2880000611767173, 
    1.2900000612717122, 1.2920000613667071, 1.294000061461702, 
    1.2960000615566969, 1.2980000616516918, 1.3000000617466867, 
    1.3020000618416816, 1.3040000619366765, 1.3060000620316714, 
    1.3080000621266663, 1.3100000622216612, 1.3120000623166561, 
    1.314000062411651, 1.3160000625066459, 1.3180000626016408, 
    1.3200000626966357, 1.3220000627916306, 1.3240000628866255, 
    1.3260000629816204, 1.3280000630766153, 1.3300000631716102, 
    1.3320000632666051, 1.3340000633616, 1.3360000634565949, 
    1.3380000635515898, 1.3400000636465847, 1.3420000637415797, 
    1.3440000638365746, 1.3460000639315695, 1.3480000640265644, 
    1.3500000641215593, 1.3520000642165542, 1.3540000643115491, 
    1.356000064406544, 1.3580000645015389, 1.3600000645965338, 
    1.3620000646915287, 1.3640000647865236, 1.3660000648815185, 
    1.3680000649765134, 1.3700000650715083, 1.3720000651665032, 
    1.3740000652614981, 1.376000065356493, 1.3780000654514879, 
    1.3800000655464828, 1.3820000656414777, 1.3840000657364726, 
    1.3860000658314675, 1.3880000659264624, 1.3900000660214573, 
    1.3920000661164522, 1.3940000662114471, 1.396000066306442, 
    1.3980000664014369, 1.4000000664964318, 1.4020000665914267, 
    1.4040000666864216, 1.4060000667814165, 1.4080000668764114, 
    1.4100000669714063, 1.4120000670664012, 1.4140000671613961, 
    1.416000067256391, 1.418000067351386, 1.4200000674463809, 
    1.4220000675413758, 1.4240000676363707, 1.4260000677313656, 
    1.4280000678263605, 1.4300000679213554, 1.4320000680163503, 
    1.4340000681113452, 1.4360000682063401, 1.438000068301335, 
    1.4400000683963299, 1.4420000684913248, 1.4440000685863197, 
    1.4460000686813146, 1.4480000687763095, 1.4500000688713044, 
    1.4520000689662993, 1.4540000690612942, 1.4560000691562891, 
    1.458000069251284, 1.4600000693462789, 1.4620000694412738, 
    1.4640000695362687, 1.4660000696312636, 1.4680000697262585, 
    1.4700000698212534, 1.4720000699162483, 1.4740000700112432, 
    1.4760000701062381, 1.478000070201233, 1.4800000702962279, 
    1.4820000703912228, 1.4840000704862177, 1.4860000705812126, 
    1.4880000706762075, 1.4900000707712024, 1.4920000708661973, 
    1.4940000709611923, 1.4960000710561872, 1.4980000711511821, 
    1.500000071246177, 1.5020000713411719, 1.5040000714361668, 
    1.5060000715311617, 1.5080000716261566, 1.5100000717211515, 
    1.5120000718161464, 1.5140000719111413, 1.5160000720061362, 
    1.5180000721011311, 1.520000072196126, 1.5220000722911209, 
    1.5240000723861158, 1.5260000724811107, 1.5280000725761056, 
    1.5300000726711005, 1.5320000727660954, 1.5340000728610903, 
    1.5360000729560852, 1.5380000730510801, 1.540000073146075, 
    1.5420000732410699, 1.5440000733360648, 1.5460000734310597, 
    1.5480000735260546, 1.5500000736210495, 1.5520000737160444, 
    1.5540000738110393, 1.5560000739060342, 1.5580000740010291, 
    1.560000074096024, 1.5620000741910189, 1.5640000742860138, 
    1.5660000743810087, 1.5680000744760036, 1.5700000745709985, 
    1.5720000746659935, 1.5740000747609884, 1.5760000748559833, 
    1.5780000749509782, 1.5800000750459731, 1.582000075140968, 
    1.5840000752359629, 1.5860000753309578, 1.5880000754259527, 
    1.5900000755209476, 1.5920000756159425, 1.5940000757109374, 
    1.5960000758059323, 1.5980000759009272, 1.6000000759959221, 
    1.602000076090917, 1.6040000761859119, 1.6060000762809068, 
    1.6080000763759017, 1.6100000764708966, 1.6120000765658915, 
    1.6140000766608864, 1.6160000767558813, 1.6180000768508762, 
    1.6200000769458711, 1.622000077040866, 1.6240000771358609, 
    1.6260000772308558, 1.6280000773258507, 1.6300000774208456, 
    1.6320000775158405, 1.6340000776108354, 1.6360000777058303, 
    1.6380000778008252, 1.6400000778958201, 1.642000077990815, 
    1.6440000780858099, 1.6460000781808048, 1.6480000782757998, 
    1.6500000783707947, 1.6520000784657896, 1.6540000785607845, 
    1.6560000786557794, 1.6580000787507743, 1.6600000788457692, 
    1.6620000789407641, 1.664000079035759, 1.6660000791307539, 
    1.6680000792257488, 1.6700000793207437, 1.6720000794157386, 
    1.6740000795107335, 1.6760000796057284, 1.6780000797007233, 
    1.6800000797957182, 1.6820000798907131, 1.684000079985708, 
    1.6860000800807029, 1.6880000801756978, 1.6900000802706927, 
    1.6920000803656876, 1.6940000804606825, 1.6960000805556774, 
    1.6980000806506723, 1.7000000807456672, 1.7020000808406621, 
    1.704000080935657, 1.7060000810306519, 1.7080000811256468, 
    1.7100000812206417, 1.7120000813156366, 1.7140000814106315, 
    1.7160000815056264, 1.7180000816006213, 1.7200000816956162, 
    1.7220000817906111, 1.7240000818856061, 1.726000081980601, 
    1.7280000820755959, 1.7300000821705908, 1.7320000822655857, 
    1.7340000823605806, 1.7360000824555755, 1.7380000825505704, 
    1.7400000826455653, 1.7420000827405602, 1.7440000828355551, 
    1.74600008293055, 1.7480000830255449, 1.7500000831205398, 
    1.7520000832155347, 1.7540000833105296, 1.7560000834055245, 
    1.7580000835005194, 1.7600000835955143, 1.7620000836905092, 
    1.7640000837855041, 1.766000083880499, 1.7680000839754939, 
    1.7700000840704888, 1.7720000841654837, 1.7740000842604786, 
    1.7760000843554735, 1.7780000844504684, 1.7800000845454633, 
    1.7820000846404582, 1.7840000847354531, 1.786000084830448, 
    1.7880000849254429, 1.7900000850204378, 1.7920000851154327, 
    1.7940000852104276, 1.7960000853054225, 1.7980000854004174, 
    1.8000000854954123, 1.8020000855904073, 1.8040000856854022, 
    1.8060000857803971, 1.808000085875392, 1.8100000859703869, 
    1.8120000860653818, 1.8140000861603767, 1.8160000862553716, 
    1.8180000863503665, 1.8200000864453614, 1.8220000865403563, 
    1.8240000866353512, 1.8260000867303461, 1.828000086825341, 
    1.8300000869203359, 1.8320000870153308, 1.8340000871103257, 
    1.8360000872053206, 1.8380000873003155, 1.8400000873953104, 
    1.8420000874903053, 1.8440000875853002, 1.8460000876802951, 
    1.84800008777529, 1.8500000878702849, 1.8520000879652798, 
    1.8540000880602747, 1.8560000881552696, 1.8580000882502645, 
    1.8600000883452594, 1.8620000884402543, 1.8640000885352492, 
    1.8660000886302441, 1.868000088725239, 1.8700000888202339, 
    1.8720000889152288, 1.8740000890102237, 1.8760000891052186, 
    1.8780000892002136, 1.8800000892952085, 1.8820000893902034, 
    1.8840000894851983, 1.8860000895801932, 1.8880000896751881, 
    1.890000089770183, 1.8920000898651779, 1.8940000899601728, 
    1.8960000900551677, 1.8980000901501626, 1.9000000902451575, 
    1.9020000903401524, 1.9040000904351473, 1.9060000905301422, 
    1.9080000906251371, 1.910000090720132, 1.9120000908151269, 
    1.9140000909101218, 1.9160000910051167, 1.9180000911001116, 
    1.9200000911951065, 1.9220000912901014, 1.9240000913850963, 
    1.9260000914800912, 1.9280000915750861, 1.930000091670081, 
    1.9320000917650759, 1.9340000918600708, 1.9360000919550657, 
    1.9380000920500606, 1.9400000921450555, 1.9420000922400504, 
    1.9440000923350453, 1.9460000924300402, 1.9480000925250351, 
    1.95000009262003, 1.9520000927150249, 1.9540000928100199, 
    1.9560000929050148, 1.9580000930000097, 1.9600000930950046, 
    1.9620000931899995, 1.9640000932849944, 1.9660000933799893, 
    1.9680000934749842, 1.9700000935699791, 1.972000093664974, 
    1.9740000937599689, 1.9760000938549638, 1.9780000939499587, 
    1.9800000940449536, 1.9820000941399485, 1.9840000942349434, 
    1.9860000943299383, 1.9880000944249332, 1.9900000945199281, 
    1.992000094614923, 1.9940000947099179, 1.9960000948049128, 
    1.9980000948999077, 2.0000000949949026, 2.0020000950898975, 
    2.0040000951848924, 2.0060000952798873, 2.0080000953748822, 
    2.0100000954698771, 2.012000095564872, 2.0140000956598669, 
    2.0160000957548618, 2.0180000958498567, 2.0200000959448516, 
    2.0220000960398465, 2.0240000961348414, 2.0260000962298363, 
    2.0280000963248312, 2.0300000964198261, 2.0320000965148211, 
    2.034000096609816, 2.0360000967048109, 2.0380000967998058, 
    2.0400000968948007, 2.0420000969897956, 2.0440000970847905, 
    2.0460000971797854, 2.0480000972747803, 2.0500000973697752, 
    2.0520000974647701, 2.054000097559765, 2.0560000976547599, 
    2.0580000977497548, 2.0600000978447497, 2.0620000979397446, 
    2.0640000980347395, 2.0660000981297344, 2.0680000982247293, 
    2.0700000983197242, 2.0720000984147191, 2.074000098509714, 
    2.0760000986047089, 2.0780000986997038, 2.0800000987946987, 
    2.0820000988896936, 2.0840000989846885, 2.0860000990796834, 
    2.0880000991746783, 2.0900000992696732, 2.0920000993646681, 
    2.094000099459663, 2.0960000995546579, 2.0980000996496528, 
    2.1000000997446477, 2.1020000998396426, 2.1040000999346375, 
    2.1060001000296324, 2.1080001001246274, 2.1100001002196223, 
    2.1120001003146172, 2.1140001004096121, 2.116000100504607, 
    2.1180001005996019, 2.1200001006945968, 2.1220001007895917, 
    2.1240001008845866, 2.1260001009795815, 2.1280001010745764, 
    2.1300001011695713, 2.1320001012645662, 2.1340001013595611, 
    2.136000101454556, 2.1380001015495509, 2.1400001016445458, 
    2.1420001017395407, 2.1440001018345356, 2.1460001019295305, 
    2.1480001020245254, 2.1500001021195203, 2.1520001022145152, 
    2.1540001023095101, 2.156000102404505, 2.1580001024994999, 
    2.1600001025944948, 2.1620001026894897, 2.1640001027844846, 
    2.1660001028794795, 2.1680001029744744, 2.1700001030694693, 
    2.1720001031644642, 2.1740001032594591, 2.176000103354454, 
    2.1780001034494489, 2.1800001035444438, 2.1820001036394387, 
    2.1840001037344337, 2.1860001038294286, 2.1880001039244235, 
    2.1900001040194184, 2.1920001041144133, 2.1940001042094082, 
    2.1960001043044031, 2.198000104399398, 2.2000001044943929, 
    2.2020001045893878, 2.2040001046843827, 2.2060001047793776, 
    2.2080001048743725, 2.2100001049693674, 2.2120001050643623, 
    2.2140001051593572, 2.2160001052543521, 2.218000105349347, 
    2.2200001054443419, 2.2220001055393368, 2.2240001056343317, 
    2.2260001057293266, 2.2280001058243215, 2.2300001059193164, 
    2.2320001060143113, 2.2340001061093062, 2.2360001062043011, 
    2.238000106299296, 2.2400001063942909, 2.2420001064892858, 
    2.2440001065842807, 2.2460001066792756, 2.2480001067742705, 
    2.2500001068692654, 2.2520001069642603, 2.2540001070592552, 
    2.2560001071542501, 2.258000107249245, 2.26000010734424, 
    2.2620001074392349, 2.2640001075342298, 2.2660001076292247, 
    2.2680001077242196, 2.2700001078192145, 2.2720001079142094, 
    2.2740001080092043, 2.2760001081041992, 2.2780001081991941, 
    2.280000108294189, 2.2820001083891839, 2.2840001084841788, 
    2.2860001085791737, 2.2880001086741686, 2.2900001087691635, 
    2.2920001088641584, 2.2940001089591533, 2.2960001090541482, 
    2.2980001091491431, 2.300000109244138, 2.3020001093391329, 
    2.3040001094341278, 2.3060001095291227, 2.3080001096241176, 
    2.3100001097191125, 2.3120001098141074, 2.3140001099091023, 
    2.3160001100040972, 2.3180001100990921, 2.320000110194087, 
    2.3220001102890819, 2.3240001103840768, 2.3260001104790717, 
    2.3280001105740666, 2.3300001106690615, 2.3320001107640564, 
    2.3340001108590513, 2.3360001109540462, 2.3380001110490412, 
    2.3400001111440361, 2.342000111239031, 2.3440001113340259, 
    2.3460001114290208, 2.3480001115240157, 2.3500001116190106, 
    2.3520001117140055, 2.3540001118090004, 2.3560001119039953, 
    2.3580001119989902, 2.3600001120939851, 2.36200011218898, 
    2.3640001122839749, 2.3660001123789698, 2.3680001124739647, 
    2.3700001125689596, 2.3720001126639545, 2.3740001127589494, 
    2.3760001128539443, 2.3780001129489392, 2.3800001130439341, 
    2.382000113138929, 2.3840001132339239, 2.3860001133289188, 
    2.3880001134239137, 2.3900001135189086, 2.3920001136139035, 
    2.3940001137088984, 2.3960001138038933, 2.3980001138988882, 
    2.4000001139938831, 2.402000114088878, 2.4040001141838729, 
    2.4060001142788678, 2.4080001143738627, 2.4100001144688576, 
    2.4120001145638525, 2.4140001146588475, 2.4160001147538424, 
    2.4180001148488373, 2.4200001149438322, 2.4220001150388271, 
    2.424000115133822, 2.4260001152288169, 2.4280001153238118, 
    2.4300001154188067, 2.4320001155138016, 2.4340001156087965, 
    2.4360001157037914, 2.4380001157987863, 2.4400001158937812, 
    2.4420001159887761, 2.444000116083771, 2.4460001161787659, 
    2.4480001162737608, 2.4500001163687557, 2.4520001164637506, 
    2.4540001165587455, 2.4560001166537404, 2.4580001167487353, 
    2.4600001168437302, 2.4620001169387251, 2.46400011703372, 
    2.4660001171287149, 2.4680001172237098, 2.4700001173187047, 
    2.4720001174136996, 2.4740001175086945, 2.4760001176036894, 
    2.4780001176986843, 2.4800001177936792, 2.4820001178886741, 
    2.484000117983669, 2.4860001180786639, 2.4880001181736588, 
    2.4900001182686538, 2.4920001183636487, 2.4940001184586436, 
    2.4960001185536385, 2.4980001186486334, 2.5000001187436283, 
    2.5020001188386232, 2.5040001189336181, 2.506000119028613, 
    2.5080001191236079, 2.5100001192186028, 2.5120001193135977, 
    2.5140001194085926, 2.5160001195035875, 2.5180001195985824, 
    2.5200001196935773, 2.5220001197885722, 2.5240001198835671, 
    2.526000119978562, 2.5280001200735569, 2.5300001201685518, 
    2.5320001202635467, 2.5340001203585416, 2.5360001204535365, 
    2.5380001205485314, 2.5400001206435263, 2.5420001207385212, 
    2.5440001208335161, 2.546000120928511, 2.5480001210235059, 
    2.5500001211185008, 2.5520001212134957, 2.5540001213084906, 
    2.5560001214034855, 2.5580001214984804, 2.5600001215934753, 
    2.5620001216884702, 2.5640001217834651, 2.56600012187846, 
    2.568000121973455, 2.5700001220684499, 2.5720001221634448, 
    2.5740001222584397, 2.5760001223534346, 2.5780001224484295, 
    2.5800001225434244, 2.5820001226384193, 2.5840001227334142, 
    2.5860001228284091, 2.588000122923404, 2.5900001230183989, 
    2.5920001231133938, 2.5940001232083887, 2.5960001233033836, 
    2.5980001233983785, 2.6000001234933734, 2.6020001235883683, 
    2.6040001236833632, 2.6060001237783581, 2.608000123873353, 
    2.6100001239683479, 2.6120001240633428, 2.6140001241583377, 
    2.6160001242533326, 2.6180001243483275, 2.6200001244433224, 
    2.6220001245383173, 2.6240001246333122, 2.6260001247283071, 
    2.628000124823302, 2.6300001249182969, 2.6320001250132918, 
    2.6340001251082867, 2.6360001252032816, 2.6380001252982765, 
    2.6400001253932714, 2.6420001254882663, 2.6440001255832613, 
    2.6460001256782562, 2.6480001257732511, 2.650000125868246, 
    2.6520001259632409, 2.6540001260582358, 2.6560001261532307, 
    2.6580001262482256, 2.6600001263432205, 2.6620001264382154, 
    2.6640001265332103, 2.6660001266282052, 2.6680001267232001, 
    2.670000126818195, 2.6720001269131899, 2.6740001270081848, 
    2.6760001271031797, 2.6780001271981746, 2.6800001272931695, 
    2.6820001273881644, 2.6840001274831593, 2.6860001275781542, 
    2.6880001276731491, 2.690000127768144, 2.6920001278631389, 
    2.6940001279581338, 2.6960001280531287, 2.6980001281481236, 
    2.7000001282431185, 2.7020001283381134, 2.7040001284331083, 
    2.7060001285281032, 2.7080001286230981, 2.710000128718093, 
    2.7120001288130879, 2.7140001289080828, 2.7160001290030777, 
    2.7180001290980726, 2.7200001291930676, 2.7220001292880625, 
    2.7240001293830574, 2.7260001294780523, 2.7280001295730472, 
    2.7300001296680421, 2.732000129763037, 2.7340001298580319, 
    2.7360001299530268, 2.7380001300480217, 2.7400001301430166, 
    2.7420001302380115, 2.7440001303330064, 2.7460001304280013, 
    2.7480001305229962, 2.7500001306179911, 2.752000130712986, 
    2.7540001308079809, 2.7560001309029758, 2.7580001309979707, 
    2.7600001310929656, 2.7620001311879605, 2.7640001312829554, 
    2.7660001313779503, 2.7680001314729452, 2.7700001315679401, 
    2.772000131662935, 2.7740001317579299, 2.7760001318529248, 
    2.7780001319479197, 2.7800001320429146, 2.7820001321379095, 
    2.7840001322329044, 2.7860001323278993, 2.7880001324228942, 
    2.7900001325178891, 2.792000132612884, 2.7940001327078789, 
    2.7960001328028738, 2.7980001328978688, 2.8000001329928637, 
    2.8020001330878586, 2.8040001331828535, 2.8060001332778484, 
    2.8080001333728433, 2.8100001334678382, 2.8120001335628331, 
    2.814000133657828, 2.8160001337528229, 2.8180001338478178, 
    2.8200001339428127, 2.8220001340378076, 2.8240001341328025, 
    2.8260001342277974, 2.8280001343227923, 2.8300001344177872, 
    2.8320001345127821, 2.834000134607777, 2.8360001347027719, 
    2.8380001347977668, 2.8400001348927617, 2.8420001349877566, 
    2.8440001350827515, 2.8460001351777464, 2.8480001352727413, 
    2.8500001353677362, 2.8520001354627311, 2.854000135557726, 
    2.8560001356527209, 2.8580001357477158, 2.8600001358427107, 
    2.8620001359377056, 2.8640001360327005, 2.8660001361276954, 
    2.8680001362226903, 2.8700001363176852, 2.8720001364126801, 
    2.8740001365076751, 2.87600013660267, 2.8780001366976649, 
    2.8800001367926598, 2.8820001368876547, 2.8840001369826496, 
    2.8860001370776445, 2.8880001371726394, 2.8900001372676343, 
    2.8920001373626292, 2.8940001374576241, 2.896000137552619, 
    2.8980001376476139, 2.9000001377426088, 2.9020001378376037, 
    2.9040001379325986, 2.9060001380275935, 2.9080001381225884, 
    2.9100001382175833, 2.9120001383125782, 2.9140001384075731, 
    2.916000138502568, 2.9180001385975629, 2.9200001386925578, 
    2.9220001387875527, 2.9240001388825476, 2.9260001389775425, 
    2.9280001390725374, 2.9300001391675323, 2.9320001392625272, 
    2.9340001393575221, 2.936000139452517, 2.9380001395475119, 
    2.9400001396425068, 2.9420001397375017, 2.9440001398324966, 
    2.9460001399274915, 2.9480001400224864, 2.9500001401174814, 
    2.9520001402124763, 2.9540001403074712, 2.9560001404024661, 
    2.958000140497461, 2.9600001405924559, 2.9620001406874508, 
    2.9640001407824457, 2.9660001408774406, 2.9680001409724355, 
    2.9700001410674304, 2.9720001411624253, 2.9740001412574202, 
    2.9760001413524151, 2.97800014144741, 2.9800001415424049, 
    2.9820001416373998, 2.9840001417323947, 2.9860001418273896, 
    2.9880001419223845, 2.9900001420173794, 2.9920001421123743, 
    2.9940001422073692, 2.9960001423023641, 2.998000142397359, 
    3.0000001424923539, 3.0020001425873488, 3.0040001426823437, 
    3.0060001427773386, 3.0080001428723335, 3.0100001429673284, 
    3.0120001430623233, 3.0140001431573182, 3.0160001432523131, 
    3.018000143347308, 3.0200001434423029, 3.0220001435372978, 
    3.0240001436322927, 3.0260001437272877, 3.0280001438222826, 
    3.0300001439172775, 3.0320001440122724, 3.0340001441072673, 
    3.0360001442022622, 3.0380001442972571, 3.040000144392252, 
    3.0420001444872469, 3.0440001445822418, 3.0460001446772367, 
    3.0480001447722316, 3.0500001448672265, 3.0520001449622214, 
    3.0540001450572163, 3.0560001451522112, 3.0580001452472061, 
    3.060000145342201, 3.0620001454371959, 3.0640001455321908, 
    3.0660001456271857, 3.0680001457221806, 3.0700001458171755, 
    3.0720001459121704, 3.0740001460071653, 3.0760001461021602, 
    3.0780001461971551, 3.08000014629215, 3.0820001463871449, 
    3.0840001464821398, 3.0860001465771347, 3.0880001466721296, 
    3.0900001467671245, 3.0920001468621194, 3.0940001469571143, 
    3.0960001470521092, 3.0980001471471041, 3.100000147242099, 
    3.1020001473370939, 3.1040001474320889, 3.1060001475270838, 
    3.1080001476220787, 3.1100001477170736, 3.1120001478120685, 
    3.1140001479070634, 3.1160001480020583, 3.1180001480970532, 
    3.1200001481920481, 3.122000148287043, 3.1240001483820379, 
    3.1260001484770328, 3.1280001485720277, 3.1300001486670226, 
    3.1320001487620175, 3.1340001488570124, 3.1360001489520073, 
    3.1380001490470022, 3.1400001491419971, 3.142000149236992, 
    3.1440001493319869, 3.1460001494269818, 3.1480001495219767, 
    3.1500001496169716, 3.1520001497119665, 3.1540001498069614, 
    3.1560001499019563, 3.1580001499969512, 3.1600001500919461, 
    3.162000150186941, 3.1640001502819359, 3.1660001503769308, 
    3.1680001504719257, 3.1700001505669206, 3.1720001506619155, 
    3.1740001507569104, 3.1760001508519053, 3.1780001509469002, 
    3.1800001510418952, 3.1820001511368901, 3.184000151231885, 
    3.1860001513268799, 3.1880001514218748, 3.1900001515168697, 
    3.1920001516118646, 3.1940001517068595, 3.1960001518018544, 
    3.1980001518968493, 3.2000001519918442, 3.2020001520868391, 
    3.204000152181834, 3.2060001522768289, 3.2080001523718238, 
    3.2100001524668187, 3.2120001525618136, 3.2140001526568085, 
    3.2160001527518034, 3.2180001528467983, 3.2200001529417932, 
    3.2220001530367881, 3.224000153131783, 3.2260001532267779, 
    3.2280001533217728, 3.2300001534167677, 3.2320001535117626, 
    3.2340001536067575, 3.2360001537017524, 3.2380001537967473, 
    3.2400001538917422, 3.2420001539867371, 3.244000154081732, 
    3.2460001541767269, 3.2480001542717218, 3.2500001543667167, 
    3.2520001544617116, 3.2540001545567065, 3.2560001546517015, 
    3.2580001547466964, 3.2600001548416913, 3.2620001549366862, 
    3.2640001550316811, 3.266000155126676, 3.2680001552216709, 
    3.2700001553166658, 3.2720001554116607, 3.2740001555066556, 
    3.2760001556016505, 3.2780001556966454, 3.2800001557916403, 
    3.2820001558866352, 3.2840001559816301, 3.286000156076625, 
    3.2880001561716199, 3.2900001562666148, 3.2920001563616097, 
    3.2940001564566046, 3.2960001565515995, 3.2980001566465944, 
    3.3000001567415893, 3.3020001568365842, 3.3040001569315791, 
    3.306000157026574, 3.3080001571215689, 3.3100001572165638, 
    3.3120001573115587, 3.3140001574065536, 3.3160001575015485, 
    3.3180001575965434, 3.3200001576915383, 3.3220001577865332, 
    3.3240001578815281, 3.326000157976523, 3.3280001580715179, 
    3.3300001581665128, 3.3320001582615077, 3.3340001583565027, 
    3.3360001584514976, 3.3380001585464925, 3.3400001586414874, 
    3.3420001587364823, 3.3440001588314772, 3.3460001589264721, 
    3.348000159021467, 3.3500001591164619, 3.3520001592114568, 
    3.3540001593064517, 3.3560001594014466, 3.3580001594964415, 
    3.3600001595914364, 3.3620001596864313, 3.3640001597814262, 
    3.3660001598764211, 3.368000159971416, 3.3700001600664109, 
    3.3720001601614058, 3.3740001602564007, 3.3760001603513956, 
    3.3780001604463905, 3.3800001605413854, 3.3820001606363803, 
    3.3840001607313752, 3.3860001608263701, 3.388000160921365, 
    3.3900001610163599, 3.3920001611113548, 3.3940001612063497, 
    3.3960001613013446, 3.3980001613963395, 3.4000001614913344, 
    3.4020001615863293, 3.4040001616813242, 3.4060001617763191, 
    3.408000161871314, 3.410000161966309, 3.4120001620613039, 
    3.4140001621562988, 3.4160001622512937, 3.4180001623462886, 
    3.4200001624412835, 3.4220001625362784, 3.4240001626312733, 
    3.4260001627262682, 3.4280001628212631, 3.430000162916258, 
    3.4320001630112529, 3.4340001631062478, 3.4360001632012427, 
    3.4380001632962376, 3.4400001633912325, 3.4420001634862274, 
    3.4440001635812223, 3.4460001636762172, 3.4480001637712121, 
    3.450000163866207, 3.4520001639612019, 3.4540001640561968, 
    3.4560001641511917, 3.4580001642461866, 3.4600001643411815, 
    3.4620001644361764, 3.4640001645311713, 3.4660001646261662, 
    3.4680001647211611, 3.470000164816156, 3.4720001649111509, 
    3.4740001650061458, 3.4760001651011407, 3.4780001651961356, 
    3.4800001652911305, 3.4820001653861254, 3.4840001654811203, 
    3.4860001655761153, 3.4880001656711102, 3.4900001657661051, 
    3.4920001658611, 3.4940001659560949, 3.4960001660510898, 
    3.4980001661460847, 3.5000001662410796, 3.5020001663360745, 
    3.5040001664310694, 3.5060001665260643, 3.5080001666210592, 
    3.5100001667160541, 3.512000166811049, 3.5140001669060439, 
    3.5160001670010388, 3.5180001670960337, 3.5200001671910286, 
    3.5220001672860235, 3.5240001673810184, 3.5260001674760133, 
    3.5280001675710082, 3.5300001676660031, 3.532000167760998, 
    3.5340001678559929, 3.5360001679509878, 3.5380001680459827, 
    3.5400001681409776, 3.5420001682359725, 3.5440001683309674, 
    3.5460001684259623, 3.5480001685209572, 3.5500001686159521, 
    3.552000168710947, 3.5540001688059419, 3.5560001689009368, 
    3.5580001689959317, 3.5600001690909266, 3.5620001691859215, 
    3.5640001692809165, 3.5660001693759114, 3.5680001694709063, 
    3.5700001695659012, 3.5720001696608961, 3.574000169755891, 
    3.5760001698508859, 3.5780001699458808, 3.5800001700408757, 
    3.5820001701358706, 3.5840001702308655, 3.5860001703258604, 
    3.5880001704208553, 3.5900001705158502, 3.5920001706108451, 
    3.59400017070584, 3.5960001708008349, 3.5980001708958298, 
    3.6000001709908247, 3.6020001710858196, 3.6040001711808145, 
    3.6060001712758094, 3.6080001713708043, 3.6100001714657992, 
    3.6120001715607941, 3.614000171655789, 3.6160001717507839, 
    3.6180001718457788, 3.6200001719407737, 3.6220001720357686, 
    3.6240001721307635, 3.6260001722257584, 3.6280001723207533, 
    3.6300001724157482, 3.6320001725107431, 3.634000172605738, 
    3.6360001727007329, 3.6380001727957278, 3.6400001728907228, 
    3.6420001729857177, 3.6440001730807126, 3.6460001731757075, 
    3.6480001732707024, 3.6500001733656973, 3.6520001734606922, 
    3.6540001735556871, 3.656000173650682, 3.6580001737456769, 
    3.6600001738406718, 3.6620001739356667, 3.6640001740306616, 
    3.6660001741256565, 3.6680001742206514, 3.6700001743156463, 
    3.6720001744106412, 3.6740001745056361, 3.676000174600631, 
    3.6780001746956259, 3.6800001747906208, 3.6820001748856157, 
    3.6840001749806106, 3.6860001750756055, 3.6880001751706004, 
    3.6900001752655953, 3.6920001753605902, 3.6940001754555851, 
    3.69600017555058, 3.6980001756455749, 3.7000001757405698, 
    3.7020001758355647, 3.7040001759305596, 3.7060001760255545, 
    3.7080001761205494, 3.7100001762155443, 3.7120001763105392, 
    3.7140001764055341, 3.7160001765005291, 3.718000176595524, 
    3.7200001766905189, 3.7220001767855138, 3.7240001768805087, 
    3.7260001769755036, 3.7280001770704985, 3.7300001771654934, 
    3.7320001772604883, 3.7340001773554832, 3.7360001774504781, 
    3.738000177545473, 3.7400001776404679, 3.7420001777354628, 
    3.7440001778304577, 3.7460001779254526, 3.7480001780204475, 
    3.7500001781154424, 3.7520001782104373, 3.7540001783054322, 
    3.7560001784004271, 3.758000178495422, 3.7600001785904169, 
    3.7620001786854118, 3.7640001787804067, 3.7660001788754016, 
    3.7680001789703965, 3.7700001790653914, 3.7720001791603863, 
    3.7740001792553812, 3.7760001793503761, 3.778000179445371, 
    3.7800001795403659, 3.7820001796353608, 3.7840001797303557, 
    3.7860001798253506, 3.7880001799203455, 3.7900001800153404, 
    3.7920001801103354, 3.7940001802053303, 3.7960001803003252, 
    3.7980001803953201, 3.800000180490315, 3.8020001805853099, 
    3.8040001806803048, 3.8060001807752997, 3.8080001808702946, 
    3.8100001809652895, 3.8120001810602844, 3.8140001811552793, 
    3.8160001812502742, 3.8180001813452691, 3.820000181440264, 
    3.8220001815352589, 3.8240001816302538, 3.8260001817252487, 
    3.8280001818202436, 3.8300001819152385, 3.8320001820102334, 
    3.8340001821052283, 3.8360001822002232, 3.8380001822952181, 
    3.840000182390213, 3.8420001824852079, 3.8440001825802028, 
    3.8460001826751977, 3.8480001827701926, 3.8500001828651875, 
    3.8520001829601824, 3.8540001830551773, 3.8560001831501722, 
    3.8580001832451671, 3.860000183340162, 3.8620001834351569, 
    3.8640001835301518, 3.8660001836251467, 3.8680001837201416, 
    3.8700001838151366, 3.8720001839101315, 3.8740001840051264, 
    3.8760001841001213, 3.8780001841951162, 3.8800001842901111, 
    3.882000184385106, 3.8840001844801009, 3.8860001845750958, 
    3.8880001846700907, 3.8900001847650856, 3.8920001848600805, 
    3.8940001849550754, 3.8960001850500703, 3.8980001851450652, 
    3.9000001852400601, 3.902000185335055, 3.9040001854300499, 
    3.9060001855250448, 3.9080001856200397, 3.9100001857150346, 
    3.9120001858100295, 3.9140001859050244, 3.9160001860000193, 
    3.9180001860950142, 3.9200001861900091, 3.922000186285004, 
    3.9240001863799989, 3.9260001864749938, 3.9280001865699887, 
    3.9300001866649836, 3.9320001867599785, 3.9340001868549734, 
    3.9360001869499683, 3.9380001870449632, 3.9400001871399581, 
    3.942000187234953, 3.9440001873299479, 3.9460001874249429, 
    3.9480001875199378, 3.9500001876149327, 3.9520001877099276, 
    3.9540001878049225, 3.9560001878999174, 3.9580001879949123, 
    3.9600001880899072, 3.9620001881849021, 3.964000188279897, 
    3.9660001883748919, 3.9680001884698868, 3.9700001885648817, 
    3.9720001886598766, 3.9740001887548715, 3.9760001888498664, 
    3.9780001889448613, 3.9800001890398562, 3.9820001891348511, 
    3.984000189229846, 3.9860001893248409, 3.9880001894198358, 
    3.9900001895148307, 3.9920001896098256, 3.9940001897048205, 
    3.9960001897998154, 3.9980001898948103 ;

 octan =
  // octan(0, 0-7)
    "X+.Y+.Z+",
  // octan(1, 0-7)
    "X+.Y+.Z-",
  // octan(2, 0-7)
    "X+.Y-.Z+",
  // octan(3, 0-7)
    "X+.Y-.Z-",
  // octan(4, 0-7)
    "X-.Y+.Z+",
  // octan(5, 0-7)
    "X-.Y+.Z-",
  // octan(6, 0-7)
    "X-.Y-.Z+",
  // octan(7, 0-7)
    "X-.Y-.Z-" ;

 qvectors_statistics =
  // qvectors_statistics(0, 0-7)
    3, 5, 3, 8, 4, 9, 6, 12,
  // qvectors_statistics(1, 0-7)
    4, 4, 6, 7, 5, 10, 5, 9,
  // qvectors_statistics(2, 0-7)
    2, 7, 8, 4, 7, 5, 6, 11,
  // qvectors_statistics(3, 0-7)
    5, 3, 4, 8, 7, 7, 9, 7,
  // qvectors_statistics(4, 0-7)
    8, 6, 3, 8, 4, 6, 8, 7,
  // qvectors_statistics(5, 0-7)
    5, 6, 6, 9, 4, 3, 8, 9,
  // qvectors_statistics(6, 0-7)
    9, 5, 6, 6, 6, 6, 7, 5,
  // qvectors_statistics(7, 0-7)
    6, 2, 7, 10, 4, 8, 5, 8,
  // qvectors_statistics(8, 0-7)
    6, 3, 5, 12, 5, 5, 9, 5,
  // qvectors_statistics(9, 0-7)
    5, 2, 6, 7, 4, 6, 10, 10 ;

 Fqt-Na =
  // Fqt-Na(0, 0-1999)
    1, 0.9998595868110316, 0.99943932389916856, 0.99874210195617363, 
    0.99777265712740371, 0.99653747141926985, 0.99504464090240008, 
    0.99330371946595286, 0.99132554411719342, 0.98912204914742874, 
    0.98670607585124015, 0.98409118252936423, 0.98129145984310762, 
    0.97832135525936925, 0.97519550860782478, 0.97192860053303087, 
    0.96853521448547886, 0.96502971410810645, 0.96142613269985111, 
    0.95773807745872686, 0.95397864633356499, 0.95016035803036003, 
    0.94629509599435291, 0.94239406465786857, 0.93846776141776189, 
    0.93452595914949255, 0.93057769916620159, 0.92663129352142659, 
    0.92269433099329756, 0.91877369011553556, 0.91487555896082462, 
    0.91100545740170125, 0.90716826690025698, 0.90336825967982648, 
    0.89960913043552815, 0.89589402864859247, 0.89222559138970925, 
    0.88860597625341176, 0.88503689433476473, 0.88151964433254115, 
    0.8780551446779874, 0.8746439688797043, 0.87128637813637955, 
    0.86798235587830286, 0.86473164071075714, 0.86153375866918624, 
    0.8583880525004135, 0.85529370996556375, 0.85224978899826431, 
    0.84925524018838816, 0.8463089251745759, 0.84340963505443411, 
    0.84055610505670864, 0.83774702828596592, 0.8349810656510237, 
    0.83225685738236765, 0.82957302893580687, 0.82692819847163368, 
    0.8243209829064837, 0.82175000382620567, 0.81921389074454576, 
    0.81671128552046346, 0.81424084609958947, 0.81180124712485802, 
    0.8093911854674235, 0.80700938385372645, 0.80465459694214703, 
    0.80232561823994653, 0.8000212864684012, 0.79774049110873146, 
    0.79548217503616825, 0.79324533568327982, 0.79102902352439097, 
    0.78883233737890857, 0.78665441974838135, 0.78449445096230486, 
    0.78235164504295074, 0.7802252444991602, 0.77811451615631488, 
    0.77601874979722796, 0.77393725403728364, 0.77186935617637276, 
    0.76981439988140699, 0.76777174494798472, 0.7657407666942313, 
    0.76372085677100299, 0.76171142246364043, 0.75971188932428602, 
    0.75772170340423484, 0.75574033244939698, 0.75376727071606853, 
    0.75180204226701808, 0.74984420378142413, 0.74789334900545645, 
    0.74594911344428716, 0.74401117835475317, 0.742079274886004, 
    0.74015318634923166, 0.73823274899999758, 0.73631785081205459, 
    0.73440842772960946, 0.73250446108733847, 0.73060597155890517, 
    0.72871301514454712, 0.7268256784612902, 0.72494407473047795, 
    0.72306833736950837, 0.72119861640984528, 0.71933507457976498, 
    0.7174778813230176, 0.71562721142690189, 0.71378324024535333, 
    0.71194614313102755, 0.71011609216183391, 0.70829325552959155, 
    0.70647779397463217, 0.70466985851603159, 0.70286958713180647, 
    0.70107710386461453, 0.69929251718582652, 0.69751592174621657, 
    0.69574740199562701, 0.69398703530582984, 0.69223489515745829, 
    0.69049105218441154, 0.6887555739914194, 0.6870285243975639, 
    0.68530996184461834, 0.68359993620158788, 0.68189848645067197, 
    0.68020563923554367, 0.67852141045158187, 0.67684580391848237, 
    0.67517881487458886, 0.67352042929492417, 0.67187062694555022, 
    0.67022938253462117, 0.66859666475584434, 0.66697243889056335, 
    0.66535666662815285, 0.66374930780222496, 0.66215032016591957, 
    0.66055965920990445, 0.65897727718261156, 0.65740312459626871, 
    0.65583714693458062, 0.65427928419566528, 0.65272946939582355, 
    0.65118762500560268, 0.6496536597165713, 0.64812746585741166, 
    0.64660891707830759, 0.64509786685254189, 0.6435941510279114, 
    0.64209758673608985, 0.64060797986048923, 0.63912512664353827, 
    0.63764881933616735, 0.63617884954463333, 0.63471501340561987, 
    0.63325711424522813, 0.63180496520880403, 0.63035839127652182, 
    0.62891723020260371, 0.62748133245224513, 0.62605055979698376, 
    0.62462478641274022, 0.62320389626867778, 0.62178778469160911, 
    0.62037635873029473, 0.61896953812889421, 0.61756725768292098, 
    0.61616946698887598, 0.61477612871431386, 0.61338721633130244, 
    0.61200271066633538, 0.61062259727412949, 0.6092468613935057, 
    0.60787548701877792, 0.60650845519110252, 0.60514574278881761, 
    0.60378732491442921, 0.60243317466619295, 0.6010832631648797, 
    0.59973756030276304, 0.59839603373471184, 0.59705864497682593, 
    0.59572534897769813, 0.5943960917524469, 0.59307080751771979, 
    0.59174941748515253, 0.59043183003497346, 0.58911794076912616, 
    0.58780763211669806, 0.58650077664293332, 0.58519724211466151, 
    0.58389689377562271, 0.58259960205828976, 0.58130524432259734, 
    0.58001370955336251, 0.57872489805569161, 0.57743872380937, 
    0.57615511598471758, 0.57487402203775184, 0.5735954049535289, 
    0.57231924851604954, 0.57104555444451699, 0.56977434246591874, 
    0.56850565043680412, 0.56723953065180088, 0.56597604869166718, 
    0.56471528053755915, 0.56345730982064557, 0.5622022243594591, 
    0.56095011281928975, 0.55970106442035006, 0.55845516406479878, 
    0.5572124915149842, 0.55597311889421486, 0.55473710884385363, 
    0.55350451147183677, 0.55227536201990013, 0.55104967984398157, 
    0.54982746591121856, 0.54860870063781564, 0.54739334408165996, 
    0.54618133543897263, 0.54497259264535369, 0.5437670132941238, 
    0.54256447520677631, 0.54136483743090524, 0.54016794149059677, 
    0.53897361057407678, 0.53778165185300109, 0.53659185687790178, 
    0.53540400346928907, 0.53421785743016603, 0.53303317677542628, 
    0.53184971478435084, 0.53066722260206067, 0.52948545526785085, 
    0.52830417302103949, 0.5271231447900554, 0.5259421500613678, 
    0.52476098247533198, 0.52357945158925157, 0.52239738823921367, 
    0.52121464441045051, 0.52003109842501671, 0.51884665637133875, 
    0.51766125426565957, 0.51647485808028648, 0.5152874617668961, 
    0.51409908759282241, 0.51290978401130094, 0.51171962486200595, 
    0.51052870986222432, 0.50933716445590704, 0.50814513885098789, 
    0.50695280731291059, 0.50576036646413536, 0.5045680334842807, 
    0.50337604057190954, 0.50218463146793002, 0.50099405400294983, 
    0.49980455567305593, 0.49861637360226557, 0.4974297316464189, 
    0.49624483373496264, 0.49506185993413476, 0.49388096459658998, 
    0.49270227415671797, 0.49152588889460863, 0.49035188493374282, 
    0.48918031471791712, 0.48801121318888513, 0.48684460234600618, 
    0.4856804937337163, 0.48451889313014473, 0.48335980420828206, 
    0.48220323083701772, 0.48104917953349025, 0.4798976622611133, 
    0.47874869706092987, 0.47760230998886499, 0.4764585363209512, 
    0.47531742039147146, 0.47417901690752684, 0.47304338916333905, 
    0.47191061151292246, 0.4707807689165634, 0.46965395796018938, 
    0.46853028541114355, 0.46740986941436147, 0.46629283856851478, 
    0.46517933122103977, 0.46406949432957245, 0.46296348259964321, 
    0.46186145436217557, 0.46076357095314213, 0.45966999195412417, 
    0.45858087123427488, 0.45749635299377073, 0.45641656835983874, 
    0.45534162957574859, 0.45427162880998967, 0.45320663319231619, 
    0.4521466846345642, 0.4510918009559336, 0.450041980255453, 
    0.44899720439250507, 0.44795744486093142, 0.44692266694071081, 
    0.4458928350902675, 0.44486791609689474, 0.44384788518188634, 
    0.44283272939419133, 0.44182244837344248, 0.44081705916003472, 
    0.4398165953116176, 0.43882110997519824, 0.43783067094784561, 
    0.43684536339069435, 0.43586528638539934, 0.43489055063332999, 
    0.43392127728255997, 0.43295759607737305, 0.43199964337354274, 
    0.43104756066807987, 0.43010149279331483, 0.42916158387333142, 
    0.4282279741892443, 0.42730079556862599, 0.42638016633042219, 
    0.42546618632112904, 0.42455893382840443, 0.4236584630263015, 
    0.42276480247905796, 0.42187795576042342, 0.42099790341731314, 
    0.42012460580423544, 0.41925800525946999, 0.41839802849780977, 
    0.41754458950842538, 0.41669758798185985, 0.41585691080364351, 
    0.41502243018621987, 0.4141940053756768, 0.41337148139881075, 
    0.41255468941202794, 0.41174344599375401, 0.4109375558836515, 
    0.41013680649565587, 0.40934096782269308, 0.40854979050031626, 
    0.40776300191815346, 0.40698030612360042, 0.40620138654273669, 
    0.40542590703220432, 0.40465351714703585, 0.40388385541850996, 
    0.40311655435277022, 0.40235124401310673, 0.40158755739123747, 
    0.40082513695758376, 0.4000636408954053, 0.3993027502373217, 
    0.39854217427825811, 0.39778165486115769, 0.3970209678449213, 
    0.39625992242536501, 0.39549835883366669, 0.39473614487475683, 
    0.39397317280203153, 0.39320935637815652, 0.39244463035854493, 
    0.391678948222694, 0.39091228171807468, 0.39014462219460977, 
    0.38937597617188957, 0.38860636520076974, 0.38783582266445915, 
    0.38706439134812015, 0.38629211873760438, 0.3855190559913016, 
    0.38474525629108897, 0.38397077106383559, 0.38319564656986188, 
    0.38241992552438453, 0.38164364389400579, 0.38086683432361562, 
    0.38008952862914153, 0.37931176268880024, 0.37853357655839354, 
    0.37775501601663092, 0.37697612729869523, 0.37619695909836359, 
    0.37541755838603202, 0.37463797149071082, 0.37385824618324021, 
    0.37307843171254579, 0.3722985822553494, 0.37151875843918103, 
    0.37073902736147279, 0.36995946060789747, 0.36918013390203219, 
    0.3684011204422018, 0.36762248925478819, 0.36684429944617319, 
    0.36606659810061759, 0.36528941562518741, 0.36451276657455095, 
    0.36373664831808683, 0.36296104379371547, 0.36218592491624657, 
    0.36141125971061971, 0.3606370188435189, 0.3598631825251708, 
    0.35908974677319139, 0.35831672767531247, 0.35754416246728127, 
    0.3567721097834905, 0.35600064501648154, 0.35522985586102901, 
    0.35445983884419863, 0.35369069256223457, 0.35292251355546372, 
    0.35215539321416939, 0.35138941588142741, 0.35062466122523073, 
    0.34986120539551135, 0.34909912706476676, 0.34833850656074444, 
    0.34757942915341677, 0.34682198217622007, 0.34606625453045531, 
    0.34531233259293592, 0.34456029971407437, 0.34381023342568634, 
    0.34306220465637893, 0.34231627576111456, 0.34157249903400344, 
    0.34083091444996932, 0.34009154898803506, 0.33935441133627153, 
    0.33861949152294185, 0.33788675723482064, 0.33715615188019554, 
    0.33642759447968429, 0.33570098193641268, 0.33497619464464368, 
    0.3342531053410373, 0.33353158844185504, 0.33281153194274565, 
    0.33209284095408692, 0.33137544257502471, 0.3306592848215365, 
    0.3299443332245714, 0.32923056759346064, 0.32851797714385084, 
    0.32780655642346346, 0.32709630105260196, 0.32638720506168512, 
    0.32567925977567558, 0.3249724556084963, 0.32426678405707654, 
    0.32356224305905695, 0.3228588411604707, 0.32215660282762393, 
    0.3214555717752553, 0.32075581399363545, 0.32005741873432553, 
    0.31936049855498944, 0.31866518688534429, 0.31797163842608722, 
    0.31728002491264085, 0.31659053257331649, 0.31590335947636328, 
    0.31521871362104509, 0.31453680555544972, 0.31385784817095053, 
    0.31318205031540031, 0.31250961422857376, 0.31184073311797894, 
    0.31117558949965474, 0.31051435430954627, 0.30985718521743921, 
    0.30920422794635699, 0.30855561402612791, 0.30791146206992553, 
    0.3072718739999224, 0.30663693658297031, 0.30600671815238323, 
    0.30538126586727932, 0.30476060679979228, 0.30414474700427901, 
    0.30353367140382748, 0.30292734649976577, 0.30232571837835026, 
    0.30172871511385374, 0.30113624348481349, 0.30054819187358323, 
    0.29996442728420614, 0.2993847946711386, 0.29880911748796818, 
    0.29823719525594466, 0.29766880724746386, 0.2971037167914487, 
    0.29654167469414977, 0.29598242745000408, 0.29542572249258947, 
    0.29487131409342043, 0.2943189670749185, 0.29376845989174288, 
    0.2932195875258029, 0.29267216461845674, 0.29212602425696743, 
    0.29158102052255264, 0.29103702866925957, 0.29049394375026016, 
    0.28995168129387067, 0.2894101736446853, 0.28886937030799209, 
    0.28832923711466918, 0.28778975549307834, 0.28725092366083482, 
    0.28671275559280812, 0.28617528052498575, 0.28563853864284561, 
    0.28510258071746125, 0.28456746258453569, 0.28403324442580713, 
    0.28349998910383478, 0.28296776185550548, 0.28243662989392515, 
    0.28190666250625845, 0.28137792906122122, 0.28085049996139372, 
    0.28032444439999304, 0.27979982785679669, 0.27927671129226933, 
    0.27875515072561352, 0.27823519527673918, 0.27771689197166205, 
    0.27720028619114934, 0.27668542432881754, 0.27617235753841163, 
    0.2756611428153477, 0.27515184395790498, 0.27464453079748141, 
    0.27413927854531001, 0.27363616409191777, 0.27313526133935023, 
    0.27263664004857441, 0.2721403592948638, 0.27164646425895561, 
    0.2711549834966156, 0.27066592714419691, 0.27017928684348164, 
    0.26969503624635549, 0.26921313417729009, 0.26873352559651315, 
    0.26825614567432859, 0.26778091907675666, 0.26730776504499387, 
    0.26683659588578934, 0.26636732119970113, 0.26589984868541916, 
    0.26543408639646998, 0.26496994375571475, 0.26450733524046804, 
    0.26404617888979753, 0.2635863997385835, 0.26312792939060736, 
    0.26267070654901908, 0.26221467719316721, 0.26175979101217062, 
    0.26130600239076235, 0.26085326485076715, 0.2604015312310583, 
    0.25995074941171903, 0.25950086188421001, 0.25905180776718556, 
    0.25860352343578791, 0.25815594658154406, 0.25770901955952347, 
    0.25726269456927908, 0.25681693448426363, 0.2563717148482812, 
    0.25592702250300331, 0.25548285398695991, 0.25503921327139084, 
    0.2545961096290032, 0.25415355504627679, 0.25371156316188115, 
    0.2532701462884675, 0.25282931418500532, 0.25238907109136788, 
    0.25194941294243528, 0.25151032528277323, 0.25107177910172884, 
    0.25063373202662748, 0.25019612655062407, 0.24975889087112413, 
    0.24932194115142187, 0.24888518606273821, 0.24844853218707841, 
    0.24801189152601338, 0.24757518675428633, 0.2471383607154822, 
    0.24670137925452271, 0.24626423455112301, 0.24582694797032281, 
    0.24538956511966456, 0.2449521548164903, 0.24451480684089402, 
    0.24407762628045787, 0.24364073003279571, 0.2432042429628109, 
    0.24276829393449778, 0.24233301147160535, 0.24189852207466889, 
    0.24146494589501841, 0.24103239512910521, 0.2406009738667208, 
    0.24017077487783631, 0.23974188123421555, 0.23931436574374021, 
    0.23888828750446897, 0.23846369312339083, 0.23804061456620085, 
    0.23761906733177365, 0.23719905125032101, 0.23678055177971172, 
    0.2363635399185727, 0.23594797672435047, 0.23553381425193018, 
    0.23512100105943765, 0.23470948208523368, 0.23429920214475228, 
    0.2338901090685705, 0.23348215096539393, 0.23307528117474155, 
    0.23266945453445842, 0.23226463062181998, 0.23186077077349418, 
    0.2314578390551566, 0.23105580243678131, 0.23065462918626511, 
    0.23025428891739869, 0.22985475206331143, 0.22945598888537574, 
    0.22905796919358193, 0.22866066138140309, 0.22826403039990228, 
    0.22786803872734507, 0.22747264398898853, 0.22707779741701065, 
    0.22668344311991045, 0.22628951600218519, 0.22589594106022379, 
    0.22550263262408379, 0.22510949557591606, 0.22471642781027448, 
    0.22432332490278684, 0.22393008270516337, 0.22353660242409623, 
    0.22314279205607496, 0.22274856991300815, 0.22235386614122729, 
    0.22195862310188438, 0.22156279783179494, 0.22116636237753245, 
    0.22076930088761634, 0.22037161030451874, 0.21997329696979195, 
    0.21957437339229544, 0.21917485419951807, 0.21877475453615386, 
    0.21837408645831488, 0.21797285485418538, 0.21757105811687363, 
    0.21716868708203646, 0.21676572680515066, 0.21636215759243693, 
    0.21595796158015121, 0.21555312732512322, 0.21514765614312606, 
    0.21474156665624078, 0.21433489976475853, 0.21392772201745316, 
    0.21352013040413359, 0.21311225377484566, 0.21270425072598784, 
    0.21229630559237017, 0.21188861937634962, 0.2114814006545761, 
    0.21107485819312605, 0.21066919534157677, 0.21026461042460168, 
    0.2098612987980033, 0.20945945333406069, 0.2090592657345437, 
    0.20866092689942292, 0.20826462442096377, 0.20787054083870579, 
    0.20747885265261701, 0.20708972446012386, 0.20670330910458978, 
    0.20631974530277897, 0.20593915513062833, 0.20556164308564126, 
    0.20518729478733375, 0.20481617668400703, 0.20444833355118902, 
    0.20408378942413624, 0.20372254695063641, 0.20336458753963058, 
    0.20300987138034832, 0.20265833951705986, 0.20230991448990701, 
    0.20196450105303831, 0.2016219873643896, 0.20128224557885419, 
    0.20094513033807754, 0.20061047876587315, 0.20027810835720178, 
    0.19994781452854635, 0.19961937286748446, 0.19929253774262401, 
    0.19896704784999086, 0.19864262794753829, 0.19831899276960391, 
    0.1979958524744477, 0.19767291388150079, 0.19734988385679766, 
    0.19702647461078496, 0.19670240788836224, 0.1963774204162641, 
    0.19605126793028041, 0.19572373282098104, 0.19539462636335961, 
    0.19506379182228242, 0.19473110557402978, 0.1943964753189763, 
    0.19405983976652369, 0.19372116407436346, 0.19338043771005503, 
    0.19303767049198833, 0.19269288929857978, 0.19234613029750203, 
    0.19199743396489297, 0.19164684043887564, 0.19129438126760559, 
    0.19094007914423949, 0.19058394423162273, 0.19022597645979891, 
    0.18986616626314518, 0.18950449791020074, 0.18914095264942948, 
    0.18877551137794341, 0.18840815816785203, 0.18803888333727264, 
    0.18766768624004582, 0.18729457755371018, 0.18691958262347053, 
    0.18654274289829822, 0.18616411572820707, 0.18578377488734146, 
    0.18540180711107099, 0.18501831015874223, 0.18463338840834775, 
    0.18424714861264163, 0.18385969713372766, 0.18347113650797869, 
    0.18308156394114963, 0.18269107100775187, 0.18229974717225705, 
    0.18190767985262379, 0.18151495831043726, 0.18112167678132579, 
    0.18072793721207928, 0.18033385054915146, 0.17993953972976012, 
    0.17954513879481132, 0.17915079446442189, 0.17875666541711127, 
    0.17836292165266007, 0.17796974435286828, 0.17757732370423934, 
    0.17718585831616657, 0.17679555097866706, 0.17640660835766125, 
    0.17601923649423495, 0.17563364145834257, 0.1752500247994353, 
    0.17486858392882659, 0.17448950893919288, 0.17411298300138198, 
    0.17373917816747697, 0.17336825691670776, 0.17300036653919815, 
    0.17263563999456744, 0.17227419152389611, 0.1719161158357928, 
    0.17156148344502214, 0.17121033783722323, 0.17086269415386574, 
    0.17051853661631663, 0.17017781467712131, 0.16984044137029641, 
    0.16950629269987361, 0.16917520780203682, 0.16884699212524321, 
    0.16852141847353616, 0.16819823246429783, 0.16787715663300945, 
    0.16755789405473345, 0.16724013165416304, 0.16692354852078417, 
    0.16660781807574743, 0.16629261293902259, 0.16597761267552014, 
    0.16566250877536801, 0.1653470079881405, 0.16503083685832506, 
    0.16471374279301682, 0.16439549343153675, 0.16407588057475286, 
    0.16375471874269454, 0.16343184887880088, 0.1631071376088607, 
    0.16278047893473072, 0.1624517913879118, 0.1621210175409396, 
    0.16178812036822432, 0.16145308237826173, 0.16111590352194397, 
    0.1607765977420533, 0.1604351907886544, 0.16009172180230427, 
    0.15974623653981604, 0.15939878922260603, 0.15904943780813299, 
    0.15869824452526171, 0.15834526952283492, 0.15799057257252422, 
    0.15763420967282613, 0.15727623255493556, 0.15691668766678191, 
    0.15655561916900299, 0.15619306992669174, 0.15582908611362495, 
    0.15546371912362611, 0.15509702876430004, 0.15472908531783042, 
    0.15435997234708118, 0.1539897837414177, 0.15361862619723665, 
    0.15324661992592867, 0.15287389866214679, 0.15250061509823268, 
    0.15212694000150193, 0.15175306590429166, 0.1513792039398078, 
    0.15100558195578367, 0.1506324418971621, 0.15026003334259647, 
    0.14988860788753489, 0.14951841523537834, 0.1491496996147017, 
    0.14878269517572534, 0.14841762271303888, 0.14805468448086681, 
    0.14769406382712075, 0.14733592325839212, 0.14698040147549629, 
    0.14662761577852002, 0.14627766210437118, 0.14593061466973437, 
    0.14558652778545517, 0.1452454354515739, 0.14490735197519219, 
    0.14457227408962944, 0.14424017656126989, 0.14391101872375028, 
    0.14358474561736773, 0.14326128961983475, 0.14294057439737815, 
    0.14262251809748366, 0.14230703571332146, 0.141994040286959, 
    0.14168344406976502, 0.1413751605277194, 0.14106910225001315, 
    0.14076518167863988, 0.14046331245433949, 0.14016340846816708, 
    0.13986538862611578, 0.13956917656122433, 0.13927470502713221, 
    0.13898191946940003, 0.13869078149078004, 0.13840127282117815, 
    0.13811340127536395, 0.1378272054032561, 0.13754275804551297, 
    0.13726017194641149, 0.13697959764982778, 0.13670122348195735, 
    0.13642527096112703, 0.13615198845187604, 0.13588164686347459, 
    0.13561453058223141, 0.13535093539984411, 0.1350911621038729, 
    0.13483551161409785, 0.13458428254179128, 0.13433776629395738, 
    0.13409624434882975, 0.13385998366607763, 0.1336292333630677, 
    0.13340422013403375, 0.13318514394831571, 0.13297217445614337, 
    0.13276544640779447, 0.13256505756279516, 0.13237106612421917, 
    0.13218348878906366, 0.1320023021390011, 0.13182744140487662, 
    0.13165880369823257, 0.13149624823992145, 0.13133959993082811, 
    0.13118865282063288, 0.13104317303792831, 0.13090290126606968, 
    0.13076755678700633, 0.13063684056657812, 0.13051043899022724, 
    0.13038803004959276, 0.13026928521069464, 0.1301538749482096, 
    0.13004147328053881, 0.12993176100371948, 0.12982442532667149, 
    0.12971916440237316, 0.12961568619309252, 0.1295137102754588, 
    0.12941296715270739, 0.12931319957875381, 0.12921416230767821, 
    0.12911562142998056, 0.12901735549711738, 0.12891915301280449, 
    0.12882081272955809, 0.12872214105285748, 0.12862295138544211, 
    0.1285230637515262, 0.12842230465840082, 0.12832050956797134, 
    0.12821752336939377, 0.12811320407913873, 0.12800742745480137, 
    0.12790008566032443, 0.12779109109167971, 0.12768037752608888, 
    0.12756790039940458, 0.12745363729887021, 0.12733758543180396, 
    0.12721976344984914, 0.12710020557131563, 0.12697896113850982, 
    0.12685609061700912, 0.12673166172378483, 0.12660574688326404, 
    0.12647841772626223, 0.12634974397657381, 0.12621979115274842, 
    0.12608862145339061, 0.12595629571708253, 0.12582287366772182, 
    0.1256884212241037, 0.12555301034136404, 0.12541672131316381, 
    0.12527964473532574, 0.12514187648557565, 0.12500351627788975, 
    0.12486466189144359, 0.12472540446201262, 0.12458582153460432, 
    0.12444597347594877, 0.12430590201036605, 0.12416562623247625, 
    0.1240251423847267, 0.12388442392276265, 0.12374341984715277, 
    0.12360205545405351, 0.12346023292737596, 0.12331783283000464, 
    0.12317471494740301, 0.12303072336554954, 0.12288568720620671, 
    0.12273943063300348, 0.12259177522780804, 0.12244254966813624, 
    0.12229159716830917, 0.12213878210564737, 0.12198399779599771, 
    0.12182717153737602, 0.12166827119109132, 0.12150730721726344, 
    0.12134433078153541, 0.12117943339511542, 0.12101273806998404, 
    0.12084439275984654, 0.12067455855057287, 0.12050340327780645, 
    0.1203310907672021, 0.12015777381854126, 0.1199835889330472, 
    0.11980865382079302, 0.11963306365354778, 0.11945689256945224, 
    0.11928019464853126, 0.11910300400971695, 0.11892533922511901, 
    0.11874720754812987, 0.11856860498115478, 0.11838952290788794, 
    0.11820995027097488, 0.11802987819792937, 0.11784930222965882, 
    0.11766822652125031, 0.11748666776030967, 0.11730465732721421, 
    0.11712224248605183, 0.11693949049916921, 0.11675648573643815, 
    0.11657332964858629, 0.11639013796267372, 0.11620703662748255, 
    0.11602415741627084, 0.11584163221481197, 0.11565959139501365, 
    0.11547815913231335, 0.11529744850670545, 0.11511756407497063, 
    0.11493859755596755, 0.11476062910466196, 0.11458372639019965, 
    0.11440794793236836, 0.11423334020180921, 0.11405994118592161, 
    0.11388778262687439, 0.11371689115800908, 0.11354729082643115, 
    0.11337900235651388, 0.11321204291571799, 0.11304642668296727, 
    0.11288216047131296, 0.11271924474403833, 0.11255766923300554, 
    0.11239740881945039, 0.1122384193211528, 0.11208063251889266, 
    0.11192395053094235, 0.11176824701694973, 0.11161336880386181, 
    0.11145913712810852, 0.11130535407184879, 0.11115180950210923, 
    0.11099828457022708, 0.11084455855120789, 0.11069041421438343, 
    0.1105356410797894, 0.11038003852200214, 0.11022341820898734, 
    0.11006560370335466, 0.10990642852120917, 0.10974573468111438, 
    0.10958337044857154, 0.10941918632855102, 0.10925303318831744, 
    0.1090847635523295, 0.10891423290651538, 0.1087413021565128, 
    0.10856584320303188, 0.10838774147326431, 0.10820689903192116, 
    0.1080232331336618, 0.10783667853301784, 0.10764718253434592, 
    0.10745470409938096, 0.10725921145342764, 0.10706067788633938, 
    0.10685908030803834, 0.10665439704258492, 0.10644660564073574, 
    0.10623568218730771, 0.1060216012636513, 0.10580433630386354, 
    0.10558386093393984, 0.1053601502742976, 0.10513318188778531, 
    0.10490293973630424, 0.10466941371180806, 0.10443260069225115, 
    0.10419250722974538, 0.10394915150177982, 0.10370256337156789, 
    0.10345278977885902, 0.10319989438883248, 0.10294396350405706, 
    0.10268510852991593, 0.10242346939411101, 0.10215921669271194, 
    0.1018925513909656, 0.10162370572595228, 0.10135293917447714, 
    0.10108053586314676, 0.10080679871804157, 0.10053204436069108, 
    0.10025659605303718, 0.099980778422317354, 0.099704912019353747, 
    0.099429307582834595, 0.099154263015780369, 0.098880060334386621, 
    0.098606962488188496, 0.098335212188427293, 0.098065031670972413, 
    0.097796621644163903, 0.097530164863772667, 0.097265823095548432, 
    0.097003742579136756, 0.096744051609087944, 0.096486861407305169, 
    0.096232267114847406, 0.095980347772197397, 0.095731165313404018, 
    0.095484769761655375, 0.095241197357540691, 0.095000477009795456, 
    0.094762630829327496, 0.094527676606891015, 0.094295628425683481, 
    0.094066497938852037, 0.093840293653248391, 0.093617021134117448, 
    0.093396683462941221, 0.093179281832663191, 0.092964814027812814, 
    0.092753274272687425, 0.092544652081676088, 0.092338930425247823, 
    0.092136083965548468, 0.091936079099028789, 0.091738872978383831, 
    0.091544412885915111, 0.09135263608942118, 0.091163472232995021, 
    0.090976843444983635, 0.090792668025417148, 0.090610863244481213, 
    0.090431345576484107, 0.090254032636091094, 0.09007884352641525, 
    0.089905696773167759, 0.08973450656712291, 0.08956518118448413, 
    0.089397622908523766, 0.089231726391336572, 0.089067381240865384, 
    0.088904472359967582, 0.08874288519324626, 0.088582504544058388, 
    0.088423217508913354, 0.088264914175301579, 0.0881074893574572, 
    0.087950842969862664, 0.087794882166487884, 0.087639524093936244, 
    0.087484700041161517, 0.087330356443861418, 0.087176461266961283, 
    0.087023003042973446, 0.086869995919290233, 0.086717478098738823, 
    0.08656551160891883, 0.086414182901534978, 0.086263600202497168, 
    0.086113890329161003, 0.085965198048337688, 0.085817681095987475, 
    0.085671507308034453, 0.085526851191858697, 0.085383891335377687, 
    0.085242804855579751, 0.08510376848494805, 0.084966955424848889, 
    0.084832536176114956, 0.084700680147826501, 0.084571555781382521, 
    0.084445329050784002, 0.084322159656022758, 0.084202197673791335, 
    0.084085577917545895, 0.083972415095712599, 0.083862804182431416, 
    0.083756814870765334, 0.083654492780197487, 0.083555857507544129, 
    0.083460901838410095, 0.083369588234243494, 0.083281848871671255, 
    0.083197582520850411, 0.083116652626139445, 0.083038892259069463, 
    0.082964102198121767, 0.082892055847388402, 0.082822501764708206, 
    0.082755170900145752, 0.082689774004257421, 0.082626008876269794, 
    0.082563560356166965, 0.082502100439496698, 0.082441291148440718, 
    0.082380781162279093, 0.082320210925126369, 0.082259213785224689, 
    0.082197417303615516, 0.082134450172859377, 0.082069946223169959, 
    0.082003549107398765, 0.081934916900453778, 0.081863724879069497, 
    0.081789668139182328, 0.081712463291327572, 0.081631850547903409, 
    0.081547597163551241, 0.081459497394251443, 0.081367378001623025, 
    0.081271096317565863, 0.081170546004796298, 0.081065652971087337, 
    0.080956377033977692, 0.080842708238620803, 0.080724663984413969, 
    0.080602284789636533, 0.08047562954436896, 0.080344774076700237, 
    0.080209802652293105, 0.080070805713617244, 0.079927873263011817, 
    0.079781091140733756, 0.079630534643236578, 0.079476271158134146, 
    0.079318356478016411, 0.079156841095790992, 0.078991773691736294, 
    0.078823203789322255, 0.078651186771582907, 0.078475786554504059, 
    0.078297076721275782, 0.078115146489668233, 0.077930099600279787, 
    0.077742060787189038, 0.077551173621751207, 0.077357600200719245, 
    0.07716151651781851, 0.076963108195722496, 0.076762568098976913, 
    0.076560087777790095, 0.076355853146449479, 0.076150036789472617, 
    0.07594279658029969, 0.075734266631735422, 0.075524553329663013, 
    0.075313730173720256, 0.075101835223475202, 0.074888870581186179, 
    0.074674805498591595, 0.074459582495221527, 0.074243124295880064, 
    0.074025346960964161, 0.073806167240267326, 0.073585516795639447, 
    0.07336334439175779, 0.073139625075709036, 0.072914355502373976, 
    0.07268755724518168, 0.072459270776394191, 0.072229551860309243, 
    0.071998466266010169, 0.071766082045018012, 0.071532467119030677, 
    0.071297680953901627, 0.071061774280862841, 0.070824782739388928, 
    0.070586730954939281, 0.070347632352875888, 0.070107494108430923, 
    0.069866322373212053, 0.06962412732278439, 0.069380928848706919, 
    0.069136763441659824, 0.0688916901356737, 0.068645801118678448, 
    0.068399225730508315, 0.06815213654654291, 0.067904749148718718, 
    0.06765731935591783, 0.0674101362388565, 0.067163519381949005, 
    0.066917811707895833, 0.06667337381171598, 0.066430581622306722, 
    0.066189819610370626, 0.065951471397416569, 0.065715917329985704, 
    0.065483524016446859, 0.065254633209934645, 0.065029557375101854, 
    0.064808569742337133, 0.064591897228105349, 0.064379714619007697, 
    0.064172144843389928, 0.063969257173431132, 0.063771072941957802, 
    0.063577570398397204, 0.063388697880816358, 0.063204382713184112, 
    0.063024544319710371, 0.062849101592410334, 0.06267798157674899, 
    0.062511119985649649, 0.062348460405789959, 0.062189953513625496, 
    0.062035552589821005, 0.061885211327437899, 0.061738888791709232, 
    0.061596545904492046, 0.061458150279759101, 0.061323674275349856, 
    0.061193091448989628, 0.061066367542445738, 0.06094345165738841, 
    0.060824267305110161, 0.060708706577811168, 0.060596625332599283, 
    0.060487846803202308, 0.060382162623712758, 0.060279335324400642, 
    0.06017911068942336, 0.06008122428447478, 0.05998541225582988, 
    0.059891420170123798, 0.059799014929156249, 0.059707985116378245, 
    0.059618142279480056, 0.059529320481473531, 0.059441370310272218, 
    0.059354155272996638, 0.059267548449287999, 0.059181428615498327, 
    0.059095681554100929, 0.059010204786722566, 0.05892490605833807, 
    0.058839710708298992, 0.058754564362587879, 0.058669434429152754, 
    0.05858431104839229, 0.058499205086929844, 0.058414143474355071, 
    0.058329163317861352, 0.058244310833548217, 0.05815963641331371, 
    0.058075191633006687, 0.057991032582554974, 0.057907221860327519, 
    0.057823830495640001, 0.057740940668823681, 0.05765864427768206, 
    0.057577039936335686, 0.05749623806434577, 0.057416354226150462, 
    0.057337511617583443, 0.057259841817677098, 0.057183483313578004, 
    0.057108582806412712, 0.057035291867534248, 0.056963769123700783, 
    0.05689417059672592, 0.056826651989716453, 0.056761360120651812, 
    0.056698430477792848, 0.056637981600869067, 0.056580109132162312, 
    0.056524885901033425, 0.056472357344127339, 0.056422541622389834, 
    0.056375426634853773, 0.056330972480260928, 0.05628911275499221, 
    0.056249753876510933, 0.056212780082683683, 0.056178056253492939, 
    0.056145440135066893, 0.05611478560042607, 0.05608595490490341, 
    0.056058825873784988, 0.056033293689320307, 0.056009276597375084, 
    0.055986713865549431, 0.055965564067898987, 0.055945804980508815, 
    0.055927428683234047, 0.055910442301654005, 0.055894867167941141, 
    0.055880734112680602, 0.055868087813303824, 0.055856982951048427, 
    0.055847488620620389, 0.055839685419548556, 0.055833665672119302, 
    0.055829535862239703, 0.055827413852061504, 0.055827431657512146, 
    0.055829732377471054, 0.055834466678546121, 0.05584179350008505, 
    0.055851870353148689, 0.055864856432649088, 0.05588090266293233, 
    0.055900152707689409, 0.055922736958470463, 0.055948772496415618, 
    0.055978363232188452, 0.056011598381155971, 0.056048551599363998, 
    0.05608927882017422, 0.056133820224951385, 0.056182194283448755, 
    0.056234396880420125, 0.05629039808371402, 0.056350141437655217, 
    0.056413545212095052, 0.056480500676525679, 0.056550879685497657, 
    0.056624532068032613, 0.056701290455748982, 0.056780974061418486, 
    0.056863390632738743, 0.05694833638657, 0.057035599278416484, 
    0.057124956500478233, 0.057216173198285855, 0.057309005493879552, 
    0.057403194513887562, 0.057498473226125592, 0.05759457044932681, 
    0.057691214712418767, 0.057788142733761233, 0.057885105931783802, 
    0.05798187440623661, 0.058078243448411143, 0.058174032904252014, 
    0.058269093663146261, 0.058363307090624268, 0.058456583729513012, 
    0.058548862117624369, 0.058640102281178226, 0.058730277489406811, 
    0.058819368634001314, 0.058907353875254857, 0.058994202541476234, 
    0.059079872537327605, 0.059164312270294069, 0.05924746736297172, 
    0.059329284932957749, 0.059409721580846085, 0.059488747104534209, 
    0.059566347997322591, 0.05964253184749458, 0.05971733198642977, 
    0.059790812951958518, 0.059863070835394536, 0.059934238058516255, 
    0.060004477876978012, 0.060073979335019831, 0.060142949505698304, 
    0.060211599726863699, 0.06028013665889189, 0.060348755305727267, 
    0.060417638145913104, 0.060486955675752276, 0.06055686970282749, 
    0.06062754051164064, 0.060699124544880273, 0.06077177046269603, 
    0.060845613828610173, 0.060920768904250931, 0.060997324983553709, 
    0.061075342489168016, 0.061154854591739236, 0.061235868898097637, 
    0.061318367632276265, 0.061402312346261867, 0.061487646226070343, 
    0.061574294914451162, 0.061662174953859096, 0.061751182861996129, 
    0.061841202459142687, 0.061932099239474882, 0.062023717739084383, 
    0.06211588166610537, 0.062208390103766532, 0.06230102047262847, 
    0.062393531870699126, 0.062485667672891272, 0.062577164187224352, 
    0.062667754399418296, 0.062757176970140743, 0.062845176684334314, 
    0.062931510489223394, 0.063015948563418522, 0.06309827616647716, 
    0.063178294638001856, 0.063255813732150043, 0.063330651108558692, 
    0.063402622987910745, 0.063471538075990638, 0.063537191156125675, 
    0.063599356620428177, 0.063657782309298139, 0.063712190991068951, 
    0.063762283052236912, 0.063807738770497113, 0.063848223867632767, 
    0.063883405931228918, 0.063912954844632483, 0.063936556930789645, 
    0.063953917024344165, 0.063964761784272614, 0.063968843742689824, 
    0.063965940355737341, 0.063955856678796524, 0.06393842259867652, 
    0.063913498786451389, 0.063880981675860343, 0.063840806447255996, 
    0.063792960338495228, 0.063737485319610807, 0.063674488180475053, 
    0.063604137261443205, 0.063526659162558105, 0.06344234030485299, 
    0.063351517539512334, 0.063254572925064409, 0.06315193461741854, 
    0.063044065336042787, 0.062931460584933985, 0.062814642003050536, 
    0.062694157696832897, 0.062570573896625833, 0.062444470338850068, 
    0.062316435343362786, 0.062187054350509453, 0.062056897497626357, 
    0.061926507932516729, 0.061796385813490777, 0.061666981061774075, 
    0.061538680616989451, 0.061411807508684003, 0.06128661739639147, 
    0.061163301105978757, 0.061041984004471909, 0.060922732507932634, 
    0.060805559876951951, 0.060690428505199817, 0.060577255037901706, 
    0.060465917858464467, 0.060356265698507161, 0.060248124466123917, 
    0.060141309396217951, 0.060035635226553377, 0.059930922054027683, 
    0.059827002877552909, 0.059723729134582383, 0.059620972739604566, 
    0.059518625660244087, 0.059416601202166061, 0.05931483625158257, 
    0.059213290934604201, 0.059111946464657929, 0.059010809163498379, 
    0.058909903741727686, 0.058809275748255833, 0.058708989293392452, 
    0.058609120738383737, 0.058509756491229033, 0.058410991196746254, 
    0.058312921578349872, 0.058215643602537157, 0.058119248284917546, 
    0.058023819337153504, 0.05792942831802364, 0.057836130934535213, 
    0.057743964854883062, 0.057652941038536659, 0.057563044613607811, 
    0.057474235737714541, 0.05738645952861178, 0.057299653298172222, 
    0.057213752137278723, 0.057128693145291565, 0.057044413943122936, 
    0.056960847878014052, 0.056877924896106567, 0.056795564195017731, 
    0.05671367813366323, 0.056632167541853837, 0.056550920504276764, 
    0.056469818943276413, 0.056388740123568586, 0.056307562008967728, 
    0.056226172458953554, 0.056144479777726262, 0.056062423279646646, 
    0.055979983606425129, 0.055897195367467969, 0.055814151276886548, 
    0.055731008125528149, 0.055647984533286232, 0.055565351947758752, 
    0.055483423500082896, 0.055402539449855702, 0.055323044281360541, 
    0.055245274103343546, 0.055169538431171596, 0.055096113262214662, 
    0.055025224682589212, 0.054957048014161104, 0.054891703882448198, 
    0.054829256065319285, 0.05476971531849225, 0.054713049466989891, 
    0.054659194017601165, 0.054608069241309593, 0.054559595317528825, 
    0.05451370244713926, 0.054470331636428448, 0.054429435416884227, 
    0.054390969423557645, 0.054354885713894775, 0.054321126713106349, 
    0.054289615075413834, 0.054260255916519132, 0.054232932737485536, 
    0.054207514011392816, 0.054183852872197784, 0.054161795029506507, 
    0.054141181629302301, 0.054121856105234116, 0.054103667362976074, 
    0.05408647785868876, 0.054070161815436571, 0.054054610403849623, 
    0.054039731231964573, 0.054025452154937544, 0.054011715134143663, 
    0.053998476646793574, 0.05398569980998761, 0.05397335626947343, 
    0.053961426381516457, 0.053949896256875976, 0.053938771731686208, 
    0.053928079882071399, 0.053917867179465326, 0.053908207844528724, 
    0.053899195959833723, 0.053890945657414799, 0.053883579068144984, 
    0.053877229932283832, 0.053872033805260712, 0.053868123373008461, 
    0.053865632356566419, 0.053864680469499444, 0.05386538357347246, 
    0.053867845623548169, 0.053872154766082772, 0.053878387808523623, 
    0.053886606956393412, 0.053896868284936179, 0.053909220338558488, 
    0.05392372042340441, 0.053940431104175963, 0.053959426459175279, 
    0.053980793414798396, 0.054004627843782516, 0.054031043517993448, 
    0.054060165404063061, 0.054092131093086179, 0.054127093994694786, 
    0.054165210056027036, 0.054206633815442606, 0.054251514544206028, 
    0.05429999319479311, 0.05435219093141113, 0.054408205633132013, 
    0.054468115508715255, 0.054531978034544827, 0.054599826097603242, 
    0.054671679255626625, 0.054747536103637646, 0.054827381919597337, 
    0.054911180404339337, 0.054998879152098182, 0.055090400775723657, 
    0.055185645044190192, 0.05528448210450778, 0.055386755568106585, 
    0.055492273053068877, 0.055600816094008604, 0.055712133146869271, 
    0.055825953609429622, 0.055941995045140525, 0.05605997566022531, 
    0.056179625772377256, 0.056300698721316718, 0.056422975095257816, 
    0.056546262435880221, 0.056670392214635261, 0.056795208356329417, 
    0.056920550790381698, 0.057046253431901756, 0.057172131621288563, 
    0.057297970452227516, 0.057423531983490476, 0.057548549379767777, 
    0.057672742942946713, 0.057795818879728296, 0.057917476677849841, 
    0.058037418276493592, 0.05815535073376165, 0.058270995437061462, 
    0.058384097779550725, 0.058494433071360236, 0.058601826509361576, 
    0.058706157950683825, 0.058807364727342992, 0.058905439909603965, 
    0.059000422611004626, 0.059092382751463765, 0.059181401670564543, 
    0.059267548439225097, 0.059350869272659132, 0.059431378429845146, 
    0.059509058798754108, 0.05958386983706733, 0.059655755007338516, 
    0.059724649545475857, 0.059790484928407009, 0.059853195907060328, 
    0.05991270783572223, 0.059968937824529819, 0.060021799982986464, 
    0.060071195496826192, 0.060117020834352608, 0.060159173786267561, 
    0.06019755910503672, 0.060232096090919243, 0.060262728821316398, 
    0.060289419098967741, 0.060312154525889457, 0.06033094511766348, 
    0.060345823834620616, 0.060356839140060674, 0.060364058732379516, 
    0.06036757084927509, 0.060367478988619015, 0.060363906968321002, 
    0.060356996932548812, 0.060346898710160787, 0.060333767548477524, 
    0.060317750054120545, 0.060298974688844868, 0.060277538606791393, 
    0.060253503452692231, 0.06022689987529331, 0.060197727762789768, 
    0.060165965443810317, 0.060131576666195535, 0.060094531807479964, 
    0.060054802857663778, 0.060012376458587015, 0.059967256828375747, 
    0.059919460732964398, 0.059869020997627913, 0.059815986115988248, 
    0.059760418635712242, 0.059702397461185788, 0.059642024822239924, 
    0.059579424080877137, 0.059514752029235833, 0.059448189150278698, 
    0.059379951685918655, 0.059310284350338444, 0.059239449566045772, 
    0.059167721777040938, 0.059095369321760557, 0.059022648399473146, 
    0.058949794911298224, 0.058877002000113011, 0.058804418745291173, 
    0.058732142363317134, 0.058660209646410798, 0.058588594133800014, 
    0.058517209789916737, 0.058445905290835688, 0.05837447668123405, 
    0.058302676903356825, 0.058230230959257986, 0.058156850242934176, 
    0.058082248647782338, 0.058006166492999785, 0.05792838407454768, 
    0.057848738575580899, 0.057767126563248582, 0.05768352093894185, 
    0.057597971500157823, 0.057510604297919078, 0.057421613877945345, 
    0.057331235317723647, 0.057239737994382985, 0.057147383429076042, 
    0.057054393443369412, 0.056960957463285097, 0.056867213970278954, 
    0.056773257393117497, 0.056679147162896182, 0.056584926933397395, 
    0.056490631962812156, 0.056396313336112058, 0.056302035207428013, 
    0.056207885507820084, 0.056113968483390085, 0.056020393939890917, 
    0.055927269913002176, 0.055834675010464296, 0.055742634216111087, 
    0.055651102932154216, 0.055559940370648951, 0.055468898024551246, 
    0.05537761487660512, 0.055285632232085644, 0.0551924042478181, 
    0.055097339247623396, 0.054999836259899328, 0.054899334823828014, 
    0.05479534636870919, 0.054687465455437102, 0.054575389714719508, 
    0.054458902474000481, 0.05433786220481255, 0.054212197295692481, 
    0.054081872180805339, 0.053946870899580002, 0.053807187490603835, 
    0.053662802876797047, 0.053513657851444296, 0.053359653293290538, 
    0.053200639969762216, 0.05303642890427572, 0.052866793301224506, 
    0.052691506125980919, 0.05251036367298071, 0.052323215981346871, 
    0.052129993145625483, 0.051930714451920761, 0.051725503093702004, 
    0.051514552270562709, 0.051298135809370357, 0.05107655009291056, 
    0.050850135899095129, 0.050619234226662042, 0.050384217023487936, 
    0.050145460411388135, 0.049903356178511035, 0.0496583028633047, 
    0.049410727396885665, 0.049161042760847803, 0.048909676335699703, 
    0.048657043015044678, 0.048403534005253122, 0.048149518074527199, 
    0.047895321640741721, 0.04764121560321162, 0.047387417547188976, 
    0.047134074607249186, 0.046881238557275579, 0.046628897472993314, 
    0.046376924140447605, 0.046125093287321589, 0.04587305788141962, 
    0.045620355904734219, 0.045366426470753472, 0.045110623044137044, 
    0.044852261046010679, 0.044590671126132048, 0.044325251636535848, 
    0.044055537384331468, 0.043781235980812551, 0.043502293168757082, 
    0.043218916909294011, 0.042931621356728331, 0.042641214895424502, 
    0.042348805585569103, 0.042055759036017368, 0.041763644991950143, 
    0.041474169344592297, 0.041189114432663494, 0.040910289058865956, 
    0.040639457829589096, 0.040378312235934105, 0.040128448545817375, 
    0.039891325943315049, 0.039668278747759925, 0.039460490841477465, 
    0.039269009736945047, 0.039094753348448787, 0.03893849146322681, 
    0.038800857442110863, 0.038682331768214777, 0.038583237067691636, 
    0.038503686744155753, 0.03844357806545879, 0.038402563588360465, 
    0.038380028977211475, 0.038375100878018938, 0.0383866357596577, 
    0.038413235320320607, 0.038453291063386401, 0.038505023793787382, 
    0.038566552122748794, 0.038635930331605117, 0.038711224906603309, 
    0.038790535765432572, 0.038872086174071903, 0.038954238035246044, 
    0.03903549230524641, 0.039114596885428538, 0.039190450730496901, 
    0.039262202697355961, 0.039329164313796787, 0.03939081619130861, 
    0.039446765526592778, 0.039496706688574801, 0.039540404738271577, 
    0.03957763067534685, 0.0396082213419219, 0.039632071054402154, 
    0.039649210545303938, 0.039659803031981161, 0.039664198584332712, 
    0.039662890459607039, 0.039656550208079067, 0.039645949456301822, 
    0.039631928467902894, 0.039615360326569288, 0.039597092952023641, 
    0.039577938776532512, 0.039558613177190068, 0.039539786933061399, 
    0.039522099351604285, 0.039506173649168981, 0.039492650312470061, 
    0.039482157341862084, 0.039475295310649403, 0.039472595926876686, 
    0.039474458037840804, 0.039481195567970723, 0.039493060074105482, 
    0.039510281480906677, 0.039533124369370252, 0.039561899044652987, 
    0.039597001094118074, 0.039638912369882352, 0.039688128350098398, 
    0.039745242192916773, 0.039810681970426295, 0.039884914654584533, 
    0.039968048914158102, 0.040059803719179193, 0.040159821871214564, 
    0.040267121852184319, 0.040380574797670543, 0.04049868875988729, 
    0.040619547269681124,
  // Fqt-Na(1, 0-1999)
    1, 0.99955259254148066, 0.99821429912965087, 0.99599677528966402, 
    0.99291910498154135, 0.98900734330458617, 0.98429391200729333, 
    0.97881688246281939, 0.9726191764032327, 0.96574771901188439, 
    0.95825257672070097, 0.95018610483745658, 0.9416021291075477, 
    0.93255517931407339, 0.923099786482521, 0.91328985145761465, 
    0.90317808827569013, 0.89281554820027498, 0.88225121284421826, 
    0.8715316648301088, 0.86070082423306304, 0.8497997511795119, 
    0.83886651274655488, 0.82793610341180324, 0.81704042465741511, 
    0.80620830449508929, 0.79546555636319616, 0.78483507019638787, 
    0.77433692139062005, 0.7639885005943724, 0.75380466275785751, 
    0.74379788112396572, 0.73397841811471254, 0.72435449190092771, 
    0.71493244581374171, 0.70571691319475605, 0.69671097842401408, 
    0.68791633128909391, 0.67933341584131579, 0.67096157367687781, 
    0.66279917716887449, 0.65484376211416462, 0.6470921468854649, 
    0.63954054959608042, 0.63218469143970901, 0.62501989329297813, 
    0.61804115728160447, 0.61124324309994893, 0.60462073257824966, 
    0.59816808797678855, 0.59187969731457979, 0.58574992164210182, 
    0.57977312880912379, 0.57394372732385623, 0.56825618818333024, 
    0.56270506944631637, 0.55728502801114665, 0.55199083152503048, 
    0.54681736711918671, 0.54175964889128081, 0.53681281752429122, 
    0.53197214310466368, 0.52723302754586554, 0.52259099879750426, 
    0.51804171796329179, 0.51358098063889202, 0.50920472498022673, 
    0.50490904226344169, 0.50069018707786483, 0.49654458534666124, 
    0.49246883748019443, 0.48845971782635678, 0.48451416942503955, 
    0.4806292921726143, 0.47680233191773469, 0.47303066867445859, 
    0.46931180603996298, 0.46564336137958484, 0.4620230571597056, 
    0.45844872040001911, 0.45491827545023289, 0.45142974700321747, 
    0.44798125905712438, 0.44457103956323574, 0.44119742367243892, 
    0.43785886208558228, 0.43455392455294889, 0.43128131040624168, 
    0.42803985361107755, 0.42482851947284378, 0.4216464059235594, 
    0.41849273595739445, 0.41536684921656319, 0.41226819546837884, 
    0.40919633104208974, 0.40615091832467365, 0.40313172189137758, 
    0.40013860603291412, 0.39717152645260151, 0.39423052066305669, 
    0.391315692862784, 0.38842720140571951, 0.38556524175368501, 
    0.38273003339299316, 0.37992180818448001, 0.37714079960401647, 
    0.37438723091004639, 0.37166130883173609, 0.36896321962523793, 
    0.36629312200685804, 0.36365114900521545, 0.361037405522591, 
    0.3584519739832262, 0.35589491254987943, 0.3533662610190208, 
    0.3508660383263647, 0.34839424072790715, 0.34595083750322109, 
    0.34353577124693901, 0.34114895545997787, 0.33879027759643277, 
    0.33645960505898209, 0.33415679014707672, 0.33188167691349979, 
    0.329634101990263, 0.32741389542737731, 0.325220879394018, 
    0.32305486477844603, 0.32091564583543986, 0.31880299568401715, 
    0.31671666414242605, 0.31465638134786628, 0.31262185823163458, 
    0.3106127906918783, 0.30862885894822095, 0.30666972853692798, 
    0.30473504892684555, 0.3028244477042491, 0.30093753111736066, 
    0.29907388229959675, 0.29723306201549665, 0.2954146082488861, 
    0.29361803637452066, 0.29184283735552768, 0.29008848011010679, 
    0.28835440617662411, 0.28664003131603483, 0.28494474206229803, 
    0.28326789433618393, 0.28160881053777892, 0.27996678034858052, 
    0.27834106338420811, 0.276730893489883, 0.27513548766043239, 
    0.27355405452228626, 0.27198581248174003, 0.27042999891515501, 
    0.26888588712036249, 0.26735279454057381, 0.26583009514349004, 
    0.26431722223161858, 0.26281367197160932, 0.26131900128943003, 
    0.25983282498516136, 0.25835480893726293, 0.25688466201223303, 
    0.25542212786886631, 0.25396697639858057, 0.25251899713505027, 
    0.25107799345817189, 0.24964378076497071, 0.24821618761407369, 
    0.24679505692380363, 0.24538024447521795, 0.24397161843104737, 
    0.24256905647098351, 0.24117244524937714, 0.23978167461056363, 
    0.23839663854575413, 0.23701723435937264, 0.23564336047338244, 
    0.23427491988526444, 0.23291182003755972, 0.23155397423768573, 
    0.23020130055588303, 0.22885372170513502, 0.22751115900334312, 
    0.22617353250734198, 0.22484075802933504, 0.22351274517257855, 
    0.22218939732917586, 0.22087061624060844, 0.21955630535670079, 
    0.21824637044650053, 0.21694072616962354, 0.21563930084370397, 
    0.21434203465438767, 0.21304888647299164, 0.21175982736872725, 
    0.21047484162970423, 0.2091939198723875, 0.20791706147607986, 
    0.20664426987159817, 0.20537555955893727, 0.20411095015433803, 
    0.20285047370856576, 0.20159417126473217, 0.20034209688912394, 
    0.19909431585572288, 0.19785090283421705, 0.19661194466587201, 
    0.19537753676166988, 0.19414778453919967, 0.19292280312228305, 
    0.1917027183923426, 0.19048767091089086, 0.18927781531296409, 
    0.1880733234214301, 0.18687438316122862, 0.18568119745407002, 
    0.18449397927700451, 0.18331294639819271, 0.18213831685384346, 
    0.18097029994058647, 0.17980909167285544, 0.1786548708333737, 
    0.17750779384584311, 0.17636799492708993, 0.17523558463887356, 
    0.17411064970304152, 0.17299325588699138, 0.17188344664695407, 
    0.17078124367100062, 0.1696866496504128, 0.16859964732097726, 
    0.16752019942466875, 0.16644824696312718, 0.16538370912222733, 
    0.16432648084963986, 0.16327642907137194, 0.16223339850387677, 
    0.1611972092688701, 0.16016766657395659, 0.15914456368059721, 
    0.15812769664868839, 0.15711686925006441, 0.15611190664301425, 
    0.15511265847977274, 0.15411900971874742, 0.15313088428668012, 
    0.15214824790492582, 0.15117110944231599, 0.15019951740094753, 
    0.14923355996313536, 0.14827336217185252, 0.14731908695994303, 
    0.1463709333314846, 0.1454291401520193, 0.14449398124455559, 
    0.143565764182773, 0.1426448231679282, 0.1417315130071482, 
    0.14082619656629047, 0.13992923188235387, 0.13904095946630196, 
    0.13816169169322753, 0.13729169479408729, 0.1364311853219142, 
    0.13558032124678854, 0.13473919964128445, 0.13390785800599081, 
    0.13308627700563674, 0.13227438873111808, 0.1314720863749948, 
    0.13067923186085195, 0.12989567009023126, 0.12912123940937764, 
    0.12835577870321002, 0.12759913441584117, 0.12685116610567157, 
    0.12611174603537942, 0.12538075886584374, 0.12465810136225677, 
    0.12394367854957503, 0.12323740285318882, 0.12253919265358, 
    0.12184897124759908, 0.1211666677276739, 0.1204922170572898, 
    0.11982556128198599, 0.11916665114480406, 0.11851544636510718, 
    0.11787191648679012, 0.11723603818809607, 0.11660779835589295, 
    0.11598719348875955, 0.11537423217108891, 0.1147689351042231, 
    0.1141713353129286, 0.11358147777709399, 0.11299941451893884, 
    0.11242520165249281, 0.11185889339511149, 0.11130053964333456, 
    0.11075017647767742, 0.1102078260966835, 0.10967349065781472, 
    0.10914714897280411, 0.10862875366781188, 0.10811823129961225, 
    0.10761548444500085, 0.10712039555050167, 0.10663283543771668, 
    0.10615267392042065, 0.10567978784562322, 0.10521407158875991, 
    0.10475544417170794, 0.1043038535459225, 0.10385927929407301, 
    0.10342173169095331, 0.1029912501469213, 0.10256789647336317, 
    0.10215175063070253, 0.10174290349809417, 0.10134144908242172, 
    0.10094747883379773, 0.10056107555968717, 0.10018231028156147, 
    0.099811236308527382, 0.099447889676756482, 0.099092285187462076, 
    0.09874441718162108, 0.098404259665343621, 0.098071766577030969, 
    0.097746872888794606, 0.097429495669385968, 0.097119533127152519, 
    0.096816866984173688, 0.096521361233413067, 0.096232863488492318, 
    0.095951205656701677, 0.095676204515618785, 0.095407662630371218, 
    0.095145371014501504, 0.094889105076852748, 0.094638628561940386, 
    0.094393686345324385, 0.094154002451396185, 0.093919272386733046, 
    0.093689156272923901, 0.093463276215640628, 0.093241215154642967, 
    0.093022512858802267, 0.092806668718641253, 0.092593143341920314, 
    0.092381359717972664, 0.092170704295953684, 0.091960534684861012, 
    0.091750186983218851, 0.091538987099806748, 0.091326265057248085, 
    0.091111363931343198, 0.090893653254109336, 0.090672541480063679, 
    0.090447488985678809, 0.090218020239392918, 0.089983732904634947, 
    0.089744306149132161, 0.089499503609946435, 0.089249171705110125, 
    0.088993237653952784, 0.088731699093393748, 0.088464620873999977, 
    0.088192122940382187, 0.087914375630106595, 0.087631591880042686, 
    0.087344020988628424, 0.08705194218647061, 0.086755660404030099, 
    0.086455497845938631, 0.08615178801007331, 0.085844872117541521, 
    0.085535090434161257, 0.085222780417175917, 0.084908273497928816, 
    0.084591894048157576, 0.084273962343650533, 0.083954791091479464, 
    0.083634691668385788, 0.083313972152793264, 0.082992935376890314, 
    0.082671876108917894, 0.08235107895130267, 0.082030816462379572, 
    0.081711352381879016, 0.081392942027744261, 0.081075837528319331, 
    0.080760287126931701, 0.080446537745004515, 0.080134837049953667, 
    0.079825432910253569, 0.079518574405022427, 0.079214508533519259, 
    0.07891347730130098, 0.078615709021171681, 0.078321410251458071, 
    0.07803075297889997, 0.077743868348696607, 0.077460834914876472, 
    0.077181673578968421, 0.076906342716339712, 0.076634735601284337, 
    0.076366680793679712, 0.076101948943244596, 0.07584025477166205, 
    0.075581268096722068, 0.075324621221814478, 0.075069916603208553, 
    0.0748167392224445, 0.074564664300619754, 0.074313270966901421, 
    0.074062150863131476, 0.073810916347456818, 0.073559210354515278, 
    0.073306713250837374, 0.073053148681554519, 0.07279829028897411, 
    0.072541966365425564, 0.072284064722353436, 0.072024539688720066, 
    0.071763413948156898, 0.071500782691676909, 0.071236809116432778, 
    0.070971721164239179, 0.070705804258983873, 0.070439389987878617, 
    0.070172841181596682, 0.069906542595185292, 0.06964088492440372, 
    0.06937625036619538, 0.069112998096396649, 0.068851449586420685, 
    0.068591874086490243, 0.068334478160817724, 0.068079391848582749, 
    0.067826659687535817, 0.067576236030158152, 0.067327976897668881, 
    0.067081642751919635, 0.066836898674288089, 0.066593325922327709, 
    0.066350436322312772, 0.066107690187416954, 0.065864518259821342, 
    0.065620340068070465, 0.065374579583389575, 0.06512667932253699, 
    0.064876106961957683, 0.064622365419064423, 0.064364997272249438, 
    0.064103590909144997, 0.063837784651423493, 0.063567272464788188, 
    0.063291806851389909, 0.063011208564196425, 0.062725369788435903, 
    0.062434261288349578, 0.06213793368761044, 0.061836515416432751, 
    0.061530212783408179, 0.061219301830384834, 0.06090412353776694, 
    0.060585073134503592, 0.060262594697635598, 0.059937173997626395, 
    0.059609330851359263, 0.059279616381860238, 0.058948607445915978, 
    0.058616906450286485, 0.058285132543835515, 0.057953923277236252, 
    0.057623924595522541, 0.05729578913525403, 0.056970169498319005, 
    0.056647713233035538, 0.056329053436965752, 0.056014801535384032, 
    0.055705536838083325, 0.055401796537357356, 0.055104064434731433, 
    0.054812758425583044, 0.054528225377130812, 0.054250731476020858, 
    0.053980457599894477, 0.053717502898336267, 0.05346188757345291, 
    0.053213557652535749, 0.052972392769793188, 0.05273820907480594, 
    0.052510761328153313, 0.05228974363716999, 0.052074791567378174, 
    0.05186548380351666, 0.051661343685790159, 0.051461845245946637, 
    0.051266420185798064, 0.051074469005883444, 0.050885376144964009, 
    0.050698523552962706, 0.050513308507142786, 0.050329155715405131, 
    0.050145530830628463, 0.049961947802402984, 0.049777975717182371, 
    0.049593244142153478, 0.049407442805804593, 0.049220318617184712, 
    0.049031673647417548, 0.048841360844668946, 0.048649278167672727, 
    0.048455365773444933, 0.048259601018743374, 0.04806199731004946, 
    0.0478626006469694, 0.047661490515031629, 0.047458776526549777, 
    0.047254597007943787, 0.047049115378017418, 0.046842512975429899, 
    0.046634987125301876, 0.046426744390658643, 0.04621800048035387, 
    0.046008978089933997, 0.045799908852088594, 0.045591030826375577, 
    0.045382590404273594, 0.045174836069430784, 0.04496802301644065, 
    0.044762406900933221, 0.044558247639180461, 0.04435581098953717, 
    0.044155372424044624, 0.043957218072348245, 0.043761651563697754, 
    0.043568991530989351, 0.043379571766262982, 0.043193738418961014, 
    0.043011843020134256, 0.042834236946969438, 0.042661261258934241, 
    0.042493238282591189, 0.042330458360241505, 0.042173167392070228, 
    0.042021558962439517, 0.041875760817404684, 0.041735830186763717, 
    0.041601749684854042, 0.041473425547929259, 0.041350693827750321, 
    0.041233324569547931, 0.041121033268875548, 0.041013485442969372, 
    0.040910307279288682, 0.040811088875147242, 0.040715395726331517, 
    0.040622772668714516, 0.040532757279628948, 0.040444887092955586, 
    0.040358713735827841, 0.040273809798263491, 0.040189777653376203, 
    0.040106252739320711, 0.040022907736877389, 0.039939454596795453, 
    0.039855643977491244, 0.039771263717437985, 0.039686136626389514, 
    0.039600120207853459, 0.039513099016286399, 0.039424984189463969, 
    0.039335708125476404, 0.039245221849598347, 0.039153495457241019, 
    0.039060515030603732, 0.038966282327595664, 0.038870813580760583, 
    0.038774139074206009, 0.038676298205363918, 0.038577337440047182, 
    0.038477305141973839, 0.038376248880579888, 0.038274214092115878, 
    0.038171238408602162, 0.038067351049539552, 0.037962571018094166, 
    0.037856903575292325, 0.037750344654041285, 0.037642878072471762, 
    0.037534479853851652, 0.037425120205426911, 0.037314764886212333, 
    0.03720338068052674, 0.037090935419097401, 0.03697739982147151, 
    0.036862750465923549, 0.036746971000110339, 0.03663005477676981, 
    0.036512007166201156, 0.036392846136306105, 0.036272608545267503, 
    0.036151343324377708, 0.036029119157382085, 0.035906018393535279, 
    0.035782133332833886, 0.03565756344662431, 0.035532411247840553, 
    0.035406776530434794, 0.03528075470849007, 0.035154431386575404, 
    0.035027881637079296, 0.034901163963035879, 0.03477431968479909, 
    0.034647365675068778, 0.034520290066428747, 0.034393045044973973, 
    0.034265538994724912, 0.03413763369553377, 0.034009142464856479, 
    0.03387982904121041, 0.033749412447309127, 0.033617573697832047, 
    0.033483960116663533, 0.033348194405155837, 0.033209886831248946, 
    0.033068643330664463, 0.032924079266071271, 0.032775829473221982, 
    0.032623562290490259, 0.032466986892000504, 0.032305864762525387, 
    0.032140016482526089, 0.031969327438903142, 0.03179375399516491, 
    0.031613325686135757, 0.031428146260554179, 0.031238393120709987, 
    0.031044313905020542, 0.030846220397779449, 0.030644480238977846, 
    0.030439507331741018, 0.030231752089969678, 0.030021686587961775, 
    0.029809796343771316, 0.029596567471923504, 0.029382477520823166, 
    0.029167989087041778, 0.028953542278324449, 0.028739546732821749, 
    0.028526375818938556, 0.028314358646317796, 0.028103769338593734, 
    0.027894819493130791, 0.027687653717989598, 0.027482354691034598, 
    0.027278950366588312, 0.027077425625647304, 0.026877736697864793, 
    0.026679823795048345, 0.026483623627072298, 0.026289077816544364, 
    0.026096139091611018, 0.025904777858577067, 0.025714976121922944, 
    0.025526724450780303, 0.025340013021996063, 0.025154822977493232, 
    0.02497111194148072, 0.02478880844367955, 0.02460780444039895, 
    0.02442794509165494, 0.024249024422993769, 0.024070778671954361, 
    0.023892885444129163, 0.023714960866259269, 0.023536564063721781, 
    0.023357211734494544, 0.023176394818717916, 0.022993605824449419, 
    0.022808365154579343, 0.022620249899544018, 0.022428916735707023, 
    0.022234123350636625, 0.022035742750550407, 0.021833765119962892, 
    0.021628290874950447, 0.021419511533972761, 0.021207684299795495, 
    0.020993110816269662, 0.020776114538922218, 0.020557032695506829, 
    0.020336206228535436, 0.020113972873726405, 0.019890661673174059, 
    0.019666586684070023, 0.019442040044747564, 0.019217286427408893, 
    0.018992561520231932, 0.018768067152894599, 0.018543973877989978, 
    0.018320420405798985, 0.018097518629090491, 0.017875357071209699, 
    0.017654002245001139, 0.017433508476003237, 0.017213913277822533, 
    0.016995245720362387, 0.016777525111978882, 0.01656076180778264, 
    0.016344953832138111, 0.016130089189827754, 0.015916141818459052, 
    0.015703072270676629, 0.015490828160126284, 0.015279350866202739, 
    0.015068579667897423, 0.014858463932660385, 0.014648974322276746, 
    0.014440107246551171, 0.014231890315347943, 0.01402438348125771, 
    0.013817669744791875, 0.013611849349835878, 0.013407028742960073, 
    0.013203314597691806, 0.013000804478712718, 0.012799583593276624, 
    0.012599721506529011, 0.012401271958734894, 0.012204272877892153, 
    0.012008748979692171, 0.011814714038892483, 0.011622173385084349, 
    0.011431122967714565, 0.011241550139616578, 0.011053429874432807, 
    0.010866722407473713, 0.010681370326278555, 0.010497297661125848, 
    0.010314408188000031, 0.010132587467865996, 0.0099517016406421785, 
    0.0097715975762472044, 0.0095921040342001641, 0.0094130267476584678, 
    0.0092341566458529929, 0.0090552658520332962, 0.0088761162433512852, 
    0.0086964607345300475, 0.008516047842030406, 0.0083346280690361953, 
    0.0081519557848122939, 0.0079677938701463377, 0.0077819165880945781, 
    0.0075941131935521999, 0.0074041896806609523, 0.0072119734532777261, 
    0.0070173147851126435, 0.0068200868055178325, 0.006620190464220391, 
    0.0064175527753414308, 0.0062121271937172623, 0.0060038978692251201, 
    0.0057928791025329517, 0.0055791177854675935, 0.0053626984880713272, 
    0.0051437399934921579, 0.0049224045222939234, 0.0046988938275676637, 
    0.0044734503349815151, 0.0042463535890776534, 0.0040179153636331153, 
    0.0037884767143404607, 0.0035583963453529139, 0.0033280475857548966, 
    0.0030978064148977245, 0.0028680466428809884, 0.002639131151233225, 
    0.0024114006640590466, 0.002185170701088964, 0.0019607257740498242, 
    0.0017383176465871975, 0.0015181625980455078, 0.001300447477394913, 
    0.0010853324483613227, 0.00087295660837593387, 0.00066344140505475652, 
    0.00045689658421252171, 0.00025341631551211016, 5.3078830168514684e-05, 
    -0.00014405586653577535, -0.00033794896267226766, 
    -0.00052858760241964852, -0.00071598336433597817, 
    -0.00090017437223532774, -0.0010812229300608141, -0.0012592183248931544, 
    -0.0014342757134558435, -0.0016065367157151631, -0.0017761709538874487, 
    -0.0019433777815201978, -0.0021083891235790918, -0.0022714682616241954, 
    -0.0024329115247111784, -0.0025930447889673689, -0.0027522238932590542, 
    -0.0029108260814318596, -0.0030692483104120794, -0.0032279008319696465, 
    -0.0033872014802229025, -0.0035475646299782922, -0.0037093945989285799, 
    -0.0038730697533397454, -0.0040389328191240779, -0.0042072752716122647, 
    -0.004378326577709769, -0.0045522484376690313, -0.0047291330390560413, 
    -0.0049090064916011257, -0.0050918325838063827, -0.0052775270219043869, 
    -0.0054659616050754612, -0.0056569789479686801, -0.005850397458893466, 
    -0.0060460194994705905, -0.0062436371617568135, -0.0064430341889329407, 
    -0.0066439887311504856, -0.0068462739043197059, -0.0070496641953724289, 
    -0.0072539366493271388, -0.0074588739634936707, -0.0076642718121912746, 
    -0.0078699394681738845, -0.0080757078361893084, -0.0082814287245189366, 
    -0.0084869818489540314, -0.0086922755335598536, -0.008897249933701442, 
    -0.0091018784031399701, -0.0093061684975982752, -0.0095101605652120873, 
    -0.0097139295240672944, -0.0099175783273309712, -0.010121234095780383, 
    -0.010325037785540527, -0.010529136358703759, -0.010733669205533765, 
    -0.010938761129069684, -0.011144510890006856, -0.011350983614539699, 
    -0.011558205674885884, -0.011766158238694089, -0.011974780224300907, 
    -0.012183962519115653, -0.012393557188260507, -0.012603378696139412, 
    -0.01281321079482076, -0.013022817610367039, -0.013231948367324803, 
    -0.013440350771942408, -0.013647776693025981, -0.013853989809079138, 
    -0.014058772146429512, -0.014261929299214073, -0.014463290385407553, 
    -0.01466270917576671, -0.014860065308943654, -0.015055261467717877, 
    -0.015248220216247136, -0.015438881400466746, -0.01562719697901541, 
    -0.01581312500310043, -0.015996620346017551, -0.016177627085903052, 
    -0.016356069699419284, -0.016531841757958177, -0.016704799250997496, 
    -0.016874754798982324, -0.017041472286913634, -0.017204668253763794, 
    -0.017364012079081555, -0.01751913401457228, -0.017669631973585422, 
    -0.017815080866144969, -0.017955044534069663, -0.018089084273430461, 
    -0.018216769712885932, -0.018337688138583524, -0.018451449628366305, 
    -0.01855769484893276, -0.018656100911829676, -0.018746383257551194, 
    -0.018828302044619646, -0.018901660990102341, -0.018966309991215784, 
    -0.019022142788972428, -0.019069095964078138, -0.01910714766135032, 
    -0.019136316504297025, -0.019156658307947095, -0.019168270316068894, 
    -0.019171292835942058, -0.019165911224279519, -0.019152352692103945, 
    -0.019130885294390887, -0.019101811738826253, -0.0190654660181463, 
    -0.019022206631521231, -0.01897241577376033, -0.018916494818634173, 
    -0.018854861533230346, -0.018787946225890056, -0.018716187603428181, 
    -0.018640028902083727, -0.018559912503650269, -0.018476278943434267, 
    -0.018389561435172889, -0.018300185661752798, -0.018208569287995382, 
    -0.018115121376047823, -0.018020238580158117, -0.017924308186873496, 
    -0.017827706799245901, -0.017730795117700725, -0.017633916651118554, 
    -0.01753739346966136, -0.017441521140807749, -0.017346562430762311, 
    -0.0172527456525382, -0.01716026219184363, -0.017069263899640533, 
    -0.016979869944236843, -0.016892165736407661, -0.016806206029225997, 
    -0.016722021293846763, -0.016639613035870603, -0.016558961075162131, 
    -0.016480024608433085, -0.016402747044465201, -0.016327059508720581, 
    -0.01625288427940003, -0.016180137207136056, -0.016108731453911035, 
    -0.016038574716095846, -0.015969570916481012, -0.015901620960992971, 
    -0.015834621768680581, -0.015768466918947736, -0.015703047631645092, 
    -0.01563825748478101, -0.015573994239651456, -0.015510163163357019, 
    -0.015446682218549628, -0.015383485740690385, -0.015320528870491007, 
    -0.015257789426328872, -0.015195268660803679, -0.015132993979371498, 
    -0.015071016118876093, -0.015009408681659618, -0.014948266949441843, 
    -0.01488770107914773, -0.014827835379889428, -0.014768802263947575, 
    -0.014710738559433261, -0.014653781846655757, -0.014598066539070394, 
    -0.014543721044503031, -0.014490863722372533, -0.014439596386541747, 
    -0.014390003757232464, -0.014342145009442225, -0.014296052960570529, 
    -0.014251728700136804, -0.014209142570466007, -0.014168234353271428, 
    -0.014128914894549077, -0.014091074134449908, -0.014054586523213208, 
    -0.014019318792506589, -0.01398514126612287, -0.013951931056400104, 
    -0.01391958410744833, -0.013888019228191639, -0.013857181377529813, 
    -0.013827043808498894, -0.013797607165200211, -0.01376889659597068, 
    -0.013740957253750631, -0.01371385273841615, -0.013687657433256556, 
    -0.013662457885587211, -0.013638347059496379, -0.013615422123748449, 
    -0.013593782309879799, -0.013573521867982908, -0.013554727482569331, 
    -0.01353747292885998, -0.013521814351657901, -0.01350778898634877, 
    -0.013495414891096293, -0.013484696343676298, -0.013475636793364321, 
    -0.013468246684062856, -0.01346256149285683, -0.013458653395546367, 
    -0.01345664321998831, -0.013456709096445824, -0.01345908576378194, 
    -0.013464064958130417, -0.013471984208962454, -0.013483215269413987, 
    -0.013498150791366037, -0.013517189134170462, -0.013540721085370728, 
    -0.013569120266412823, -0.013602736032014721, -0.0136418916623891, 
    -0.013686880402326506, -0.013737965300539594, -0.01379538073774546, 
    -0.013859327041648059, -0.013929967929942748, -0.014007423663936465, 
    -0.014091765313048676, -0.014183003887979367, -0.014281082015142351, 
    -0.014385868029207351, -0.014497150146364969, -0.014614634370366236, 
    -0.014737947427367983, -0.014866641562797656, -0.015000197410074721, 
    -0.015138035056011136, -0.015279517027789166, -0.015423960473246514, 
    -0.015570645929143822, -0.015718831889200938, -0.015867768982435956, 
    -0.016016714441611044, -0.016164951328650527, -0.016311804653867747, 
    -0.01645665531287982, -0.016598951879948913, -0.01673822403204471, 
    -0.016874087922750972, -0.017006252539403497, -0.017134519434811511, 
    -0.017258775184544963, -0.017378987360729917, -0.017495189934011546, 
    -0.017607472959727678, -0.017715972281333984, -0.017820861747958945, 
    -0.017922349988766517, -0.0180206742566551, -0.018116098394874675, 
    -0.018208905699564754, -0.018299389884223506, -0.018387845659866186, 
    -0.018474556377242046, -0.018559781023316103, -0.018643744269072771, 
    -0.018726625452559265, -0.018808551528346464, -0.018889591526444316, 
    -0.018969752216304734, -0.019048979258464181, -0.019127159217773314, 
    -0.019204126824621286, -0.019279669334546692, -0.019353539285028119, 
    -0.019425460004045408, -0.019495133436119819, -0.019562249004104221, 
    -0.019626486924890947, -0.019687522015403719, -0.019745029338970835, 
    -0.019798687759164883, -0.019848185879038006, -0.01989322887239214, 
    -0.019933548062088108, -0.01996890381738553, -0.019999099657640389, 
    -0.020023981937763183, -0.020043448032334751, -0.02005744633259627, 
    -0.020065974219438121, -0.020069078343834552, -0.020066847841992749, 
    -0.020059414437917679, -0.020046946806940191, -0.020029646232606099, 
    -0.020007739151656486, -0.019981473733119787, -0.019951108894041655, 
    -0.019916908192745768, -0.019879130470283075, -0.019838024630444043, 
    -0.019793821884191397, -0.019746731196088413, -0.019696935301161865, 
    -0.019644586453490334, -0.019589804480744478, -0.019532674497108889, 
    -0.01947324668244586, -0.01941153566039365, -0.01934751915760893, 
    -0.019281140914281718, -0.019212312934723912, -0.01914092199568828, 
    -0.019066833903811496, -0.018989900513682004, -0.018909967674766839, 
    -0.018826882741813652, -0.018740501488426747, -0.01865069593637016, 
    -0.018557358443511557, -0.01846040753891328, -0.018359791931396512, 
    -0.018255493998871559, -0.018147529906387825, -0.018035953006021802, 
    -0.0179208511145433, -0.017802346345664511, -0.017680589515556865, 
    -0.017555758841202845, -0.017428050347022012, -0.01729767433437851, 
    -0.017164847726466991, -0.017029789146580977, -0.016892713872113253, 
    -0.016753831358956809, -0.01661334285396282, -0.016471442058379412, 
    -0.016328316939188636, -0.016184150370799361, -0.016039125886218471, 
    -0.0158934294377523, -0.01574725232423952, -0.015600793707210379, 
    -0.015454261419343395, -0.015307872329290208, -0.015161851653858333, 
    -0.01501643074281216, -0.014871846657475662, -0.014728340575145767, 
    -0.014586157039580378, -0.014445541754402963, -0.014306741258799327, 
    -0.014170001920191168, -0.014035571589709585, -0.013903697367833718, 
    -0.013774629268931377, -0.013648616583853345, -0.013525909611638857, 
    -0.013406759113597223, -0.013291408735363389, -0.013180090247488395, 
    -0.013073021123553063, -0.012970391649210062, -0.012872362276268371, 
    -0.012779057762499086, -0.012690563869882224, -0.012606928219709782, 
    -0.012528156172837181, -0.012454215892903336, -0.012385029689901683, 
    -0.012320477258679994, -0.012260393101890886, -0.012204559039156496, 
    -0.012152708245059275, -0.012104522274807222, -0.012059635419416338, 
    -0.012017641444739586, -0.011978100820794358, -0.01194055542236858, 
    -0.01190453748095097, -0.01186958522238205, -0.011835250602916588, 
    -0.011801111379189174, -0.01176677435943631, -0.011731881935584177, 
    -0.011696110217159631, -0.011659168363251243, -0.011620793495069427, 
    -0.011580747542170663, -0.011538811149808972, -0.011494781124525398, 
    -0.011448466975926936, -0.011399692317152151, -0.01134829649589564, 
    -0.011294142750291357, -0.011237125116189111, -0.011177179152271649, 
    -0.011114289236775285, -0.011048495204056877, -0.010979895106732458, 
    -0.010908643675563474, -0.010834947668005168, -0.010759056899646636, 
    -0.010681251963956737, -0.010601832033418504, -0.010521105526014631, 
    -0.010439373834677801, -0.010356922356372441, -0.010274014231372855, 
    -0.010190878818709365, -0.010107712328299942, -0.010024671712680108, 
    -0.0099418757439352703, -0.0098594043626708747, -0.0097772998308753543, 
    -0.0096955653246318021, -0.009614168577227732, -0.0095330394293807932, 
    -0.0094520743076572621, -0.0093711360571428343, -0.0092900609323660031, 
    -0.0092086618815495312, -0.0091267349466690236, -0.0090440608008825023, 
    -0.008960416278124406, -0.0088755751683295397, -0.0087893139707439193, 
    -0.0087014211722813914, -0.008611698214603657, -0.0085199676105720684, 
    -0.0084260721489706116, -0.0083298771928989688, -0.0082312681291689463, 
    -0.0081301487821686946, -0.008026440106563365, -0.0079200782123848984, 
    -0.0078110128522567131, -0.0076992055750061527, -0.0075846257500702336, 
    -0.0074672439385975115, -0.0073470315854476552, -0.0072239521776964457, 
    -0.0070979647895876852, -0.006969023972963821, -0.0068370924293588622, 
    -0.006702152334881771, -0.0065642154161859156, -0.0064233393364441227, 
    -0.0062796298437913477, -0.0061332520242504528, -0.0059844328985925298, 
    -0.0058334659386358864, -0.0056807052687515448, -0.0055265639937068988, 
    -0.0053715026625008357, -0.0052160190766131617, -0.0050606311131931227, 
    -0.0049058680805471686, -0.0047522619860123558, -0.0046003386500073776, 
    -0.004450613023390634, -0.0043035805748234063, -0.0041597138307322085, 
    -0.0040194592977208666, -0.003883230739451534, -0.0037514128539474839, 
    -0.003624356354040867, -0.0035023848011705968, -0.0033857981346577205, 
    -0.0032748787266012025, -0.0031698974913649787, -0.0030711266625961997, 
    -0.0029788460376112312, -0.0028933520524807967, -0.0028149596879533147, 
    -0.0027439984280719339, -0.0026808048494848975, -0.0026257103212800437, 
    -0.0025790273357848732, -0.0025410380088459993, -0.0025119852386626439, 
    -0.0024920660368759591, -0.0024814305399441178, -0.002480180159262651, 
    -0.0024883668748364104, -0.0025059919360752173, -0.0025330088172131207, 
    -0.002569319067805719, -0.0026147752044585778, -0.0026691733701825794, 
    -0.0027322520208945956, -0.0028036907581961167, -0.0028831020372718443, 
    -0.0029700319803819893, -0.0030639548050440018, -0.0031642724136839496, 
    -0.0032703135065470655, -0.003381334432401096, -0.0034965254328092892, 
    -0.0036150155779932423, -0.003735883843792392, -0.0038581724389337583, 
    -0.0039809000114956654, -0.0041030773372467567, -0.004223723033147676, 
    -0.0043418764974675599, -0.0044566097418953709, -0.0045670369159139124, 
    -0.0046723231602999833, -0.0047716870649789416, -0.00486441339581068, 
    -0.004949854405173643, -0.0050274410364789489, -0.0050966884088569555, 
    -0.0051572013340760725, -0.0052086723227867055, -0.0052508795644321477, 
    -0.0052836814656528818, -0.0053070081495086513, -0.0053208526533039275, 
    -0.00532526245089313, -0.005320330547021899, -0.0053061939931620412, 
    -0.0052830225651740231, -0.0052510150271469084, -0.005210395256669045, 
    -0.0051613977343549717, -0.0051042614150469271, -0.0050392175027023913, 
    -0.0049664852930332995, -0.0048862582350681655, -0.004798704463637663, 
    -0.0047039612625393327, -0.0046021342664308573, -0.0044933034862865307, 
    -0.00437753099591154, -0.0042548624609658756, -0.0041253384644862699, 
    -0.0039890020746410331, -0.0038458983269322317, -0.0036960767434079935, 
    -0.0035395896692124069, -0.0033764939975644125, -0.0032068463758620925, 
    -0.0030307073399557997, -0.0028481394188217082, -0.0026592177227096154, 
    -0.0024640320217883815, -0.0022626958195506837, -0.002055356167337344, 
    -0.0018421980616877415, -0.0016234442548290907, -0.0013993581594425979, 
    -0.0011702369185051889, -0.00093640470458584068, -0.00069820857245380297, 
    -0.00045601038610489238, -0.00021018507474514182, 3.8879241265903867e-05, 
    0.00029078207074026007, 0.00054510925228533585, 0.00080142488265237135, 
    0.0010592706386264791, 0.0013181569556724171, 0.0015775614816125247, 
    0.0018369274992795007, 0.0020956598675593557, 0.0023531379836588756, 
    0.0026087165227453371, 0.0028617365650741057, 0.0031115285402660894, 
    0.0033574208921107896, 0.0035987397731730422, 0.0038348196075376302, 
    0.0040650103382114623, 0.0042886830400977868, 0.0045052438108096164, 
    0.0047141470397461518, 0.0049149052903303056, 0.00510709935038878, 
    0.0052903893151055982, 0.0054645139824734713, 0.0056292979187557383, 
    0.0057846448355862159, 0.0059305307491519244, 0.0060669940833098079, 
    0.0061941285799965865, 0.0063120661220857702, 0.006420971038643225, 
    0.0065210351450730852, 0.0066124695949232488, 0.0066955091186076529, 
    0.0067704125858021732, 0.0068374726391828584, 0.0068970156605134766, 
    0.0069494119731885609, 0.0069950775413850164, 0.0070344729048735961, 
    0.0070680963987357712, 0.0070964771990354716, 0.0071201652221583719, 
    0.007139719626335389, 0.0071557003144240901, 0.007168664714600894, 
    0.0071791646487148943, 0.0071877444295024764, 0.00719494043543024, 
    0.0072012860728649635, 0.0072073136079346366, 0.0072135600599814841, 
    0.0072205681023999949, 0.0072288925460938522, 0.0072391038978967667, 
    0.0072517851250278363, 0.0072675280211241065, 0.0072869277902569991, 
    0.007310570961619074, 0.007339019412954919, 0.0073727931153820814, 
    0.0074123574271223206, 0.0074581081035434036, 0.0075103608282925949, 
    0.0075693461621385016, 0.0076352059787654965, 0.0077079960754531697, 
    0.0077876976834300804, 0.0078742221955521198, 0.0079674251221157257, 
    0.0080671214624112898, 0.0081730985001658412, 0.0082851316109806943, 
    0.0084029997442485113, 0.008526505825782054, 0.0086554905229758537, 
    0.0087898474901707043, 0.0089295317321164761, 0.0090745589282704223, 
    0.0092249950486167458, 0.009380935924555937, 0.0095424886396271603, 
    0.009709752791878903, 0.0098828115048098554, 0.010061719443975697, 
    0.010246502485281073, 0.010437156390038031, 0.010633642392903583, 
    0.010835889645644709, 0.01104378866631889, 0.011257190690652985, 
    0.011475901565170471, 0.011699679087770646, 0.011928226025725894, 
    0.012161191784256415, 0.01239816850367464, 0.01263869342186119, 
    0.01288225517649484, 0.013128304698372794, 0.013376259457069304, 
    0.013625518452543089, 0.01387547222809851, 0.014125508765535109, 
    0.014375019592486396, 0.014623403671237004, 0.014870066600837253, 
    0.015114420505379648, 0.01535588014683412, 0.015593867757457941, 
    0.015827815141141302, 0.016057169735528402, 0.016281402269177039, 
    0.016500009721251305, 0.016712528977883757, 0.016918534978004669, 
    0.017117661698438768, 0.017309608599407153, 0.01749415139988892, 
    0.017671144769943675, 0.017840527375971506, 0.018002324973313041, 
    0.01815664945818965, 0.018303699708634446, 0.018443756093653563, 
    0.018577173391167288, 0.018704374548739838, 0.018825829820303789, 
    0.018942047844668387, 0.019053551390402074, 0.019160860515908408, 
    0.019264477386929085, 0.019364863174047543, 0.019462434310652827, 
    0.01955755724290037, 0.019650540906471118, 0.019741645358268441, 
    0.019831072730243007, 0.019918966023870797, 0.020005404052420322, 
    0.020090396484125583, 0.020173886204506428, 0.020255749135996943, 
    0.020335807173108837, 0.02041383906210938, 0.020489600889818955, 
    0.020562843724386631, 0.020633328804553167, 0.02070084015016135, 
    0.020765195797932293, 0.020826255099264078, 0.020883922935671088, 
    0.020938153569406426, 0.020988952646552782, 0.021036374576942681, 
    0.021080526286404212, 0.021121560438258451, 0.02115967134380025, 
    0.021195081627254791, 0.021228033039914388, 0.021258763960928181, 
    0.021287495439507718, 0.021314402976326301, 0.021339609611959579, 
    0.021363159780047637, 0.021385008351949449, 0.021405007674073707, 
    0.021422908459672308, 0.021438360976628022, 0.021450917441992193, 
    0.02146004609207593, 0.021465145227157097, 0.021465564242509196, 
    0.021460625942154237, 0.021449640159778315, 0.021431935705607835, 
    0.021406873930711969, 0.02137386857912385, 0.021332395756145862, 
    0.021282000426965767, 0.021222304122466101, 0.021153001166960856, 
    0.021073852576544826, 0.020984680179663911, 0.020885357169119323, 
    0.020775808593438628, 0.020656012961262103, 0.020526020076261909, 
    0.020385967599694962, 0.020236100760955378, 0.020076785763137681, 
    0.019908510174360104, 0.019731877915623936, 0.019547590441853401, 
    0.019356435014306141, 0.019159259333144846, 0.018956954353211427, 
    0.018750425285205763, 0.018540574554764103, 0.018328286171805, 
    0.018114405754777019, 0.017899732315100416, 0.017685013821519741, 
    0.017470948467220561, 0.017258178147321977, 0.017047291998916029, 
    0.016838811390862674, 0.016633187367871061, 0.016430784768972258, 
    0.016231875666851654, 0.01603663202349492, 0.015845125198133858, 
    0.015657330966413412, 0.015473139505847968, 0.015292376946692658, 
    0.015114824493562726, 0.01494024175144871, 0.014768388559768626, 
    0.014599044062974903, 0.014432018423125217, 0.014267160175226485, 
    0.014104361985188323, 0.013943559202618031, 0.013784723181450225, 
    0.013627862779483243, 0.01347302634556702, 0.013320300055454579, 
    0.01316981423094526, 0.013021744178311267, 0.012876309539268226, 
    0.012733766855346929, 0.012594402695714978, 0.012458520404296184, 
    0.012326424274635431, 0.012198407443921123, 0.012074733884452488, 
    0.011955632513411968, 0.011841282267369834, 0.011731817907201975, 
    0.011627325313965136, 0.011527845664105755, 0.011433380881626423, 
    0.011343901801036322, 0.011259354084553917, 0.011179673693775911, 
    0.0111047861171449, 0.011034615819160576, 0.010969064258450624, 
    0.010907987209854125, 0.010851166975416382, 0.010798295479768339, 
    0.010748964854557242, 0.010702680562633579, 0.010658871147721686, 
    0.010616902440265653, 0.010576095401328171, 0.01053573639310885, 
    0.010495097805393374, 0.01045345052628876, 0.010410082711096761, 
    0.010364311758845089, 0.010315489599960394, 0.010263009292887221, 
    0.01020630213691171, 0.010144831943838695, 0.010078088443622426, 
    0.010005592155341409, 0.0099268864996150258, 0.0098415483924606771, 
    0.0097491907422015515, 0.0096494803938356761, 0.0095421546011845836, 
    0.0094270304992987858, 0.0093040188801080236, 0.0091731344657418855, 
    0.0090344972384846772, 0.0088883411888155909, 0.0087350102175204978, 
    0.0085749654175909969, 0.0084087807154331218, 0.0082371443650141613, 
    0.0080608484635742855, 0.0078807717859913015, 0.0076978489785397676, 
    0.0075130418878599876, 0.0073273097555341601, 0.0071415895982051532, 
    0.006956790212320707, 0.00677379196748862, 0.0065934512838067335, 
    0.0064166034425955226, 0.0062440650960681032, 0.0060766339242184289, 
    0.0059150855840261647, 0.0057601615895681805, 0.0056125648686458224, 
    0.0054729460239442071, 0.0053418910979270116, 0.0052199166429057892, 
    0.0051074696206240876, 0.0050049177260572701, 0.0049125591148549384, 
    0.004830623594873816, 0.0047592801703893331, 0.0046986424618429652, 
    0.004648772260855613, 0.0046096944601046602, 0.0045813886198336788, 
    0.0045637942250709388, 0.0045568172480578793, 0.0045603259806715618, 
    0.0045741594198497239, 0.0045981273703573043, 0.0046320178058360294, 
    0.0046755955273369192, 0.004728609076649474, 0.0047907870435154832, 
    0.0048618395397698336, 0.0049414615565911268, 0.0050293325682317681, 
    0.0051251200936389268, 0.005228493398883852, 0.0053391158388296093, 
    0.0054566645072182413, 0.0055808249213760023, 0.0057113132734966368, 
    0.0058478750872240906, 0.0059903054567333009, 0.006138457651555438, 
    0.0062922447756882452, 0.0064516377282499999, 0.0066166504375430686, 
    0.0067873355513524934, 0.0069637622580637284, 0.0071459876444674086, 
    0.0073340498750187715, 0.00752793296002305, 0.0077275505147843598, 
    0.0079327364602035447, 0.008143234778658727, 0.0083586926596653614, 
    0.0085786644441626092, 0.0088026126919309861, 0.0090299187683989864, 
    0.0092598848342390887, 0.0094917560468888527, 0.0097247266872241365, 
    0.0099579658502936767, 0.010190635180186019, 0.010421925333657791, 
    0.010651073747761301, 0.010877395349834696, 0.011100294114629776, 
    0.011319286005568599, 0.011534001102667526, 0.011744192568778336, 
    0.011949741012305989, 0.012150666520436898, 0.012347120977003993, 
    0.012539400751088468, 0.012727931569166153, 0.012913263899182565, 
    0.013096060879758262, 0.01327707707279142, 0.013457152345745092, 
    0.013637187936807564, 0.013818147122141163, 0.01400101995161155, 
    0.014186841710554168, 0.014376666245165214, 0.014571553378076462, 
    0.014772567666491725, 0.014980772408038015, 0.015197217406376223, 
    0.015422938565195372, 0.015658945018639042, 0.015906215088598335, 
    0.016165673610408268, 0.016438174186476993, 0.016724480544266153, 
    0.01702523506554968, 0.017340950765102132, 0.017671982507961162, 
    0.018018516872867239, 0.018380552689211471, 0.018757905011621466, 
    0.019150180101401536, 0.019556765848403629, 0.019976825311419776, 
    0.020409298268652905, 0.020852895358768057, 0.02130611090067238, 
    0.021767238478583112, 0.022234406995331212, 0.022705603178874462, 
    0.023178713322950194, 0.023651556899103789, 0.024121913085280684, 
    0.02458755461633368, 0.02504626992871203, 0.025495878445460141, 
    0.025934245746811919, 0.026359298165682079, 0.026769042712050346, 
    0.027161560939848329, 0.027535025798165018, 0.027887707082094031, 
    0.02821798620896368, 0.02852436099387156, 0.028805456025625092, 
    0.029060044222524777, 0.029287054961884978, 0.029485593187530076, 
    0.02965495910805897, 0.029794663660673192, 0.029904442078738873, 
    0.029984267229996624, 0.030034357181997096, 0.030055161985143512, 
    0.030047360761729383, 0.030011839411325517, 0.029949664132006972, 
    0.029862038754697721, 0.029750277465530814, 0.029615776692337063, 
    0.029459984241863059, 0.029284386916923415, 0.029090488169940525, 
    0.028879809307504879, 0.028653883293340832, 0.028414237023549494, 
    0.028162397774383563, 0.027899880564998713, 0.027628187491874182, 
    0.027348800814688073, 0.027063188612593679, 0.026772794039499254, 
    0.026479031524399239, 0.026183273182076097, 0.025886841433692694, 
    0.025590984827753599, 0.02529686503588361, 0.025005530230870605, 
    0.024717904357531122, 0.024434747422422208, 0.024156630409555981, 
    0.023883906210803475, 0.023616686678143595, 0.023354840170018612, 
    0.023097972387031422, 0.02284545549694323, 0.022596444995619303, 
    0.02234991760605028, 0.022104721263748527, 0.021859623140054733, 
    0.02161336569748535, 0.021364730023643898, 0.021112563421068337, 
    0.020855832479676591, 0.020593637601013993, 0.020325255448204772, 
    0.02005015051157346, 0.019767986492401437, 0.019478643914144413, 
    0.019182244273756657, 0.018879160336012685, 0.018570047920108617, 
    0.018255854946701181, 0.017937788401738496, 0.01761730315471674, 
    0.017296023108912557, 0.016975654110181683, 0.016657899551586718, 
    0.016344391852109307, 0.016036645281564902, 0.015736013759093628, 
    0.015443673621155212, 0.015160592937146725, 0.014887508267720267, 
    0.014624904753501131, 0.014373002247745282, 0.01413176787705756, 
    0.013900921428115326, 0.013679985182289071, 0.013468303018408519, 
    0.013265109007954343, 0.013069554417265396, 0.012880750898381274, 
    0.01269779775686369, 0.012519823311946999, 0.012345991294765081, 
    0.012175530717546049, 0.012007748255707822, 0.011842054749867062, 
    0.011677952659014107, 0.011515076364275909, 0.01135317445076834, 
    0.011192113783658543, 0.01103186590353223, 0.010872518906428416, 
    0.010714260518802369, 0.010557358334074706, 0.010402161068550467, 
    0.010249074633122555, 0.010098534863396553, 0.0099510043311175061, 
    0.0098069667762548662, 0.009666922890269802, 0.0095314063872866568, 
    0.0094009716592678219, 0.009276182022906157, 0.0091575843655073205, 
    0.009045681552172528, 0.008940918948985032, 0.0088436504789501345, 
    0.0087541232784568747, 0.0086724744505525045, 0.0085986926189532947, 
    0.0085326419405770508, 0.0084740280248779103, 0.0084223965443590756, 
    0.0083771023727316589, 0.0083373398834524631, 0.0083021004794409468, 
    0.0082701963626150114, 0.0082402491788699742, 0.0082107127137669121, 
    0.008179882000944709, 0.0081459400410697647, 0.008106981534437091, 
    0.008061075462139378, 0.0080063241718455538, 0.007940928329395084, 
    0.0078632362630997234, 0.0077718376516493761, 0.0076656102302578482, 
    0.00754376086725571, 0.0074058650470062957, 0.0072518761732252119, 
    0.0070821248082984321, 0.0068972936983292881, 0.0066983638167050228, 
    0.0064865582974995718, 0.006263246340830044, 0.006029849885558331, 
    0.0057877594622386362, 0.0055382699024062506, 0.0052825372927147096, 
    0.0050216006629216006, 0.0047564121251672488, 0.0044878528235037735, 
    0.0042168256069915677, 0.0039442734246051625, 0.0036712493653070621, 
    0.0033989305173691142, 0.0031286452442470802, 0.0028618429306801222, 
    0.0026001461278685979, 0.0023452415865572204, 0.0020989120246296582, 
    0.0018629531008646344, 0.0016391900688358424, 0.0014294332343477618, 
    0.0012354676827946976, 0.0010590254391373312, 0.0009018084882452856, 
    0.00076544351233394413, 0.00065147771506177468, 0.00056139349902307382, 
    0.00049657998421726631, 0.00045839106620080877, 0.00044810317669028137, 
    0.00046700229592946366, 0.00051635770058200154, 0.00059750534490066697, 
    0.00071180016731183134, 0.0008606698080941221, 0.0010455716046061739, 
    0.0012679299885568771, 0.0015291040973606034, 0.0018302521330808665, 
    0.0021722102457757352, 0.0025554132595294048, 0.0029797858762832504, 
    0.0034446633583923737, 0.0039487763975558053, 0.0044902041915386879, 
    0.0050664521754938529, 0.0056744772264307238, 0.0063107716636720476, 
    0.0069714800054325697, 0.0076524788514225391, 0.0083494936868144728, 
    0.0090582016209602625, 0.0097743522610979627, 0.010493868167504944, 
    0.011212971623027538, 0.01192829154054429, 0.012636963068009301, 
    0.013336724683596743, 0.014025997316054202, 0.014703989980056861, 
    0.015370678615632318, 0.016026823293313414, 0.01667392642451225, 
    0.017314024746986477, 0.017949458545323295, 0.018582595025836559, 
    0.019215516155294488, 0.01984959416645166, 0.02048540940490275, 
    0.021122521791042258, 0.021759557670516124, 0.022394365162327699, 
    0.023024183134191849, 0.02364590095296672, 0.024256345699700598, 
    0.024852589775201654, 0.025432086297146664, 0.025992846725186144, 
    0.026533473500569935, 0.027052887635190061, 0.027550147862070332, 
    0.02802410196719465, 0.028473000221212956, 0.028894431747796975, 
    0.029284895637113187, 0.029639833542769431, 0.029954147177426171, 
    0.030222116726952374, 0.030437852700958758, 0.030595917416404876, 
    0.030690929660422722, 0.030718073061851106, 0.030673037308019666,
  // Fqt-Na(2, 0-1999)
    1, 0.99912105988048761, 0.99649431430235447, 0.99214939633524424, 
    0.98613454766767183, 0.97851526931981658, 0.9693725482592509, 
    0.9588007641194114, 0.94690537480768566, 0.93380048829018536, 
    0.91960641990040382, 0.90444731509693077, 0.88844891025498252, 
    0.87173648602140041, 0.85443304746199167, 0.83665775251747188, 
    0.81852459601410166, 0.80014135550659859, 0.78160876769897525, 
    0.7630199404667487, 0.74445996876020182, 0.72600573781107203, 
    0.70772589584663115, 0.6896809640586431, 0.67192357429325611, 
    0.65449879402794287, 0.63744452420884645, 0.62079195230581852, 
    0.6045660355523621, 0.58878600595762021, 0.57346589674994952, 
    0.55861505722554006, 0.54423867668133763, 0.53033827835587766, 
    0.51691219446922876, 0.50395600763635762, 0.49146295901773734, 
    0.47942432188046352, 0.46782973581201248, 0.45666751505348668, 
    0.44592491575779963, 0.43558838476850109, 0.42564377517341118, 
    0.41607654370198743, 0.40687191975576731, 0.39801505432691042, 
    0.38949114564790704, 0.38128554942113274, 0.37338386848151278, 
    0.36577202899813011, 0.35843633381709128, 0.35136351549024669, 
    0.34454076719148152, 0.33795577284561928, 0.33159672017762143, 
    0.3254523157535017, 0.31951178823757886, 0.31376488516183609, 
    0.30820186978239744, 0.30281351485266739, 0.29759108180995564, 
    0.29252630652294187, 0.28761138102753125, 0.28283892215877715, 
    0.27820195157505417, 0.273693865265279, 0.26930840545613621, 
    0.26503963840377281, 0.2608819273602378, 0.25682991277540324, 
    0.25287849395801554, 0.24902280737492538, 0.2452582141847599, 
    0.24158028062799161, 0.23798476675957911, 0.23446761495289165, 
    0.23102494197384016, 0.22765303259620912, 0.2243483333355222, 
    0.22110745684516564, 0.21792717453664534, 0.21480442386727791, 
    0.21173630712311722, 0.20872009727591748, 0.20575324433987349, 
    0.20283338486560767, 0.19995834763950848, 0.19712616602665903, 
    0.19433508725384629, 0.19158356954593395, 0.18887028780429704, 
    0.18619412987665473, 0.18355419056258207, 0.18094976792444784, 
    0.17838035680335645, 0.17584564640758024, 0.17334550591961984, 
    0.17087997560404111, 0.16844924578108703, 0.16605363923903277, 
    0.16369358641518239, 0.16136960259279443, 0.15908226225065356, 
    0.15683217667243296, 0.15461997543772982, 0.15244628690822126, 
    0.15031172083822672, 0.14821685644480276, 0.14616223649289212, 
    0.14414835719396785, 0.1421756686407446, 0.14024457188137146, 
    0.13835542424927072, 0.13650853786186035, 0.13470418341675461, 
    0.13294258766972664, 0.13122392431436877, 0.129548305574995, 
    0.12791577634775864, 0.12632630536352948, 0.12477978290050029, 
    0.12327602106347224, 0.1218147541369794, 0.12039564310348384, 
    0.11901827548629813, 0.11768216569121048, 0.11638675360276542, 
    0.11513140084048022, 0.11391538663162518, 0.11273790106827408, 
    0.11159804112695292, 0.11049481178625804, 0.10942712600696167, 
    0.10839380456938535, 0.10739357432575777, 0.1064250695376051, 
    0.10548683218147963, 0.10457731564640593, 0.10369489500347505, 
    0.10283788056463103, 0.10200453471892679, 0.10119309114662685, 
    0.10040177496624808, 0.099628818161406063, 0.098872478593829985, 
    0.098131047187515447, 0.097402865538574718, 0.096686328444433284, 
    0.095979892297920991, 0.09528207836496827, 0.094591476897142174, 
    0.093906748893847106, 0.093226629881098033, 0.092549928292810363, 
    0.091875528332355377, 0.091202393847521671, 0.090529566403360351, 
    0.089856172550052613, 0.089181426820213919, 0.088504641076780438, 
    0.087825227747875934, 0.087142707454558557, 0.086456706459864099, 
    0.08576695402844059, 0.085073270705506188, 0.084375556632757295, 
    0.083673772837915689, 0.082967924590354389, 0.082258047473518892, 
    0.081544192581480185, 0.08082642587677899, 0.080104826875119384, 
    0.079379496969531643, 0.078650562131526283, 0.077918182085402035, 
    0.077182553185198594, 0.076443916397359438, 0.075702559928552626, 
    0.074958821611633752, 0.074213092806722045, 0.073465817160229555, 
    0.072717490533762738, 0.071968658510261393, 0.071219912729760165, 
    0.070471878671950941, 0.069725212360709332, 0.068980584064405798, 
    0.068238673170119224, 0.06750015747015875, 0.066765709644550544, 
    0.066035990560501148, 0.065311653938404643, 0.064593343979113191, 
    0.063881693059251413, 0.063177321644652396, 0.062480832608961548, 
    0.061792803332056577, 0.061113778640685158, 0.060444254489074381, 
    0.059784666966546648, 0.059135373993322672, 0.05849665395649295, 
    0.057868688676299546, 0.057251567819145338, 0.056645285195199409, 
    0.056049747361784766, 0.055464776416247835, 0.05489012567755186, 
    0.054325489777460927, 0.053770518289954494, 0.053224834616606126, 
    0.052688048226062892, 0.052159773785439498, 0.051639646666968332, 
    0.051127337032586963, 0.050622564450003862, 0.050125106226947269, 
    0.049634803778034094, 0.049151563063741709, 0.048675352501711178, 
    0.048206194759850052, 0.047744159973731846, 0.047289354261854981, 
    0.04684191008983872, 0.046401975930812848, 0.045969708924964249, 
    0.045545262562720179, 0.045128783344508643, 0.044720400992703219, 
    0.044320218900353328, 0.04392831376491417, 0.043544721321218477, 
    0.043169435659408006, 0.042802402573075937, 0.042443514294861574, 
    0.042092601914058878, 0.041749428475104718, 0.041413688129447186, 
    0.041084997510049709, 0.040762896967191875, 0.040446861176774623, 
    0.040136305566859889, 0.039830610573219072, 0.039529137947589985, 
    0.039231264995997814, 0.03893640096713237, 0.03864401283160282, 
    0.038353639010321926, 0.038064901585414451, 0.037777513533737386, 
    0.037491278691656457, 0.037206095656130769, 0.03692195317222579, 
    0.036638926027235452, 0.036357172727263333, 0.036076935968301617, 
    0.035798533797378886, 0.03552236296377851, 0.035248886268979603, 
    0.034978621712293718, 0.034712125100334619, 0.034449967667106854, 
    0.034192713943332571, 0.033940890322907716, 0.03369496204121903, 
    0.033455313191721341, 0.033222223799836609, 0.032995867246074818, 
    0.032776303966557001, 0.032563487583546179, 0.032357278218220611, 
    0.03215745203423253, 0.031963720612461187, 0.031775743903200884, 
    0.03159314900387223, 0.031415544753749178, 0.031242535811405438, 
    0.031073735761289051, 0.030908778454553608, 0.030747329592805392, 
    0.030589094069638039, 0.030433823277282432, 0.03028131746419508, 
    0.030131426822595384, 0.029984052492249214, 0.029839141112491713, 
    0.029696683051047754, 0.029556703172973885, 0.029419256216595663, 
    0.029284417270626133, 0.029152269640803159, 0.029022898298845662, 
    0.028896377176371502, 0.028772759948969835, 0.028652079392059847, 
    0.028534340105817627, 0.028419521733805533, 0.028307576451651807, 
    0.028198430317221291, 0.028091979954103199, 0.027988086009381505, 
    0.027886566573471057, 0.027787186954326078, 0.027689654907100882, 
    0.027593611708561481, 0.027498633100909928, 0.027404225529528915, 
    0.027309830467722524, 0.027214824467061909, 0.027118529383112561, 
    0.027020215191193513, 0.026919114188448015, 0.026814433994195974, 
    0.026705377076106061, 0.026591158826197756, 0.026471032945826457, 
    0.026344314500039951, 0.026210401277726059, 0.026068796740027277, 
    0.025919129309309372, 0.025761165184845582, 0.025594822705853452, 
    0.025420182581703574, 0.025237491329972852, 0.025047163701266095, 
    0.024849776376042378, 0.024646057096128018, 0.024436871621371363, 
    0.024223200974167781, 0.024006124249598186, 0.023786795892463349, 
    0.023566431273800589, 0.023346289810962949, 0.023127663001654534, 
    0.022911865894134974, 0.022700223480077615, 0.022494058615477746, 
    0.022294673922669275, 0.022103333198882014, 0.021921236243612873, 
    0.021749494497132638, 0.021589103672357671, 0.021440918983323239, 
    0.021305633573773502, 0.021183755573003362, 0.021075594214323118, 
    0.020981244357683868, 0.020900578981842256, 0.020833249492842151, 
    0.020778684668247869, 0.020736105267695593, 0.020704538481113352, 
    0.020682838171943461, 0.020669710698107465, 0.02066374146196194, 
    0.020663422826387896, 0.020667181981310224, 0.020673407304866987, 
    0.02068047589074079, 0.020686781114570913, 0.020690757367679977, 
    0.020690902847327775, 0.020685803608075589, 0.020674157287878539, 
    0.020654795528156782, 0.020626701399766554, 0.02058902455268102, 
    0.020541089136426858, 0.020482396097356987, 0.020412620767156206, 
    0.020331603637867308, 0.020239338716564081, 0.020135959230763015, 
    0.020021722569378512, 0.01989699288875782, 0.019762224793054981, 
    0.019617951164963857, 0.019464770112957497, 0.019303335720232628, 
    0.01913435338697432, 0.018958574546346224, 0.018776797287663884, 
    0.018589864532031021, 0.01839866313948452, 0.018204121942863753, 
    0.018007202889823097, 0.017808897965710453, 0.017610211683164557, 
    0.017412154387368029, 0.017215727862466133, 0.017021918694666235, 
    0.016831691382745644, 0.016645981247930319, 0.016465686247196649, 
    0.016291654744041581, 0.016124672097747959, 0.015965446975628787, 
    0.015814598598942058, 0.015672649591276646, 0.01554002073043163, 
    0.015417028512631695, 0.015303890351634679, 0.015200725245077821, 
    0.015107555377808862, 0.015024307813183608, 0.014950811441773066, 
    0.014886796450637329, 0.014831897351230895, 0.014785658225193146, 
    0.014747539553942639, 0.014716929260558486, 0.014693150429309878, 
    0.014675474790050552, 0.014663134514784758, 0.014655331235777898, 
    0.014651249677985867, 0.014650069756004885, 0.014650979458538783, 
    0.014653189896132244, 0.014655946967614058, 0.014658546006831188, 
    0.014660340692965425, 0.014660752753912928, 0.014659281831935704, 
    0.014655512222126261, 0.014649117507761867, 0.014639867955032467, 
    0.014627631666127024, 0.014612377774988621, 0.014594176503533503, 
    0.014573194989330129, 0.014549692008691231, 0.014524009109492137, 
    0.014496563558200335, 0.014467839975234273, 0.014438376922080234, 
    0.014408751935601712, 0.014379569230918985, 0.014351439380463784, 
    0.014324957680888262, 0.014300683138415822, 0.014279120803418836, 
    0.014260701890453505, 0.014245775319568747, 0.014234599865617852, 
    0.014227338884391833, 0.014224064723834341, 0.014224758159394349, 
    0.014229316093432953, 0.014237553503592033, 0.014249206367325878, 
    0.014263937929503714, 0.014281337077177851, 0.014300924748826629, 
    0.014322162349020867, 0.014344461773586527, 0.014367198206275404, 
    0.014389723189252777, 0.01441137915215273, 0.014431508842917551, 
    0.014449470746634819, 0.014464645015976383, 0.014476440904693331, 
    0.014484304558880501, 0.014487726972667994, 0.014486246902943494, 
    0.014479460698732885, 0.014467025799621315, 0.014448663576708033, 
    0.014424161491953559, 0.014393371174070232, 0.014356207211302992, 
    0.014312637403480356, 0.014262680973705073, 0.014206404042920886, 
    0.014143914026708334, 0.014075359764228263, 0.014000931630882122, 
    0.013920862566924068, 0.013835429846965657, 0.013744960112955704, 
    0.013649828381485258, 0.01355046049531905, 0.013447331214732792, 
    0.013340961694979149, 0.013231909881445141, 0.01312076290606992, 
    0.013008124121078001, 0.01289459704981828, 0.012780773399136249, 
    0.012667216344234665, 0.012554453952723532, 0.01244297013811577, 
    0.012333202837746547, 0.01222554560132926, 0.012120352385035517, 
    0.012017935543456273, 0.011918565690963674, 0.011822465129327286, 
    0.011729798102881637, 0.01164066449902167, 0.011555085710178123, 
    0.011473004126969791, 0.011394280115265958, 0.011318692264122977, 
    0.0112459453080699, 0.0111756807464993, 0.011107488993400349, 
    0.011040924636074097, 0.010975521757863939, 0.010910809539987893, 
    0.010846331194427737, 0.010781656008958354, 0.010716396395618737, 
    0.010650219798476636, 0.010582855531384815, 0.010514098511539088, 
    0.010443809238229032, 0.01037190934734687, 0.010298374224868619, 
    0.010223220462330481, 0.010146497418218119, 0.010068270373994518, 
    0.0099886079008477437, 0.0099075750651532301, 0.0098252243810658772, 
    0.0097415990516257663, 0.0096567361348382664, 0.0095706705200893118, 
    0.0094834473521255257, 0.0093951220359743699, 0.009305770719440512, 
    0.0092154874691223482, 0.0091243915955818971, 0.0090326234639058426, 
    0.008940343919382485, 0.008847728340256723, 0.0087549681490745063, 
    0.0086622646623198719, 0.0085698294087724197, 0.0084778824218756099, 
    0.0083866558375580783, 0.0082963895022248775, 0.0082073316360996296, 
    0.0081197346711254156, 0.0080338514466874837, 0.007949927968875798, 
    0.0078681929806889393, 0.0077888526045021148, 0.0077120772480969461, 
    0.0076379926035776658, 0.0075666662165022949, 0.0074980957955654935, 
    0.0074322015775273483, 0.0073688183165847403, 0.0073076931300142482, 
    0.0072484897016654726, 0.0071907909057648111, 0.0071341139246269506, 
    0.0070779217777131084, 0.0070216435255088996, 0.0069646882224591875, 
    0.0069064623579152759, 0.0068463817638404981, 0.0067838838322729052, 
    0.0067184414443697705, 0.0066495774391862805, 0.0065768763658277983, 
    0.0065000047427474193, 0.0064187209270435957, 0.0063328896617207923, 
    0.0062424875424783024, 0.0061476111033753125, 0.0060484755689869316, 
    0.0059454181973273325, 0.0058388873680258087, 0.0057294401881384299, 
    0.0056177277331306919, 0.005504481928152536, 0.0053904989503166263, 
    0.0052766209895310848, 0.0051637152200444056, 0.0050526580366589864, 
    0.0049443125141299862, 0.0048395138791301195, 0.0047390512216646296, 
    0.0046436510017430106, 0.0045539600366878638, 0.004470529288249073, 
    0.0043938004250046753, 0.0043240921684310936, 0.0042615958735117126, 
    0.0042063657455159191, 0.0041583241061604881, 0.004117266951667602, 
    0.0040828761318629832, 0.0040547383206190352, 0.0040323634795055695, 
    0.0040152082453869253, 0.0040026976846115562, 0.0039942464783452722, 
    0.0039892801324899665, 0.0039872548528377474, 0.0039876684725918491, 
    0.0039900752775986273, 0.0039940890306146837, 0.0039993825803050984, 
    0.0040056820576706408, 0.0040127593817053308, 0.0040204201988022787, 
    0.0040284927338598581, 0.0040368240141338742, 0.004045266165138426, 
    0.004053673042711277, 0.0040618948872593735, 0.0040697711065304266, 
    0.0040771258578191708, 0.004083762053102017, 0.0040894536345671504, 
    0.0040939363139127763, 0.0040969012711851178, 0.0040979874430922599, 
    0.0040967752182423404, 0.0040927845761901567, 0.0040854736810598336, 
    0.0040742423149432109, 0.004058439823913791, 0.0040373769042843597, 
    0.004010333127719411, 0.0039765712609276666, 0.0039353527636944614, 
    0.0038859509823684188, 0.0038276695488895589, 0.0037598624925365047, 
    0.0036819535483127181, 0.0035934548179082215, 0.0034939841780846663, 
    0.0033832766612166242, 0.0032611914255935145, 0.0031277193946144272, 
    0.0029829788819948247, 0.002827214848444227, 0.0026607886320083709, 
    0.0024841732410529967, 0.0022979420264510556, 0.0021027602051493658, 
    0.001899377864634792, 0.001688615745870292, 0.0014713614885826795, 
    0.0012485544814621662, 0.0010211806696003413, 0.00079026182118146723, 
    0.00055684769629697891, 0.00032200755795378389, 8.6820216336335604e-05, 
    -0.0001476360995902161, -0.00038029835040865223, -0.00061013685545186847, 
    -0.00083617778240387564, -0.0010575265769635889, -0.0012734005492026526, 
    -0.0014831475333274859, -0.0016862663593682067, -0.0018824062833128837, 
    -0.0020713644238249218, -0.0022530727616403672, -0.0024275796210578363, 
    -0.0025950350320303921, -0.0027556733181881739, -0.0029098002886982395, 
    -0.0030577833312898459, -0.0032000388909264304, -0.0033370285559407046, 
    -0.0034692483030512983, -0.003597224898808479, -0.0037215061153627548, 
    -0.0038426649621196005, -0.0039612892994424194, -0.0040779806439835238, 
    -0.004193355702301213, -0.0043080407135116378, -0.0044226708066318213, 
    -0.0045378869635228029, -0.0046543296253078606, -0.0047726281596437541, 
    -0.0048933839102865582, -0.0050171485098935032, -0.0051443992724999887, 
    -0.0052755156778153687, -0.0054107606178576372, -0.0055502702241919926, 
    -0.0056940433947107131, -0.0058419413138329698, -0.0059937011957283343, 
    -0.0061489519498843549, -0.0063072492724086694, -0.0064681104905218618, 
    -0.006631054840775653, -0.0067956404066665871, -0.0069614881434771313, 
    -0.0071283054762251337, -0.0072959010467620522, -0.0074641942185381012, 
    -0.0076332195596432329, -0.0078031267968312456, -0.0079741740723949222, 
    -0.0081467164629476646, -0.0083211918640250515, -0.0084980998014824744, 
    -0.0086779834552233211, -0.0088614054012399295, -0.0090489231411312078, 
    -0.0092410735282890642, -0.0094383460222495427, -0.0096411727218808519, 
    -0.0098499098320790728, -0.010064826618688936, -0.010286095120950644, 
    -0.010513780239366468, -0.010747831428415009, -0.010988078258458107, 
    -0.011234222684667675, -0.011485838638801253, -0.011742370060766744, 
    -0.012003137944276585, -0.012267344364408017, -0.012534087119250147, 
    -0.012802376398603607, -0.013071154066226585, -0.013339320156399015, 
    -0.013605756056164825, -0.013869352850950194, -0.014129029089965463, 
    -0.014383754727195245, -0.014632572212606696, -0.014874610369289096, 
    -0.015109101057163381, -0.015335393941195609, -0.015552966629298682, 
    -0.015761435007440146, -0.015960555725557306, -0.016150231002437898, 
    -0.016330504945651379, -0.016501560774180992, -0.016663719717989696, 
    -0.016817433458281482, -0.016963275335179828, -0.017101924536088511, 
    -0.017234146365496823, -0.01736076699431547, -0.017482643209992866, 
    -0.017600637825684523, -0.017715584660800098, -0.017828262660683152, 
    -0.017939361985229683, -0.018049461067173339, -0.018158999368903708, 
    -0.018268259629398553, -0.018377355279521647, -0.018486223623647408, 
    -0.01859462740863491, -0.018702162581819406, -0.018808273850730819, 
    -0.018912277587194069, -0.019013387292613159, -0.019110742858079829, 
    -0.019203441328862376, -0.019290562557876024, -0.019371194658961546, 
    -0.019444458362081918, -0.019509524849294215, -0.019565627864825366, 
    -0.019612073429163972, -0.019648243689218147, -0.019673599675820719, 
    -0.019687682336680806, -0.019690108222869235, -0.019680570988575192, 
    -0.019658839883343226, -0.019624762859539312, -0.019578267576490466, 
    -0.019519359840426201, -0.019448125249302187, -0.019364722397318301, 
    -0.019269381893795727, -0.019162394286057181, -0.019044104575550551, 
    -0.018914902077472102, -0.01877520592729514, -0.018625460860444983, 
    -0.018466125047954494, -0.018297665767243856, -0.018120552220794096, 
    -0.017935252742750089, -0.017742239234180099, -0.017541985157707607, 
    -0.017334975934700042, -0.017121716564522649, -0.016902740941267768, 
    -0.016678617928574838, -0.016449956863681635, -0.016217411518088656, 
    -0.015981674680042062, -0.015743474775585558, -0.015503571326244192, 
    -0.015262747951851523, -0.015021806897065889, -0.014781562275720708, 
    -0.014542829626768457, -0.014306416007591619, -0.014073110006962847, 
    -0.013843664248346444, -0.013618784311303641, -0.013399115019828087, 
    -0.013185225858916589, -0.012977599195548637, -0.012776620712399, 
    -0.012582570527717114, -0.012395615566662809, -0.012215807563162009, 
    -0.012043076984965411, -0.01187723147578554, -0.011717956699797904, 
    -0.011564815728144414, -0.011417259060793801, -0.01127462960290466, 
    -0.011136178804436018, -0.011001082511533341, -0.010868457803530905, 
    -0.010737388950335172, -0.010606943874101722, -0.010476197874476142, 
    -0.01034425176036903, -0.010210252683566243, -0.010073413178888695, 
    -0.0099330267722957128, -0.0097884821904641716, -0.0096392803870536808, 
    -0.0094850411135086327, -0.0093255123889794886, -0.0091605718351285576, 
    -0.0089902269771765155, -0.008814612376709963, -0.008633984903314372, 
    -0.0084487146931487428, -0.0082592729061243455, -0.0080662217428389381, 
    -0.0078701990251133277, -0.0076719039531601731, -0.0074720799814074219, 
    -0.0072715073322813916, -0.0070709908433623488, -0.00687134931035812, 
    -0.0066734143446038428, -0.0064780190999295479, -0.0062859959192832649, 
    -0.0060981643582098677, -0.0059153199423109711, -0.0057382174229003904, 
    -0.0055675527333121835, -0.0054039434894363574, -0.0052479107031839136, 
    -0.0050998658758431821, -0.0049600981482575803, -0.0048287673223042869, 
    -0.00470590285753846, -0.004591404216596707, -0.0044850476475524117, 
    -0.0043864913927437509, -0.0042952880215943656, -0.0042108942525419454, 
    -0.0041326862151050033, -0.0040599764524607675, -0.0039920299897861188, 
    -0.0039280842002776574, -0.0038673693142087869, -0.0038091248751502089, 
    -0.0037526130846045891, -0.0036971308517183121, -0.0036420156149922465, 
    -0.0035866508463071782, -0.0035304675893278559, -0.0034729443128078737, 
    -0.0034136058302363112, -0.0033520215894146596, -0.0032878039253872084, 
    -0.00322060353343963, -0.0031501135552170437, -0.0030760632124411528, 
    -0.0029982220503553805, -0.0029163938412776255, -0.0028304211834277279, 
    -0.0027401848980616022, -0.0026456041376517435, -0.0025466423240205751, 
    -0.0024433081459896153, -0.0023356648482307121, -0.0022238306014002798, 
    -0.0021079830932045672, -0.0019883583386902095, -0.0018652458624164527, 
    -0.0017389806437777776, -0.0016099333063340508, -0.0014784940856847908, 
    -0.0013450587375085268, -0.0012100112353764713, -0.0010737095723267842, 
    -0.00093647480001137428, -0.00079858534841475667, 
    -0.00066028144967200946, -0.0005217783690110952, -0.00038328165485558259, 
    -0.00024500532966714185, -0.00010718814693641077, 2.9897961980814534e-05, 
    0.00016594382536566513, 0.00030060296075150295, 0.00043349467605984589, 
    0.00056420755971994265, 0.00069230401745853107, 0.00081732599772374047, 
    0.00093880277315988537, 0.001056257732046027, 0.0011692183353404224, 
    0.0012772274366697762, 0.0013798496962048872, 0.0014766833239780479, 
    0.00156736882128997, 0.0016515937422441956, 0.0017291028774336502, 
    0.0017996998488634802, 0.0018632537268334507, 0.0019197020991424168, 
    0.0019690513859487195, 0.0020113785973423859, 0.0020468307107084642, 
    0.0020756200486205974, 0.0020980191241608531, 0.0021143603177208687, 
    0.0021250297850639514, 0.0021304657828638981, 0.0021311502655944714, 
    0.0021276058768831046, 0.0021203875621511291, 0.002110069990358121, 
    0.0020972377881207549, 0.0020824737266679104, 0.0020663470566189891, 
    0.0020494043979509035, 0.0020321618366709523, 0.0020150975712582165, 
    0.0019986458317030427, 0.0019831912843119846, 0.00196906406256484, 
    0.0019565373764489774, 0.0019458205206931429, 0.0019370549377269162, 
    0.0019303045885549113, 0.0019255522605818259, 0.0019226931022623362, 
    0.0019215310672544967, 0.0019217852003759689, 0.0019230898964113774, 
    0.0019250054832600336, 0.0019270263681905645, 0.0019285914394276172, 
    0.0019290962850563047, 0.001927902180392472, 0.0019243501826038238, 
    0.0019177740992144441, 0.001907515053258811, 0.0018929363760748024, 
    0.0018734364879603696, 0.0018484717167375603, 0.0018175640198495374, 
    0.0017803156056866581, 0.0017364172320732997, 0.0016856539800010402, 
    0.0016278999197164446, 0.0015631149548274224, 0.0014913302365043418, 
    0.0014126359515139997, 0.0013271628600052981, 0.0012350651372189405, 
    0.0011365065067626139, 0.0010316455009320121, 0.00092062795308527198, 
    0.00080358056263420954, 0.00068060502066151322, 0.00055178204945192173, 
    0.00041717227683982596, 0.00027682868398527121, 0.00013080754076994828, 
    -2.0818919982420244e-05, -0.0001779461887925003, -0.00034042160279715674, 
    -0.00050803292220826793, -0.00068049437676615703, 
    -0.00085743611790532043, -0.001038394542130305, -0.0012228045652400176, 
    -0.001409994763497037, -0.0015991853836977016, -0.0017894956307052347, 
    -0.0019799529672776617, -0.0021695120411721514, -0.002357078870264805, 
    -0.0025415403619769451, -0.0027217930473897997, -0.0028967757349409088, 
    -0.0030654914350475649, -0.0032270278620521922, -0.0033805701239705164, 
    -0.0035254125574309498, -0.003660965550510467, -0.0037867629024635977, 
    -0.0039024571018782556, -0.0040078213565038264, -0.0041027384933678291, 
    -0.0041871848855593611, -0.0042612186323752761, -0.0043249589617534914, 
    -0.0043785671814827835, -0.0044222287994194883, -0.0044561403748578261, 
    -0.004480494856210859, -0.0044954743887769127, -0.0045012453468623159, 
    -0.0044979540330404716, -0.0044857319595085357, -0.0044646971714159146, 
    -0.0044349605599685749, -0.0043966348527184835, -0.004349842443038052, 
    -0.0042947252694152472, -0.0042314561166706833, -0.004160241792551117, 
    -0.0040813314705008775, -0.0039950180957935141, -0.0039016409516833745, 
    -0.0038015810814104847, -0.0036952583609433497, -0.0035831262497905817, 
    -0.0034656651649613629, -0.0033433755630881959, -0.0032167681961641882, 
    -0.0030863565558719671, -0.0029526473891917822, -0.0028161335994483176, 
    -0.0026772901422899994, -0.0025365716065720812, -0.002394413669439501, 
    -0.0022512386407321336, -0.0021074647659900256, -0.0019635164777209464, 
    -0.001819835405081812, -0.0016768929208249347, -0.0015351966931837291, 
    -0.0013952918113041622, -0.001257763906371554, -0.0011232339586071836, 
    -0.00099235472823330068, -0.00086580823189429373, 
    -0.00074430105214389147, -0.00062855897102324031, 
    -0.00051932236314210407, -0.00041733255531835344, 
    -0.00032332155885456734, -0.00023799515403925917, 
    -0.00016201700196143251, -9.5986502192151361e-05, 
    -4.0421567371691849e-05, 4.2608944519767489e-06, 3.7759776187584043e-05, 
    5.9895684334576875e-05, 7.0618568845255453e-05, 6.9998270124870866e-05, 
    5.8219325711507603e-05, 3.556179770362552e-05, 2.3826275619895625e-06, 
    -4.0903587979888964e-05, -9.3845253127374266e-05, 
    -0.00015596907720396116, -0.00022679175815658412, 
    -0.00030582274315557384, -0.00039256414380424681, 
    -0.00048650488244301494, -0.00058711298101772819, 
    -0.00069383029232814616, -0.00080606869281638397, 
    -0.00092320780683834743, -0.0010445934376953053, -0.001169536919097085, 
    -0.0012973099550004611, -0.0014271372071720028, -0.0015581948233519384, 
    -0.0016896058086293166, -0.0018204367181283525, -0.0019497005756477521, 
    -0.0020763555508053122, -0.002199308237928071, -0.002317419375585523, 
    -0.0024295123215479376, -0.0025343839665776507, -0.0026308196945143839, 
    -0.0027176172068818262, -0.0027936024504715351, -0.0028576590939048308, 
    -0.0029087488651005529, -0.002945936832351679, -0.0029684139493513315, 
    -0.0029755155618761834, -0.0029667426255875575, -0.002941775812759233, 
    -0.0029004934782827473, -0.0028429802743198118, -0.0027695372077005255, 
    -0.0026806848001932927, -0.00257716092961661, -0.0024599141281565888, 
    -0.0023300921387077473, -0.0021890238585578689, -0.0020381960799721118, 
    -0.0018792292629499726, -0.0017138447230736799, -0.0015438375526304828, 
    -0.0013710423354861257, -0.0011973070887451019, -0.0010244657633209607, 
    -0.00085431246053802577, -0.00068857842252367297, 
    -0.00052891258013532572, -0.00037686344291082337, 
    -0.00023385990378157887, -0.00010120229122670291, 1.9944270125330182e-05, 
    0.00012855996668834275, 0.00022376775158826346, 0.00030483405160952045, 
    0.0003711651339638099, 0.00042230311342016601, 0.00045791750888858607, 
    0.00047780214919723458, 0.00048186654061374459, 0.00047013177620526178, 
    0.00044272851018160961, 0.00039989088298874551, 0.00034195357078565473, 
    0.00026934662097969416, 0.00018258565936731872, 8.2266774401685818e-05, 
    -3.0946882205885802e-05, -0.00015633342800374235, 
    -0.00029311991363962977, -0.00044048786491455777, 
    -0.00059757878702225453, -0.00076349625269004056, 
    -0.00093731098772688814, -0.0011180627027493691, -0.0013047638749393137, 
    -0.0014964044280832173, -0.001691964837197159, -0.001890424645912025, 
    -0.0020907758538588833, -0.00229204164275182, -0.0024932888811589789, 
    -0.0026936463685056054, -0.0028923207161712801, -0.003088606390981899, 
    -0.0032818970037410237, -0.0034716953752911006, -0.0036576120872289218, 
    -0.0038393660452344441, -0.0040167781830304219, -0.0041897655824816782, 
    -0.0043583249573565805, -0.004522523146094499, -0.0046824870126796836, 
    -0.0048383905369924094, -0.0049904497678220317, -0.0051389163502690996, 
    -0.0052840671783418117, -0.0054261954383913362, -0.0055655994679683829, 
    -0.0057025709937984018, -0.0058373778582607415, -0.0059702525528231498, 
    -0.0061013813402673624, -0.0062308956706761025, -0.0063588655862413853, 
    -0.0064852974300859531, -0.0066101354776925639, -0.0067332606298259974, 
    -0.0068544926798761183, -0.0069735846481295887, -0.0070902244268860508, 
    -0.0072040280065905583, -0.0073145445173502278, -0.0074212532957255457, 
    -0.0075235730048304854, -0.0076208713800281691, -0.0077124820371449925, 
    -0.0077977231517325236, -0.0078759173013196095, -0.0079464141352533404, 
    -0.0080086033142082215, -0.008061928882267087, -0.0081058980574297591, 
    -0.0081400851998205716, -0.0081641367706241901, -0.0081777699899622594, 
    -0.0081807744521037937, -0.0081730090830080798, -0.008154401504509563, 
    -0.0081249457600863963, -0.0080847010718670936, -0.0080337889475587711, 
    -0.0079723888726366213, -0.0079007345130788272, -0.0078191026364173369, 
    -0.0077278066417711616, -0.0076271903813955079, -0.0075176161222659243, 
    -0.0073994598765568511, -0.0072731076525900549, -0.0071389470192158239, 
    -0.0069973714374784767, -0.0068487685430414537, -0.0066935257336052162, 
    -0.0065320220070866925, -0.0063646324888990023, -0.0061917231780022333, 
    -0.00601365892107515, -0.0058308053984592887, -0.0056435354646368931, 
    -0.0054522373243362024, -0.0052573190582502396, -0.0050592165929208548, 
    -0.0048583920787814341, -0.0046553351690358999, -0.0044505589620116581, 
    -0.004244590485650096, -0.0040379612994558165, -0.0038311952427674979, 
    -0.003624799050870806, -0.0034192466335863647, -0.003214969995390836, 
    -0.003012346813215847, -0.0028116937791586496, -0.0026132615664844518, 
    -0.0024172294969704907, -0.0022237167428324424, -0.0020327879210299553, 
    -0.0018444815198019513, -0.0016588169954818057, -0.0014758223136081467, 
    -0.0012955451644422441, -0.0011180481590546967, -0.00094340571184804744, 
    -0.00077168657276267512, -0.00060293079831950501, 
    -0.00043713064677697907, -0.00027421840959640167, 
    -0.00011405944879112881, 4.3541307975498167e-05, 0.00019883089603189825, 
    0.00035208814136532496, 0.00050360335553467736, 0.00065365902086384972, 
    0.00080251470385477659, 0.00095039201139467241, 0.0010974659709191068, 
    0.0012438614980296173, 0.001389649539186973, 0.0015348501121982543, 
    0.0016794325873524564, 0.0018233212181739142, 0.0019663919343765666, 
    0.0021084833011030392, 0.0022493937606918122, 0.0023888897161875797, 
    0.0025267065309647493, 0.0026625520080012198, 0.0027961088702830486, 
    0.0029270363360656051, 0.0030549755754310042, 0.0031795526745821861, 
    0.0033003870366657712, 0.0034170978720085006, 0.0035293104786865473, 
    0.0036366573374326618, 0.003738783898296559, 0.0038353524593988772, 
    0.0039260426027367045, 0.0040105594119880681, 0.0040886379805234298, 
    0.0041600467562932309, 0.0042246043554039804, 0.0042821841717421939, 
    0.0043327229704936514, 0.0043762286384091461, 0.0044127790659613478, 
    0.0044425251896736276, 0.0044656790230930086, 0.0044825068906203108, 
    0.0044933170955556963, 0.004498446213872939, 0.0044982488280437766, 
    0.0044930907348634539, 0.0044833398317527849, 0.0044693694278879481, 
    0.0044515584785882883, 0.0044302916522241734, 0.0044059676225348537, 
    0.0043789980145459593, 0.0043498047506334986, 0.0043188132351617168, 
    0.0042864413865255045, 0.0042530804653482385, 0.0042190863547884681, 
    0.0041847653047666885, 0.0041503725341571953, 0.0041161092572732216, 
    0.004082137743353133, 0.0040485895405434034, 0.0040155797055914455, 
    0.0039832227103260799, 0.003951646085383168, 0.0039210011940587356, 
    0.0038914712344323005, 0.0038632699669803646, 0.0038366449336406363, 
    0.0038118689958507928, 0.0037892313662728199, 0.0037690380114499969, 
    0.0037515975090353457, 0.0037372120349031639, 0.0037261632611974584, 
    0.0037186985573836717, 0.0037150131500010724, 0.0037152341585992201, 
    0.0037194132129864739, 0.0037275132491714404, 0.0037394102191376849, 
    0.0037548973210294531, 0.0037736845995099484, 0.0037954157803077758, 
    0.0038196617616863362, 0.0038459373970282746, 0.0038736962385846297, 
    0.0039023405869924041, 0.0039312214226661863, 0.0039596501562502041, 
    0.0039869023663629656, 0.004012231540547825, 0.0040348812664380805, 
    0.0040541022963173721, 0.0040691633135310342, 0.0040793654768314378, 
    0.0040840494283324287, 0.004082607457360889, 0.0040744842873316261, 
    0.0040591837138198132, 0.0040362639760381652, 0.0040053370788547954, 
    0.0039660641580274722, 0.0039181475363833894, 0.0038613293693151429, 
    0.0037953859816329356, 0.0037201304839086548, 0.0036354185841864601, 
    0.0035411535982003903, 0.0034373018190572476, 0.00332389852379195, 
    0.0032010573627248018, 0.003068975779385408, 0.0029279333282503876, 
    0.0027782887105927139, 0.0026204645518253665, 0.0024549378093468815, 
    0.0022822145444728937, 0.0021028289318880539, 0.0019173307326896321, 
    0.0017262936663747087, 0.0015303217870553188, 0.0013300569984076387, 
    0.0011261904525244229, 0.00091945964640752947, 0.00071064914660790154, 
    0.00050058061784030293, 0.00029009952672588051, 8.0063433277246339e-05, 
    -0.00012867270364402047, -0.00033527247005618903, 
    -0.00053892449614469215, -0.00073885938022233161, 
    -0.00093435149721023841, -0.0011247255881210363, -0.0013093640549853671, 
    -0.0014877005258621416, -0.0016592228820582287, -0.0018234545475485273, 
    -0.0019799533350929391, -0.0021283002944429276, -0.0022680887017414871, 
    -0.002398927202764307, -0.0025204423933132452, -0.0026322931064464133, 
    -0.0027341885093207334, -0.0028258975491593668, -0.0029072651905869403, 
    -0.0029782132102327973, -0.0030387488823711986, -0.0030889576115594015, 
    -0.0031289975033109542, -0.0031590965143959288, -0.0031795484296568946, 
    -0.0031907072619877302, -0.0031929951138696942, -0.0031868948240349974, 
    -0.0031729481299114784, -0.0031517527543978349, -0.0031239393809973427, 
    -0.0030901704059665778, -0.0030511125486734399, -0.0030074327769168538, 
    -0.0029597814857237528, -0.0029087977608707374, -0.0028550929207457189, 
    -0.0027992566907046688, -0.0027418515022204055, -0.0026834122873795798, 
    -0.0026244336958675977, -0.002565367503571084, -0.0025066050931630062, 
    -0.0024484747628516529, -0.0023912224617104578, -0.0023349992843547389, 
    -0.0022798503183833808, -0.0022257028922587465, -0.0021723565501568383, 
    -0.0021194858998355693, -0.0020666444820956835, -0.0020132842795069481, 
    -0.0019587906348500221, -0.0019025261644707932, -0.0018438776372209028, 
    -0.0017823053085384668, -0.001717370198295858, -0.0016487538584732636, 
    -0.0015762636797860524, -0.0014998356309862864, -0.0014195280631564893, 
    -0.0013355165909164914, -0.001248083508739082, -0.0011576060877390734, 
    -0.0010645419660481963, -0.00096941321585831844, -0.00087278732410163494, 
    -0.00077526704911746189, -0.00067747597008692634, 
    -0.00058005413067089607, -0.00048365434478699716, 
    -0.00038893582207064591, -0.00029655767151030323, 
    -0.00020716886462109085, -0.00012139054575045392, 
    -3.9794530194029744e-05, 3.7112139922993392e-05, 0.00010890377711020392, 
    0.00017524143617568425, 0.00023587103730080114, 0.00029060970867514108, 
    0.00033933183601956597, 0.00038195972701842557, 0.00041845413951380769, 
    0.00044881820190270346, 0.00047311095417022341, 0.00049145727132615322, 
    0.0005040635687095892, 0.00051122148302421683, 0.00051329577294396392, 
    0.00051070803776237126, 0.00050391031232193957, 0.00049335534502271624, 
    0.00047947650234354822, 0.0004626811202559256, 0.00044333279290061968, 
    0.00042175441213225594, 0.00039822680818373988, 0.00037298504083103077, 
    0.00034621779372771838, 0.00031806254363140658, 0.00028860866755478232, 
    0.00025789120105070397, 0.00022589817233611455, 0.00019257473639044812, 
    0.00015782213482130219, 0.00012151205006176446, 8.3492301769519644e-05, 
    4.3590431992949097e-05, 1.6243389609140076e-06, -4.2591326628117348e-05, 
    -8.9245736055422047e-05, -0.00013851990370623626, 
    -0.00019058368279315521, -0.00024559047586753414, -0.0003036671157323525, 
    -0.00036491323352627581, -0.0004294092278419492, -0.0004972221653332193, 
    -0.00056841504885727268, -0.00064306531029090079, 
    -0.00072127035439758657, -0.00080315707819160356, 
    -0.00088888477598396301, -0.0009786353522431685, -0.0010726077696418086, 
    -0.0011710047845175969, -0.0012740121228851506, -0.0013817755148048854, 
    -0.0014943821645896545, -0.001611840807309826, -0.0017340585817883008, 
    -0.0018608373269747951, -0.0019918660938818924, -0.0021267254117239643, 
    -0.0022648985832371088, -0.0024057877179170972, -0.0025487394217996737, 
    -0.0026930614417222647, -0.0028380516092302997, -0.0029830157823221033, 
    -0.0031272884244074343, -0.0032702559508194229, -0.0034113708178256296, 
    -0.0035501677692682527, -0.0036862753001187035, -0.0038194152295473001, 
    -0.0039493970107052174, -0.0040760975937162089, -0.0041994355234903696, 
    -0.0043193331001091864, -0.0044356882411713738, -0.0045483379092283241, 
    -0.0046570426302831747, -0.0047614653340780702, -0.0048611891594383654, 
    -0.0049557301423674262, -0.0050445741829729177, -0.0051272211529425141, 
    -0.0052032235817332743, -0.0052722164014844166, -0.0053339410818367926, 
    -0.0053882542855768845, -0.0054351342282288311, -0.0054746988143650919, 
    -0.0055072110538537901, -0.0055330800492586251, -0.0055528623692443586, 
    -0.0055672476518727762, -0.0055770273651091018, -0.0055830732395433366, 
    -0.0055862891967338396, -0.0055875721636078303, -0.0055877677077251307, 
    -0.0055876375243379718, -0.0055878212780184917, -0.0055888193799679626, 
    -0.0055909748082231927, -0.0055944631358763319, -0.0055992875171550043, 
    -0.005605296036629937, -0.0056121969451662472, -0.0056195900484010816, 
    -0.0056270004329328502, -0.0056339153648809351, -0.0056398031019323468, 
    -0.0056441340062257832, -0.0056463885416236544, -0.0056460514309141915, 
    -0.0056426207372241499, -0.0056356096187100456, -0.0056245548258528509, 
    -0.0056090286027650569, -0.0055886537520946711, -0.0055631274756742146, 
    -0.0055322348080967176, -0.0054958810185302513, -0.0054541095581317322, 
    -0.0054071199085189876, -0.0053552704135947857, -0.0052990762161906017, 
    -0.0052391813680666066, -0.0051763327729119216, -0.0051113430704589711, 
    -0.0050450446950981772, -0.00497825657591245, -0.0049117511593230754, 
    -0.0048462239088773833, -0.0047822792123584455, -0.0047204278019455839, 
    -0.0046610864274810818, -0.0046045880090003367, -0.0045511970548604173, 
    -0.0045011142176016395, -0.0044544945766748605, -0.0044114389656633116, 
    -0.0043720066943202665, -0.0043362189750026005, -0.0043040764664739354, 
    -0.0042755739923088084, -0.0042507261095492644, -0.0042295908597345085, 
    -0.0042122892511027837, -0.0041990190423686988, -0.0041900572423348038, 
    -0.0041857578988913624, -0.0041865410843386335, -0.0041928832843494378, 
    -0.004205292801427311, -0.0042242968667132496, -0.0042504097280632487, 
    -0.0042841104388236162, -0.0043258253032364361, -0.0043758880970463133, 
    -0.0044345309637539264, -0.0045018580333614387, -0.004577833928782471, 
    -0.0046622822136221567, -0.0047548901806979387, -0.004855208673719801, 
    -0.0049626777431256387, -0.0050766292746233631, -0.0051963184134951618, 
    -0.0053209304151504086, -0.0054495967600972899, -0.0055814134041880523, 
    -0.0057154537078700938, -0.0058507782415443835, -0.0059864529403971549, 
    -0.0061215601207373314, -0.006255216943841466, -0.0063865934709749338, 
    -0.0065149243685225251, -0.0066395317272972187, -0.0067598271497199981, 
    -0.0068753083275469055, -0.0069855515346723294, -0.0070901778237646611, 
    -0.0071888338061131957, -0.0072811727181740175, -0.0073668386453895913, 
    -0.0074454670961679086, -0.0075166875740987184, -0.0075801440432201285, 
    -0.0076355033357996252, -0.0076824875150379255, -0.0077208891942394655, 
    -0.0077506034958473233, -0.0077716260801820479, -0.0077840604964748471, 
    -0.0077881083398150487, -0.0077840519187840542, -0.0077722303418170892, 
    -0.0077530202003454531, -0.0077268205510625954, -0.0076940399099031448, 
    -0.0076551049994377967, -0.007610454045313372, -0.0075605641147013479, 
    -0.0075059600152347179, -0.0074472400215323158, -0.0073850791530269064, 
    -0.0073202377901693989, -0.0072535388164067854, -0.0071858557227391694, 
    -0.0071180849876901252, -0.0070511039522884915, -0.0069857510029698129, 
    -0.0069227789786981053, -0.0068628377990997786, -0.0068064394212342672, 
    -0.0067539482474123051, -0.0067055743367002195, -0.0066613762872651501, 
    -0.0066212700719555243, -0.0065850530941906453, -0.0065524193214370335, 
    -0.0065229880235470701, -0.0064963217674293538, -0.0064719512838035736, 
    -0.0064494031501501252, -0.0064282361458038728, -0.0064080822889971039, 
    -0.0063886838295297062, -0.0063699201051918963, -0.0063518175550802674, 
    -0.0063345196351848269, -0.0063182519584643439, -0.0063032649625731274, 
    -0.006289785852504913, -0.0062779761960957232, -0.0062678912767211784, 
    -0.0062594681549962734, -0.0062525137533513929, -0.006246709428584166, 
    -0.0062416245091101805, -0.0062367362645543798, -0.0062314493261666441, 
    -0.0062251186860081253, -0.0062170838763835664, -0.0062066778862657612, 
    -0.0061932473488399654, -0.0061761591108206249, -0.0061548113979157711, 
    -0.0061286350438245684, -0.0060971034536137173, -0.0060597422202137647, 
    -0.006016152778012292, -0.0059660320979874303, -0.0059091951164216214, 
    -0.0058455900318919052, -0.005775299560981037, -0.0056985404740100181, 
    -0.0056156499057260188, -0.0055270624377213697, -0.0054332945927274851, 
    -0.0053349214967213458, -0.0052325707837029738, -0.0051269255482860199, 
    -0.0050187227644079109, -0.0049087659195910247, -0.0047979321011285669, 
    -0.0046871708668502193, -0.0045774836638157613, -0.0044698954571497345, 
    -0.0043654160103236703, -0.0042650017413498617, -0.004169513336224972, 
    -0.0040796809446311012, -0.0039960782078848796, -0.0039191125856117273, 
    -0.0038490212443079578, -0.0037858911333724567, -0.0037296697381604335, 
    -0.0036801986461583395, -0.0036372290959168201, -0.0036004425907011032, 
    -0.0035694659871458147, -0.003543865444854878, -0.0035231439404577606, 
    -0.0035067408670563056, -0.0034940197673703302, -0.0034842692835144956, 
    -0.0034767169493062073, -0.0034705235328582511, -0.0034647963414480326, 
    -0.0034585941631041098, -0.003450927900856438, -0.0034407635799743493, 
    -0.0034270449169730142, -0.0034086999162138607, -0.0033846526203380163, 
    -0.0033538442456403353, -0.0033152361847376688, -0.0032678202838754547, 
    -0.0032106313759868279, -0.0031427655298602321, -0.0030634224845402453, 
    -0.00297192958980855, -0.0028677939613997211, -0.0027507298162174013, 
    -0.0026206848986258979, -0.0024778603070951099, -0.0023227067764953571, 
    -0.0021559082145603549, -0.0019783683754150821, -0.0017911627513995652, 
    -0.0015955175038262384, -0.0013927539774866776, -0.0011842445107631283, 
    -0.00097137343205587934, -0.00075548946721578822, 
    -0.00053788933304317957, -0.00031979758558619453, -0.000102368549095301, 
    0.0001133009048179649, 0.00032616429539540637, 0.00053519943872649229, 
    0.00073941949638523256, 0.00093786382366790812, 0.0011296114813072419, 
    0.0013138005271166632, 0.0014896404105298948, 0.0016564288218070744, 
    0.0018135585155933879, 0.0019605415255262242, 0.0020970070177222869, 
    0.0022227092540985384, 0.0023375453940000148, 0.0024415277128259404, 
    0.0025347864579045409, 0.0026175553265153305, 0.0026901302252861619, 
    0.0027528354262025679, 0.0028059843602352775, 0.0028498407609973226, 
    0.0028845756899858657, 0.0029102343765888159, 0.0029267197459687481, 
    0.0029337564216188731, 0.0029308988861377503, 0.0029175226487870693, 
    0.0028928429541192247, 0.0028559367788576584, 0.0028057846981754926, 
    0.002741321502952703, 0.0026614857674529058, 0.0025652761014933931, 
    0.0024518188897652096, 0.002320409688558765, 0.0021705429998500041, 
    0.002001974708072919, 0.0018147347948791715, 0.0016091793143922632, 
    0.0013860218730721476, 0.0011463523523276517, 0.00089168097290241873, 
    0.0006239481142310525, 0.00034554334085618813, 5.9305978197923001e-05, 
    -0.00023150598334278894, -0.00052332406366706948, 
    -0.00081238479256268592, -0.0010949676163314703, -0.0013675921902807811, 
    -0.0016271898060939507, -0.0018712119830320176, -0.0020976656127120728, 
    -0.0023050877826566859, -0.0024925007248982707, -0.0026593481926854082, 
    -0.0028054374492916608, -0.0029308686294820252, -0.0030359882192813811, 
    -0.003121332632549322, -0.0031876230431166276, -0.0032357139632609344, 
    -0.0032666164480857586, -0.0032814688070904883, -0.0032815278056362567, 
    -0.0032681277807701304, -0.0032426439957250956, -0.0032064478169623791, 
    -0.0031608584599224841, -0.0031071465060184024, -0.0030465187448986105, 
    -0.002980153426547733, -0.0029092402126259216, -0.0028350060610087399, 
    -0.0027587437513732983, -0.0026818118700546916, -0.0026056109803353051, 
    -0.0025315746128803766, -0.0024611220020206845, -0.0023956540782384991, 
    -0.0023365135950355869, -0.0022849444296177681, -0.0022420823264071156, 
    -0.0022089079908175551, -0.0021862353197761092, -0.0021746776366824015, 
    -0.0021746451352926098, -0.0021863597671150444, -0.0022098543366286679, 
    -0.0022450186500619848, -0.0022916350253081282, -0.0023494339154822123, 
    -0.0024181480369184823, -0.0024975597228156354, -0.0025875492204194173, 
    -0.0026880889838166526, -0.0027992137425110909, -0.0029210102997245433, 
    -0.0030535315201085894, -0.0031967929719798806, -0.0033507142816622958, 
    -0.0035151348654920474, -0.0036897846572793865, -0.0038743005336922005, 
    -0.0040682573080235906, -0.0042711659699067976, -0.004482519132355531, 
    -0.0047017894381811776, -0.0049284665313616355, -0.0051620562155467549, 
    -0.0054020948015033009, -0.0056481359044819679, -0.0058997146451354853, 
    -0.006156296077854383, -0.0064172468448250447, -0.0066817632769042975, 
    -0.0069488211095641928, -0.0072171441365798871, -0.0074852041015572102, 
    -0.0077512414955731614, -0.0080133105289066971, -0.0082693416714755066, 
    -0.0085171896101788568, -0.0087546542087461598, -0.0089795017172113294, 
    -0.0091894560773890244, -0.0093821623549991771, -0.0095551970784189828, 
    -0.0097060741680782027, -0.0098322774311703706, -0.0099313125966973385, 
    -0.010000781669182602, -0.010038453609592837, -0.010042365381873712, 
    -0.010010866832618011, -0.0099426967240144881, -0.009837062994654637, 
    -0.0096936684324388962, -0.0095128128534441962, -0.0092954171451344776, 
    -0.0090430989830053102, -0.0087581985635052581, -0.0084438180786581517, 
    -0.0081038435301544042, -0.0077428742663446098, -0.0073662114295159377, 
    -0.0069797237915283222, -0.0065897284292771446, -0.0062028189023100736, 
    -0.0058256991243889108, -0.0054650709528812364, -0.0051274497317671634, 
    -0.0048190314957873969, -0.004545587024189118, -0.0043123249562318239, 
    -0.0041237859914260303, -0.0039837796500085416, -0.0038952573758940694, 
    -0.0038603131119386118, -0.0038800924556783656, -0.0039548174598263664, 
    -0.0040837540330193774, -0.0042652596888688183, -0.0044967624520198674, 
    -0.0047747897163219009, -0.0050949593064622545, -0.0054520633584610014, 
    -0.0058400841526172354, -0.0062522531976854454, -0.0066811671980403437, 
    -0.0071188606604538586, -0.0075570532677994105, -0.0079872958128049971, 
    -0.0084012719322968769, -0.008790981981839174, -0.0091490902201012969, 
    -0.0094690596301069494, -0.0097454468032648223, -0.0099739673281124801, 
    -0.010151673805086376, -0.010277067322474485, -0.010350102070487279, 
    -0.010372175886370242, -0.010346050825485308, -0.010275744094552678, 
    -0.01016641202222463, -0.010024022439508746, -0.0098551725523853256, 
    -0.0096667195249149594, -0.0094654220837936068, -0.0092576724911452163, 
    -0.0090494275814509192, -0.0088461304704607422, -0.0086527342456397954, 
    -0.0084737763793303056, -0.0083130452502616255, -0.0081735935125854843, 
    -0.0080572932871869687, -0.0079649304618234166, -0.0078959633580688374, 
    -0.0078487178672614778, -0.0078205854507964381, -0.0078081181376425642, 
    -0.0078074347098812946, -0.0078143208704164538, -0.0078250677226508365, 
    -0.0078361750748916336, -0.0078454795774851611, -0.0078518918219181756, 
    -0.0078561457885194946, -0.007860370620537226, -0.0078694102604162687, 
    -0.0078893839999277619,
  // Fqt-Na(3, 0-1999)
    1, 0.99846482694426086, 0.9938827389734467, 0.9863229989511253, 
    0.97589820359091062, 0.96276042697130748, 0.94709618373548377, 
    0.92912053315927645, 0.90907064736150378, 0.88719917774416068, 
    0.8637677257361146, 0.83904066686042111, 0.81327953445488843, 
    0.78673810883253026, 0.75965829145817332, 0.73226680236255481, 
    0.70477268883701483, 0.67736561628162129, 0.65021484787537542, 
    0.62346886239467414, 0.59725549926865507, 0.57168255032140036, 
    0.5468387065497734, 0.52279476007050085, 0.499605002026556, 
    0.47730871558309446, 0.45593172865474957, 0.43548797501634312, 
    0.41598102100722795, 0.39740553341768814, 0.37974867635663112, 
    0.36299139755362192, 0.34710962037786963, 0.33207530775194116, 
    0.3178574094996699, 0.30442268539268186, 0.29173641439692716, 
    0.27976299647220881, 0.2684664530067678, 0.25781085036082441, 
    0.24776064160769573, 0.2382809573998558, 0.22933783564533344, 
    0.2208984192451583, 0.21293110106974691, 0.20540564285549273, 
    0.19829325632664743, 0.19156665971115044, 0.18520010581384053, 
    0.17916939260620932, 0.17345184329009883, 0.1680262843317927, 
    0.16287300116813241, 0.15797369163070479, 0.15331140487011499, 
    0.148870481692086, 0.14463648904633419, 0.14059614847094945, 
    0.13673726788488696, 0.1330486775918571, 0.12952015255535054, 
    0.12614234395945439, 0.12290671087329594, 0.11980543656326806, 
    0.11683134752978153, 0.11397782078934582, 0.11123868453765332, 
    0.10860812780473504, 0.10608060746202826, 0.10365077817107632, 
    0.10131344162978577, 0.099063509474687617, 0.096895989494831247, 
    0.094805979020700024, 0.092788673935982682, 0.090839381445768724, 
    0.088953533919489111, 0.087126707314729226, 0.085354634092288051, 
    0.083633225367916092, 0.081958578001260454, 0.080326995217229163, 
    0.078734997428138248, 0.077179341527736839, 0.075657035607005041, 
    0.074165358335909329, 0.072701875202589861, 0.071264457541105414, 
    0.069851293816424131, 0.068460889013745238, 0.067092072367935726, 
    0.065743989418299675, 0.064416097534579608, 0.063108159225626834, 
    0.061820230156955189, 0.060552649554747949, 0.059306012157169526, 
    0.058081138349515879, 0.056879027025522229, 0.055700811421359839, 
    0.054547707771276911, 0.053420967491777979, 0.052321832656368153, 
    0.051251497422623929, 0.050211079487508109, 0.049201592550199069, 
    0.048223929946149817, 0.047278848686170195, 0.0463669678167382, 
    0.045488762628402353, 0.044644568775236149, 0.043834587357260507, 
    0.043058893772126128, 0.042317440661409057, 0.041610066667071087, 
    0.040936498642944401, 0.040296349264969285, 0.039689114989088281, 
    0.039114176406989901, 0.038570803438297496, 0.038058157242377641, 
    0.037575302786221544, 0.037121213663086149, 0.036694787697223591, 
    0.036294848983017526, 0.035920153652419975, 0.035569390580181159, 
    0.035241176706025779, 0.034934055748322014, 0.034646492332888336, 
    0.034376870249500098, 0.034123503673313245, 0.033884639777676431, 
    0.03365846879245591, 0.033443133636859315, 0.033236745193777013, 
    0.03303739447349209, 0.032843175828835558, 0.032652212267727063, 
    0.032462686978929886, 0.032272875504260785, 0.032081180937883515, 
    0.031886162097418444, 0.031686557797913691, 0.031481302863850563, 
    0.031269530647317696, 0.031050577580784791, 0.030823970643597161, 
    0.03058941611361992, 0.030346784422139957, 0.0300960942341372, 
    0.029837488820274188, 0.029571224634655394, 0.029297644757682074, 
    0.029017163547486201, 0.028730248350321615, 0.028437398524797531, 
    0.028139134977574386, 0.027835989173296098, 0.027528505947881067, 
    0.027217244990451993, 0.026902798250508224, 0.026585799252977223, 
    0.026266935880112134, 0.025946952244195198, 0.025626648250398416, 
    0.025306861021172879, 0.024988440368928565, 0.024672223213255427, 
    0.024358998952957581, 0.024049487135700352, 0.023744319861190504, 
    0.023444031724741608, 0.023149047816453112, 0.02285968030945059, 
    0.022576124819805678, 0.022298461238164702, 0.022026654301735921, 
    0.021760555074465768, 0.021499907396677249, 0.021244350295534252, 
    0.020993430739131874, 0.020746610830941051, 0.020503296629148321, 
    0.020262853184996692, 0.020024641835354899, 0.019788048029414331, 
    0.019552514539922565, 0.019317576259193888, 0.019082892944232547, 
    0.018848278003996632, 0.018613727884059954, 0.018379438726103398, 
    0.018145811390546648, 0.017913444798938496, 0.017683112345159478, 
    0.017455730089751879, 0.017232318510250373, 0.017013952505228139, 
    0.016801716670888985, 0.016596655317511155, 0.016399732933436599, 
    0.016211789366528378, 0.016033510534767297, 0.015865401155254651, 
    0.015707767775882012, 0.015560708632276014, 0.015424112823698885, 
    0.015297665788967038, 0.015180860919010259, 0.015073016204735062, 
    0.014973295037168891, 0.014880733383104607, 0.01479426568925769, 
    0.014712752304266493, 0.014635011302179608, 0.014559844463820382, 
    0.014486065645683508, 0.014412519669464522, 0.014338103836263666, 
    0.014261779484292027, 0.014182587649969377, 0.014099656683379213, 
    0.014012213632212072, 0.013919592651040842, 0.013821245484699636, 
    0.013716745008816712, 0.013605797191476086, 0.013488239708018088, 
    0.01336404214545397, 0.013233311579415354, 0.013096280342697567, 
    0.012953302692975602, 0.012804845646429072, 0.012651475117982687, 
    0.01249384214003354, 0.01233266270656206, 0.012168702998073429, 
    0.012002755794880133, 0.011835622620156638, 0.011668094877177975, 
    0.011500936755529035, 0.011334870861251222, 0.011170568804987633, 
    0.011008647685822506, 0.01084966412373814, 0.010694115104864782, 
    0.010542435982083674, 0.010395000767595208, 0.010252125279308655, 
    0.010114064665845137, 0.0099810233328042394, 0.0098531617529019275, 
    0.0097306007597145975, 0.009613439661652087, 0.009501768991345012, 
    0.0093956856130004048, 0.0092953185286603172, 0.0092008444125694522, 
    0.0091125006260112332, 0.0090305969366944339, 0.0089555153855737975, 
    0.0088877045476873171, 0.0088276611554927061, 0.0087759062304921254, 
    0.0087329628369139742, 0.0086993233755650289, 0.0086754324025292047, 
    0.0086616598417842208, 0.0086582924525852329, 0.0086655240384455774, 
    0.008683450059141418, 0.0087120719863352618, 0.0087512976624262336, 
    0.0088009563789853661, 0.00886080891639646, 0.0089305639086198728, 
    0.0090098951780847591, 0.0090984561124017559, 0.0091958935337207968, 
    0.0093018579147714445, 0.0094160050171805711, 0.0095379961444493795, 
    0.0096674925122093164, 0.0098041493986192867, 0.0099476056192556207, 
    0.01009747003765077, 0.010253308606055103, 0.01041462640235777, 
    0.010580855920837734, 0.010751329841897649, 0.010925273452036536, 
    0.011101780216053724, 0.011279809400876603, 0.011458181841403629, 
    0.011635583808333013, 0.011810579156483201, 0.011981626827642797, 
    0.012147100388229738, 0.012305311031542417, 0.01245452767480114, 
    0.012592995433077431, 0.012718953017955482, 0.012830654077224763, 
    0.012926381015982154, 0.01300446466249423, 0.013063298196618651, 
    0.013101353659934733, 0.013117190287831714, 0.01310946916481916, 
    0.013076957723975564, 0.013018540600437157, 0.012933232334234504, 
    0.01282019768575563, 0.012678775045403535, 0.012508513931374234, 
    0.012309212383344491, 0.012080953001264228, 0.011824135727547922, 
    0.011539503495094637, 0.011228145395417029, 0.010891495868279116, 
    0.010531312868989602, 0.010149646340222312, 0.0097487932790849222, 
    0.0093312460304532819, 0.0088996392284977494, 0.0084566982976193028, 
    0.0080051878174466091, 0.0075478721222176125, 0.0070874805584756305, 
    0.0066266873084598575, 0.0061680972097269337, 0.0057142397492369627, 
    0.0052675692113128489, 0.004830464991071151, 0.0044052247384603581, 
    0.0039940505495951479, 0.0035990375968426584, 0.0032221456079574973, 
    0.0028651754856786958, 0.0025297447587149481, 0.0022172667008663501, 
    0.0019289387584066192, 0.001665726557131343, 0.001428358005827706, 
    0.0012173133477426821, 0.0010328143449223029, 0.00087481804121276223, 
    0.00074300663486786297, 0.00063678726150902623, 0.00055529118265573068, 
    0.0004973930667049205, 0.00046173317603011424, 0.00044675981667685702, 
    0.00045077359136672237, 0.0004719831403249597, 0.00050855617193069794, 
    0.00055866746730884483, 0.00062053791289336257, 0.00069246664465563192, 
    0.00077285168443557274, 0.00086020621122780204, 0.00095316328631639478, 
    0.0010504830849284532, 0.0011510505139903306, 0.001253878148500865, 
    0.0013581081379481943, 0.0014630151415566325, 0.0015680113265146693, 
    0.001672648499368423, 0.0017766222977392979, 0.0018797683241598714, 
    0.0019820623479046475, 0.0020836105714616302, 0.0021846359247911255, 
    0.0022854676668117501, 0.0023865229816742426, 0.0024882907394504243, 
    0.0025913193243358836, 0.0026962013264833651, 0.0028035569975536556, 
    0.0029140219219333501, 0.003028219579287005, 0.0031467471037613429, 
    0.0032701490585909905, 0.0033988969427270407, 0.0035333684697578583, 
    0.0036738310322193429, 0.0038204280075809149, 0.0039731725265176347, 
    0.0041319427018872111, 0.0042964782911363965, 0.0044663862205433988, 
    0.0046411403742174385, 0.0048200884181435703, 0.0050024612376259681, 
    0.0051873814227860679, 0.0053738827301436061, 0.0055609179855315863, 
    0.0057473767705974125, 0.0059321021580973467, 0.0061139026121728862, 
    0.0062915634532112359, 0.0064638573569906392, 0.0066295530836343085, 
    0.0067874202177596451, 0.006936235493254032, 0.0070747927320239847, 
    0.0072019128126439699, 0.0073164541341719739, 0.0074173317915860147, 
    0.0075035376938692219, 0.0075741668130560463, 0.0076284422539838704, 
    0.007665738792041822, 0.0076855962846785883, 0.0076877337086237382, 
    0.0076720448908386982, 0.0076385940517656016, 0.0075876075540234622, 
    0.00751946514124329, 0.0074346988869894454, 0.0073339916117494703, 
    0.0072181809642924127, 0.0070882659470135482, 0.0069454135611056811, 
    0.0067909643749590239, 0.0066264293797820683, 0.0064534836919925053, 
    0.0062739532325685873, 0.0060897920583245302, 0.0059030604026529517, 
    0.0057158974385907863, 0.0055304884404164048, 0.0053490246428518498, 
    0.0051736619180707318, 0.0050064731864746951, 0.0048494037378575203, 
    0.0047042261448620361, 0.0045725052689599829, 0.0044555725353641797, 
    0.0043545052601202767, 0.0042701172283974463, 0.0042029612301611235, 
    0.00415332880714588, 0.0041212651286815088, 0.0041065802413987936, 
    0.0041088652570979442, 0.0041275068076790699, 0.0041617050607539122, 
    0.0042104880196956506, 0.0042727248215074778, 0.0043471416779711867, 
    0.004432345270213793, 0.0045268508461762903, 0.0046291167112119443, 
    0.0047375842249026004, 0.0048507185333955365, 0.0049670376175257706, 
    0.0050851456700816049, 0.005203751293306717, 0.0053216779374516479, 
    0.0054378721154908424, 0.005551403315217307, 0.0056614655181851372, 
    0.0057673750242014325, 0.005868566842461097, 0.0059645912027806447, 
    0.0060551054118542051, 0.0061398677875567926, 0.0062187289042429815, 
    0.00629162324729128, 0.0063585600988165791, 0.0064196192515804011, 
    0.0064749522792028882, 0.0065247750063053443, 0.0065693740146137254, 
    0.0066091016570623291, 0.0066443729955770522, 0.0066756589057831448, 
    0.0067034810494558204, 0.0067283945621529374, 0.0067509745336180255, 
    0.0067717963627597424, 0.0067914117538886275, 0.0068103169272790941, 
    0.0068289250406163293, 0.0068475332581629774, 0.0068662933995742919, 
    0.006885191577778919, 0.0069040345390172404, 0.0069224489941588736, 
    0.0069398995578537574, 0.0069557109523258895, 0.0069691036002816151, 
    0.0069792235189781631, 0.00698517539084457, 0.0069860481131174147, 
    0.0069809353457922331, 0.0069689504388714789, 0.0069492420047435116, 
    0.0069210078181783643, 0.006883518832578735, 0.0068361373738661428, 
    0.0067783507140749405, 0.0067097969221974682, 0.0066302913210252784, 
    0.0065398458221668735, 0.0064386837639754321, 0.0063272498187487113, 
    0.0062062167006949887, 0.0060764864018724692, 0.0059391862591859062, 
    0.005795662947373768, 0.0056474636041261598, 0.0054963134780385437, 
    0.0053440806509711721, 0.0051927429878948477, 0.0050443438112664192, 
    0.0049009477606778507, 0.0047646001232948794, 0.0046372799112202757, 
    0.0045208581662045666, 0.0044170583418858588, 0.0043274223036008719, 
    0.0042532822313449473, 0.0041957437701969375, 0.0041556674922750975, 
    0.004133664495552085, 0.0041300868108391994, 0.0041450202656992891, 
    0.0041782808343284392, 0.00422941269215487, 0.0042976896582931053, 
    0.0043821190295042847, 0.004481448726700938, 0.0045941803338845431, 
    0.0047185861384834386, 0.00485274056174443, 0.0049945598042340188, 
    0.00514185866308676, 0.0052924090386890187, 0.0054440101817756397, 
    0.0055945548313119505, 0.0057420906340587934, 0.0058848698315257684, 
    0.0060213870058484706, 0.006150404807391676, 0.0062709644699445247, 
    0.0063823900675911835, 0.0064842779732012679, 0.0065764832872661468, 
    0.0066591033127456241, 0.0067324524873721651, 0.006797035677557824, 
    0.0068535186208633758, 0.0069026925951926697, 0.0069454367485725296, 
    0.006982681201668884, 0.0070153717325921686, 0.007044435717643298, 
    0.0070707569800873438, 0.007095150307614739, 0.0071183418668934809, 
    0.0071409574913882763, 0.0071635165003526291, 0.0071864293168806027, 
    0.0072100078019143449, 0.0072344652078855038, 0.0072599284178417427, 
    0.0072864472551180653, 0.007314008233705138, 0.0073425473562546383, 
    0.0073719658855176213, 0.0074021439688921799, 0.0074329597478478377, 
    0.0074642999214780126, 0.0074960731673325435, 0.0075282155025305983, 
    0.0075607042344496035, 0.0075935565648847332, 0.0076268289726979504, 
    0.0076606085521122736, 0.0076950053461026912, 0.0077301316584448988, 
    0.0077660813400871904, 0.0078029007490451729, 0.0078405697666735167, 
    0.0078789809701186909, 0.0079179176027970224, 0.0079570558041559287, 
    0.0079959569892461141, 0.0080340807858281845, 0.0080707997891200211, 
    0.0081054269663061295, 0.0081372420108015223, 0.0081655224874578013, 
    0.0081895699519807241, 0.0082087275888030158, 0.0082223927488526728, 
    0.0082300203932702577, 0.0082311239105141848, 0.0082252677052092275, 
    0.008212060498932177, 0.0081911489352345344, 0.0081622110051223183, 
    0.0081249546431197226, 0.0080791190220737483, 0.0080244810065105195, 
    0.0079608670580150042, 0.0078881662583906321, 0.0078063467235873736, 
    0.0077154739999756895, 0.0076157224095203075, 0.0075073900455159851, 
    0.0073909010505824576, 0.0072668040991532828, 0.0071357659007788244, 
    0.0069985500693455268, 0.0068559980544229951, 0.0067090044351921056, 
    0.0065584898059252205, 0.0064053761847373963, 0.0062505625256641158, 
    0.0060949048873627943, 0.005939198697887978, 0.0057841687736374268, 
    0.005630456560746358, 0.0054786225555457499, 0.0053291482837259842, 
    0.005182441452178662, 0.0050388503128181153, 0.0048986753837095675, 
    0.0047621884689128544, 0.0046296499253810639, 0.0045013267595900453, 
    0.0043775088953381504, 0.0042585159137215178, 0.0041447010860446208, 
    0.0040364419386518611, 0.0039341307109682791, 0.0038381477683679015, 
    0.0037488441698602729, 0.0036665193823399046, 0.0035914086331159181, 
    0.0035236786548234183, 0.0034634256001372502, 0.0034106847254072353, 
    0.0033654366908328461, 0.0033276176459553597, 0.0032971256910771332, 
    0.0032738309585893391, 0.0032575757055106785, 0.0032481805485030956, 
    0.0032454430653100067, 0.0032491326492181641, 0.0032589867443618315, 
    0.0032747015216186013, 0.0032959154712536498, 0.0033221940965091692, 
    0.0033530171272593543, 0.0033877722542903026, 0.003425761952862275, 
    0.0034662236728191841, 0.0035083588773861143, 0.0035513755099099041, 
    0.0035945260615830471, 0.0036371451941391887, 0.0036786805869313492, 
    0.0037187058398326211, 0.0037569280718359535, 0.0037931722506287539, 
    0.0038273719399338096, 0.0038595389651224282, 0.0038897421308035402, 
    0.0039180787546864706, 0.0039446539367440523, 0.0039695565042504538, 
    0.0039928406017745981, 0.0040145069373537304, 0.0040344949884233289, 
    0.0040526723553119502, 0.0040688479582609615, 0.004082779881005633, 
    0.0040941968967642389, 0.0041028242919416476, 0.0041084076446512288, 
    0.0041107303696200836, 0.0041096266328744645, 0.0041049799159644344, 
    0.004096724062922821, 0.0040848323195011799, 0.0040693033757938837, 
    0.0040501506181255947, 0.0040273842560914598, 0.0040009959104806859, 
    0.003970934141715403, 0.0039370759845339578, 0.0038992116474378725, 
    0.0038570197801946768, 0.0038100628397811959, 0.0037577948153044642, 
    0.0036995728727066057, 0.0036346872075497436, 0.0035623875433192747, 
    0.00348192114618554, 0.0033925650653045432, 0.0032936599341637789, 
    0.0031846349880111985, 0.0030650350243476825, 0.0029345373636601004, 
    0.0027929602793506053, 0.0026402764325071534, 0.0024766047462783224, 
    0.0023022126649509889, 0.0021175004763195776, 0.0019229912310625861, 
    0.0017193135829948508, 0.001507184591234069, 0.0012873915599746798, 
    0.0010607755911090236, 0.00082821663920441715, 0.00059062176752924106, 
    0.00034892047534918191, 0.00010406468160220817, -0.00014296771402030743, 
    -0.0003911618064571644, -0.00063945680320420914, -0.00088673588992662451, 
    -0.0011318232027049252, -0.0013734825690520087, -0.0016104224851985645, 
    -0.0018413127540474015, -0.0020648015241357346, -0.002279536418787525, 
    -0.0024841848385178875, -0.0026774555330952719, -0.0028581184380080996, 
    -0.0030250227652304381, -0.0031771174390194568, -0.003313476676245204, 
    -0.0034333259827876348, -0.0035360684167934989, -0.003621316673802286, 
    -0.0036889128225551572, -0.0037389449426619439, -0.0037717466351534219, 
    -0.0037878882165085408, -0.0037881466218576609, -0.0037734785102786239, 
    -0.0037449812027414149, -0.0037038569653618436, -0.0036513838051121564, 
    -0.0035888828019110205, -0.0035177045817896785, -0.0034392035413907513, 
    -0.0033547265179169846, -0.0032655996392673471, -0.0031731129157531587, 
    -0.0030785119623534299, -0.0029829857819162536, -0.0028876642547367047, 
    -0.0027936087120169002, -0.002701814181977544, -0.0026132001155697729, 
    -0.0025286128120375786, -0.0024488184176428688, -0.0023745013749883106, 
    -0.0023062607612600976, -0.0022446096013605146, -0.0021899681619420843, 
    -0.0021426654390768762, -0.0021029411135077315, -0.0020709464122859417, 
    -0.0020467562760202477, -0.0020303744788629325, -0.0020217480445441846, 
    -0.0020207725767578994, -0.0020273034649034316, -0.0020411609670251411, 
    -0.0020621379965010418, -0.0020899971618543976, -0.0021244737659139867, 
    -0.0021652749340551869, -0.0022120762519719072, -0.0022645220281832432, 
    -0.0023222220901553802, -0.0023847484120896028, -0.0024516413311098792, 
    -0.0025224021617503479, -0.0025964994419242805, -0.0026733652073232762, 
    -0.0027524036939676204, -0.0028329890262522852, -0.0029144789677661956, 
    -0.0029962188638850197, -0.0030775541053517643, -0.0031578385151974702, 
    -0.0032364439874250847, -0.0033127680947563371, -0.0033862441375216729, 
    -0.003456350180159851, -0.0035226236558077713, -0.0035846699340371349, 
    -0.0036421778937131485, -0.0036949280741625768, -0.0037427986215346808, 
    -0.0037857702064817882, -0.0038239229734599867, -0.0038574297258544103, 
    -0.0038865458348982525, -0.0039116009754168943, -0.0039329883173656816, 
    -0.0039511555910039181, -0.0039665976194722058, -0.0039798470260838078, 
    -0.0039914648004283834, -0.0040020266287950556, -0.0040121153279208694, 
    -0.0040222961652524999, -0.004033103291063149, -0.0040450203835977402, 
    -0.0040584561208605111, -0.004073724332407898, -0.0040910245121970508, 
    -0.0041104258348987465, -0.0041318592602364208, -0.0041551127072955649, 
    -0.004179830569728489, -0.0042055257353760134, -0.0042315832105495116, 
    -0.0042572779429131099, -0.0042817859000102917, -0.0043042001710440403, 
    -0.0043235435719440165, -0.0043387874340098075, -0.004348869502436516, 
    -0.0043527190011577949, -0.0043492839974667921, -0.0043375629292731381, 
    -0.0043166391434084758, -0.0042857174427245607, -0.0042441562019010677, 
    -0.0041915025765887556, -0.0041275120449626879, -0.004052170437965982, 
    -0.0039657060252814369, -0.0038685882124283011, -0.0037615229477399783, 
    -0.0036454384010227805, -0.0035214641007920611, -0.0033909066902084238, 
    -0.0032552179963432175, -0.0031159595979590826, -0.0029747764028648666, 
    -0.0028333534381508826, -0.0026933796555962852, -0.0025565083166381318, 
    -0.0024243078314299025, -0.0022982210283595101, -0.0021795168513834727, 
    -0.0020692490117426576, -0.0019682193665543114, -0.0018769463320722822, 
    -0.0017956460623780302, -0.0017242317775197386, -0.0016623155460560339, 
    -0.0016092329322045711, -0.0015640731481184166, -0.0015257221988106149, 
    -0.0014929155310103826, -0.0014642873840262317, -0.0014384204760047922, 
    -0.0014138932740400474, -0.001389317140737851, -0.0013633635692199028, 
    -0.0013347844058717953, -0.0013024222889025591, -0.0012652146663203168, 
    -0.0012221937414921985, -0.0011724805980817031, -0.0011152802465167102, 
    -0.0010498761408226018, -0.00097562554603044106, -0.00089196170755503207, 
    -0.00079839348357120174, -0.0006945107847990071, -0.00057999486196331509, 
    -0.00045462488866474806, -0.00031828590927998336, 
    -0.00017097980476434683, -1.2830762284515116e-05, 0.00015590912658866406, 
    0.00033485672196066044, 0.00052349910255181271, 0.0007211944844304481, 
    0.00092718091879964856, 0.00114057722638165, 0.0013603974080668895, 
    0.001585555520485961, 0.0018148746389904653, 0.0020470942292526153, 
    0.0022808790020890247, 0.0025148277287338617, 0.0027474934405274667, 
    0.0029774005700431015, 0.0032030721793766094, 0.0034230574195114327, 
    0.0036359546027195464, 0.0038404341812185504, 0.0040352513888642048, 
    0.0042192533335167126, 0.00439138181566949, 0.004550675333850728, 
    0.0046962612148380052, 0.004827350338422411, 0.0049432228125075349, 
    0.0050432137121574783, 0.0051267039555842279, 0.0051931095669041187, 
    0.0052418784357842326, 0.0052724920790089566, 0.0052844744316234999, 
    0.0052773996811930823, 0.0052509010783516122, 0.0052046812827221522, 
    0.0051385153588681537, 0.0050522517056704819, 0.0049458086058394466, 
    0.0048191761960604583, 0.0046724156356261932, 0.0045056685596835573, 
    0.0043191625380990112, 0.0041132303657708492, 0.0038883207377303827, 
    0.0036450212410855977, 0.0033840692267156566, 0.0031063664026880831, 
    0.0028129833767476164, 0.0025051677940853695, 0.002184339005457061, 
    0.0018520836643112519, 0.0015101473667380307, 0.0011604255984452262, 
    0.00080494669376154297, 0.00044585670310545505, 8.5391190546222663e-05, 
    -0.00027415463217585136, -0.00063046158001540877, 
    -0.00098123135532891597, -0.0013242235168355815, -0.001657295168602005, 
    -0.0019784322207930466, -0.0022857859994333844, -0.0025776855059219286, 
    -0.0028526574971672164, -0.0031094291585532707, -0.0033469305961822795, 
    -0.0035642847486479583, -0.0037608008012074519, -0.0039359607573468281, 
    -0.0040893964557663157, -0.0042208767777317888, -0.0043302853995337703, 
    -0.0044175993736374859, -0.0044828753048638077, -0.0045262329130101205, 
    -0.0045478499436077792, -0.0045479536478080819, -0.0045268215159579312, 
    -0.0044847812773632202, -0.0044222121058606588, -0.0043395550785115767, 
    -0.004237324243263561, -0.0041161183096157924, -0.0039766382647541841, 
    -0.0038197064728907829, -0.0036462773994915812, -0.0034574563588773604, 
    -0.0032545109946709857, -0.0030388726714667639, -0.0028121436206525446, 
    -0.0025760852563620888, -0.002332605427033156, -0.0020837374893962479, 
    -0.001831619283052041, -0.0015784644363379804, -0.0013265328755640068, 
    -0.0010780965507708803, -0.0008354059432276247, -0.00060065062552046907, 
    -0.000375923801327989, -0.00016318268140928316, 3.5792139388686126e-05, 
    0.00021942667072965476, 0.00038638500239859905, 0.00053558906954174535, 
    0.0006662304495985811, 0.00077777458312436472, 0.00086995103684452211, 
    0.00094274185781205162, 0.00099636173888634195, 0.001031232567890219, 
    0.0010479627960855973, 0.0010473218615598464, 0.0010302210871758633, 
    0.00099770056818943476, 0.00095091139130546419, 0.00089109893365469468, 
    0.00081957117839802623, 0.00073766818905157986, 0.00064671477018105029, 
    0.00054797639588755965, 0.00044262401883969063, 0.00033170531541184276, 
    0.00021613103606736399, 9.6672515967977232e-05, -2.6028507194024615e-05, 
    -0.00015144426958091785, -0.00027913955215958853, 
    -0.00040875095720045132, -0.00053996452870889869, 
    -0.00067249250487710411, -0.00080605532382645639, 
    -0.00094035862229836233, -0.0010750759084722312, -0.0012098237356489609, 
    -0.0013441488017621403, -0.0014775084233393681, -0.0016092626020941555, 
    -0.0017386689720061094, -0.0018648802778117746, -0.0019869509671978426, 
    -0.0021038476298590315, -0.0022144667557753616, -0.0023176623286835047, 
    -0.0024122706629933722, -0.0024971437247892003, -0.0025711800306192738, 
    -0.0026333507064596161, -0.0026827235037847389, -0.0027184826840684329, 
    -0.0027399435729830875, -0.0027465647600507272, -0.0027379622697088503, 
    -0.0027139177491983073, -0.0026743909006324501, -0.0026195345841218349, 
    -0.0025496953570685599, -0.0024654213381460127, -0.0023674583545093067, 
    -0.0022567388332213685, -0.0021343668472980858, -0.0020015949852450602, 
    -0.0018597922015391143, -0.0017104128229844273, -0.0015549610904376748, 
    -0.0013949598480601378, -0.0012319219500808907, -0.0010673292868020406, 
    -0.00090262094018278571, -0.00073918056321668388, 
    -0.00057833256491517907, -0.00042133576370002423, 
    -0.00026938326841060363, -0.00012359201439294404, 1.5002472607575324e-05, 
    0.00014545521973107557, 0.00026691991244497657, 0.00037865790565621584, 
    0.0004800457979950289, 0.00057058000023262035, 0.00064988249245972649, 
    0.00071770742078713045, 0.00077394255993118108, 0.00081861321572327208, 
    0.00085188438135544767, 0.00087405628392080311, 0.00088556304290902965, 
    0.00088696563035773766, 0.00087894459998670398, 0.00086228590386555138, 
    0.00083786649834205365, 0.00080664091655969496, 0.00076960890810579951, 
    0.00072779367704206034, 0.00068221330804412589, 0.00063385062107167416, 
    0.00058363313259302278, 0.00053241195904841132, 0.00048095491816191755, 
    0.00042993871236403906, 0.00037994742586600826, 0.00033148161475172935, 
    0.00028496511879000732, 0.00024076060252622023, 0.00019919036516356353, 
    0.00016055991894264377, 0.00012518182321504017, 9.339380052384859e-05, 
    6.5570537334169331e-05, 4.2122277360709284e-05, 2.3491770157159125e-05, 
    1.0130344254070847e-05, 2.4753076776168836e-06, 9.1813825400761462e-07, 
    5.7724916861568213e-06, 1.7240370166498085e-05, 3.538302127794197e-05, 
    6.010423768671446e-05, 9.1133899411849492e-05, 0.00012803177080463634, 
    0.00017019531474283425, 0.0002168725050474362, 0.00026718594756824313, 
    0.00032016157510645493, 0.00037475824045890994, 0.00042990176759635177, 
    0.00048452352585521917, 0.00053759473399455672, 0.0005881632295015541, 
    0.00063538257818395848, 0.0006785345348381054, 0.00071705694244459837, 
    0.00075055109591630649, 0.00077879633362603544, 0.00080175254978527414, 
    0.00081956424317929338, 0.00083255769691244327, 0.00084123792568133789, 
    0.00084628234402396336, 0.00084853045469863617, 0.00084896409941225741, 
    0.00084868065072643572, 0.00084886060540102239, 0.00085072901076382336, 
    0.00085550988578224829, 0.00086437772606517808, 0.00087841131743029066, 
    0.00089854266421802824, 0.00092551410376013883, 0.00095984445473151336, 
    0.0010018002389763098, 0.0010513836615987752, 0.0011083228484539698, 
    0.0011720757655304314, 0.0012418396411076962, 0.0013165667093970018, 
    0.0013949854260031363, 0.0014756216717747141, 0.0015568320645957009, 
    0.0016368383299851274, 0.001713764948117993, 0.001785688870606356, 
    0.0018506828776197924, 0.0019068641221019502, 0.0019524425735502476, 
    0.0019857644533761098, 0.0020053501929599327, 0.0020099306624250576, 
    0.0019984746933229009, 0.0019702089861629614, 0.0019246372286841193, 
    0.0018615472147219289, 0.0017810074262139552, 0.0016833623801031229, 
    0.0015692128564117535, 0.0014393930616291839, 0.0012949386984779188, 
    0.0011370536034588136, 0.00096707732115971145, 0.00078644561651510013, 
    0.00059665482207737705, 0.00039922169443338504, 0.00019565018685537586, 
    -1.2607501598947365e-05, -0.00022418082425916083, 
    -0.00043780165323140991, -0.00065232252697102855, -0.0008667169577483006, 
    -0.0010800792037225109, -0.0012916100679925546, -0.0015006040038675545, 
    -0.0017064262299111566, -0.0019084998156724843, -0.0021062950436426253, 
    -0.0022993235245118361, -0.0024871429520522828, -0.0026693611757168411, 
    -0.0028456471099676008, -0.0030157398699258565, -0.0031794590077041046, 
    -0.0033367030512979714, -0.0034874542449183951, -0.0036317737250634013, 
    -0.0037697994395436757, -0.0039017467032707066, -0.0040278997971208283, 
    -0.0041486164607540833, -0.0042643263681404371, -0.0043755275652555582, 
    -0.0044827875453194929, -0.0045867340135440967, -0.004688046382706949, 
    -0.0047874350169660237, -0.0048856244770310196, -0.0049833247799406042, 
    -0.0050812104278506638, -0.0051798968398467857, -0.0052799247262088579, 
    -0.0053817498092135468, -0.0054857365533549432, -0.0055921588847706889, 
    -0.0057011998609001868, -0.0058129559712447928, -0.0059274325290193507, 
    -0.0060445457446829118, -0.0061641137838995682, -0.0062858590038509876, 
    -0.0064093977714671929, -0.0065342449029119941, -0.0066598181796553102, 
    -0.0067854465142285648, -0.0069103851884757218, -0.0070338385091849214, 
    -0.0071549802576378451, -0.0072729799983152635, -0.0073870283038315514, 
    -0.0074963624884290857, -0.0076002803294134879, -0.0076981626572298926, 
    -0.007789486414074444, -0.0078738416944105806, -0.0079509430383272496, 
    -0.0080206469545475566, -0.0080829519474381242, -0.0081380084403304236, 
    -0.0081861084631528226, -0.0082276721476789924, -0.0082632212607715704, 
    -0.0082933516180178583, -0.0083186990774816137, -0.0083399054107042743, 
    -0.008357587991372312, -0.0083723134022763695, -0.008384579031290907, 
    -0.0083947984116298537, -0.0084033006078770931, -0.0084103383701850595, 
    -0.008416114338980922, -0.0084208156216167545, -0.0084246466776278922, 
    -0.0084278626938903457, -0.0084307972296072554, -0.0084338758098452104, 
    -0.0084376233833730416, -0.0084426557767123631, -0.0084496616194341175, 
    -0.0084593643490073218, -0.008472484616017021, -0.0084896915570844226, 
    -0.0085115663155856374, -0.0085385599101471584, -0.0085709671092808921, 
    -0.0086089069504283501, -0.0086523133761848437, -0.0087009254887301553, 
    -0.0087542929247456519, -0.008811779374538007, -0.0088725670936494038, 
    -0.0089356814009202076, -0.009000006696757188, -0.0090643234424496073, 
    -0.0091273457886958537, -0.0091877712562404464, -0.009244327612725145, 
    -0.0092958231713221595, -0.0093411815620804573, -0.0093794746196197588, 
    -0.0094099385662918221, -0.0094319782898107905, -0.0094451682265601165, 
    -0.0094492418958647753, -0.0094440711401953658, -0.0094296530575537114, 
    -0.0094060812125584346, -0.0093735195449135885, -0.0093321608797444708, 
    -0.0092822013189744167, -0.0092238066079770448, -0.0091570817067844115, 
    -0.0090820565405355155, -0.0089986676845019153, -0.0089067555827857473, 
    -0.0088060720185966813, -0.0086962972218366918, -0.0085770609680019295, 
    -0.0084479745045240775, -0.0083086638096892852, -0.0081588004992916904, 
    -0.0079981370520959411, -0.0078265239907633673, -0.0076439314714275043, 
    -0.0074504610475303861, -0.0072463423035352727, -0.0070319289594759395, 
    -0.006807699885928999, -0.0065742436268748806, -0.006332266158238271, 
    -0.006082555817179286, -0.0058259635706069835, -0.00556335405772399, 
    -0.0052955570900238471, -0.0050233273593901437, -0.0047473157828897905, 
    -0.0044680560557595625, -0.0041859622697986735, -0.0039013524646249204, 
    -0.0036144647401257549, -0.0033254787414614194, -0.00303454168059451, 
    -0.0027417884525039269, -0.0024473665090513574, -0.0021514530840261786, 
    -0.0018542887882325256, -0.0015561942229539829, -0.0012576015020954942, 
    -0.00095906729490139635, -0.00066129311794992671, 
    -0.00036513416352228776, -7.1608423110971521e-05, 0.00021811437930696967, 
    0.00050272204772990547, 0.00078078388715685726, 0.0010507781879560917, 
    0.0013111327247213506, 0.0015602550396707797, 0.0017965670061786078, 
    0.0020185224440597777, 0.0022246276421118501, 0.0024134442968235352, 
    0.002583596800040631, 0.0027337677421784851, 0.0028627072116217517, 
    0.002969241304757475, 0.0030522861454349544, 0.0031108629462887494, 
    0.0031441028211336374, 0.0031512606109555404, 0.0031317178963017958, 
    0.0030849837942597473, 0.0030107029388858064, 0.0029086694471970368, 
    0.0027788314269578114, 0.0026213155394235036, 0.0024364370534466434, 
    0.0022247120619325717, 0.0019868634222358745, 0.0017238133240049247, 
    0.0014366795955518706, 0.0011267449969312457, 0.00079544236314421657, 
    0.00044433397055147208, 7.5088337309511875e-05, -0.00031054121423529737, 
    -0.0007107368455115294, -0.0011236257874116008, -0.0015473088076170128, 
    -0.001979879149529463, -0.0024194440450375576, -0.0028641482793860559, 
    -0.0033121883947610556, -0.0037618338947617786, -0.0042114325501888712, 
    -0.0046594203151183455, -0.0051043165085172572, -0.005544714926914174, 
    -0.0059792751470966691, -0.0064067001496302626, -0.006825728528057325, 
    -0.0072351260792785496, -0.0076336841584132573, -0.0080202271797521329, 
    -0.0083936221698044031, -0.0087527892360338075, -0.0090967085129776346, 
    -0.0094244330215040393, -0.0097350942214022157, -0.010027905843117458, 
    -0.010302167093039391, -0.010557262984383515, -0.010792665225483465, 
    -0.011007931448489938, -0.011202709052122679, -0.011376732900715532, 
    -0.011529832064211131, -0.011661929892564215, -0.011773054535025775, 
    -0.011863339138377473, -0.011933030136516018, -0.011982486378311268, 
    -0.012012181848564516, -0.012022699358700187, -0.012014720298945932, 
    -0.011989004533921382, -0.011946363506712661, -0.011887627745217674, 
    -0.011813613201989155, -0.011725087416291823, -0.011622747066376843, 
    -0.011507195278364274, -0.011378927532492256, -0.01123833084177267, 
    -0.011085682145256454, -0.010921160794160988, -0.010744854720834304, 
    -0.010556788788706669, -0.010356942918313055, -0.010145277741647859, 
    -0.0099217662693639637, -0.0096864238309281869, -0.0094393278512433839, 
    -0.0091806518283600053, -0.0089106883752814465, -0.0086298728971072186, 
    -0.0083388044242154735, -0.0080382543160917776, -0.0077291817548578593, 
    -0.0074127353447819835, -0.0070902471661671851, -0.0067632308413169417, 
    -0.0064333655203688521, -0.0061024753391917298, -0.0057725091022802063, 
    -0.0054455057069437759, -0.0051235642191560567, -0.0048088076927417294, 
    -0.0045033405613414037, -0.004209223074975922, -0.0039284370818953073, 
    -0.0036628689578528575, -0.0034142924526273963, -0.0031843630433963559, 
    -0.0029746181987470154, -0.0027864701023607224, -0.0026212097226586493, 
    -0.00247998919463041, -0.0023638130964772665, -0.0022735115582410009, 
    -0.0022097199724928226, -0.0021728549508043061, -0.0021630886481800401, 
    -0.0021803315168245083, -0.0022242180941481893, -0.0022941102697140378, 
    -0.0023891010007050183, -0.0025080392879414663, -0.0026495507315590751, 
    -0.0028120748070957912, -0.0029939045530133698, -0.003193219598985692, 
    -0.0034081246757008423, -0.0036366975790987897, -0.0038770215600467768, 
    -0.0041272403738180155, -0.0043856064550987723, -0.004650520233844403, 
    -0.004920555320310183, -0.0051944738890378908, -0.0054712119672613172, 
    -0.005749856046565519, -0.0060296050812742585, -0.0063097385611405763, 
    -0.0065895807273109227, -0.0068684695748703816, -0.0071457385789094087, 
    -0.0074206869430962089, -0.0076925905161032556, -0.0079606830531577244, 
    -0.0082241645864573002, -0.0084822118307658102, -0.0087339863471132748, 
    -0.0089786574446693752, -0.0092154196399368334, -0.0094435256277641821, 
    -0.0096623059330752919, -0.009871209065571214, -0.01006983079009191, 
    -0.010257939851735587, -0.010435513038378278, -0.010602749507992297, 
    -0.010760071026400949, -0.010908111351483217, -0.011047678159670081, 
    -0.011179708881028406, -0.011305201648382687, -0.011425154458672595, 
    -0.011540506636121273, -0.01165207395772814, -0.01176052519492778, 
    -0.011866356458456769, -0.011969882812556204, -0.012071257846212886, 
    -0.012170491400133506, -0.012267471441177047, -0.012362007277572354, 
    -0.012453829740392965, -0.012542605352464027, -0.012627916283047611, 
    -0.0127092402746508, -0.012785923861211084, -0.012857171027704804, 
    -0.012922025384469241, -0.012979388409228612, -0.013028026726995327, 
    -0.013066591620942772, -0.013093646466994409, -0.013107682052595901, 
    -0.013107139082211668, -0.013090424155096793, -0.013055941766263235, 
    -0.013002129697246846, -0.012927486818858651, -0.012830627004503175, 
    -0.012710330285839143, -0.012565583544802616, -0.01239564654087875, 
    -0.01220008367206294, -0.011978808525810507, -0.011732108906755101, 
    -0.011460668212059778, -0.011165571023149735, -0.010848303866087178, 
    -0.010510733631663532, -0.010155084225901662, -0.0097838941661091156, 
    -0.0093999751972165223, -0.0090063512069180687, -0.008606181468144734, 
    -0.0082026868615041951, -0.0077990360191946455, -0.0073982279640493641, 
    -0.0070029669422930017, -0.0066155387496054426, -0.0062377143660336427, 
    -0.0058706820059960712, -0.0055150493383801201, -0.0051708851206910128, 
    -0.0048378259985061341, -0.0045152230550086483, -0.0042022739252901209, 
    -0.003898159951842737, -0.0036021051786847796, -0.0033134068415954891, 
    -0.0030314241312778055, -0.0027555676560805154, -0.0024852660853409165, 
    -0.0022199505875808148, -0.0019590418676825724, -0.00170195977091521, 
    -0.0014481364919421201, -0.0011970621035696646, -0.00094832169066733432, 
    -0.00070167549993569822, -0.00045709818303710584, 
    -0.00021484124628368104, 2.4561853537147439e-05, 0.00026029411758035577, 
    0.00049129146185309302, 0.00071630522196633592, 0.00093397036213749458, 
    0.0011428825957230421, 0.001341673666228089, 0.001529080267078708, 
    0.0017039951929557625, 0.0018655132321045433, 0.0020129694827949766, 
    0.0021459555399809551, 0.0022643315612464101, 0.0023682234523712022, 
    0.0024580068482604918, 0.0025342848582024847, 0.0025978527156674488, 
    0.0026496569314730955, 0.0026907427025437422, 0.0027222169703087339, 
    0.0027452026397749674, 0.0027607928685475128, 0.0027700332082964685, 
    0.0027739023791027951, 0.0027733052934356831, 0.0027690627432138699, 
    0.0027619181987103957, 0.0027525266645993789, 0.0027414511708076907, 
    0.002729169590045463, 0.0027160684320044638, 0.0027024462107829031, 
    0.0026885267140666948, 0.0026744532974266452, 0.0026602921396751333, 
    0.0026460282143467139, 0.0026315592057906505, 0.0026166863454990825, 
    0.0026011089982786854, 0.0025844159705926896, 0.002566075323955498, 
    0.0025454312998847164, 0.0025216944123971244, 0.0024939507651200303, 
    0.0024611928947024242, 0.0024223890834269702, 0.002376571057668018, 
    0.0023229228148962779, 0.0022608546468353675, 0.0021900581789722046, 
    0.0021105114139048737, 0.002022483884457262, 0.0019265176603177245, 
    0.0018234120356489709, 0.0017141945621982919, 0.0016000869917559334, 
    0.0014824859620759332, 0.0013629067151387712, 0.0012429536093360545, 
    0.001124264149730779, 0.0010084797170312396, 0.00089719582164385424, 
    0.00079194005046169871, 0.00069415795722058094, 0.00060520148414858926, 
    0.00052632223981323705, 0.00045867617045106492, 0.00040330352855528416, 
    0.00036111642422840135, 0.00033288271672913866, 0.00031921080137533203, 
    0.00032053850739402251, 0.00033715044489810461, 0.00036918552734664363, 
    0.00041667995353106339, 0.00047959049720597193, 0.00055782659984588464, 
    0.00065128852521011691, 0.00075987766837972944, 0.00088349100525391485, 
    0.0010220213062088802, 0.0011753015271680114, 0.0013430533286622065, 
    0.0015248326778710549, 0.0017199786977589234, 0.0019275835476584104, 
    0.0021464872807944639, 0.0023752932991168022, 0.0026124118220490363, 
    0.0028561092273859511, 0.0031045715426374692, 0.0033559749050493916, 
    0.0036085444143455479, 0.0038606121977754651, 0.0041106441416554713, 
    0.0043572505922244032, 0.0045991836019579815, 0.0048352951512590763, 
    0.005064513371299372, 0.0052858136502662838, 0.0054981663773067237, 
    0.0057005417441713382, 0.0058919016101529218, 0.0060712104166401144, 
    0.0062374537597153605, 0.0063896518001093734, 0.006526874666364515, 
    0.0066482391458093197, 0.006752915138781207, 0.0068401334991593839, 
    0.0069091732755363726, 0.0069593892688092794, 0.0069902280541970542, 
    0.0070012644385873644, 0.0069922294573419126, 0.0069630529924947903, 
    0.0069138754579476987, 0.0068450593597473471, 0.0067571824721701524, 
    0.0066510212910940421, 0.0065275279640902087, 0.0063877778567760614, 
    0.0062329552223377585, 0.0060643045891673854, 0.0058830971146825173, 
    0.0056905931824514852, 0.0054879897276898038, 0.0052763962441767509, 
    0.0050568105307581927, 0.0048301220520714887, 0.0045971098261069661, 
    0.0043584459765336862, 0.0041147280853973374, 0.0038664878838492955, 
    0.0036142520348003116, 0.0033585843395999306, 0.0031001497616084811, 
    0.0028397930352680933, 0.00257857276632497, 0.0023178272359849856, 
    0.0020591853253991176, 0.0018045978475556544, 0.0015563214442137845, 
    0.0013169050248204666, 0.0010891378587128825, 0.00087598346602237444, 
    0.00068049043698093794, 0.00050568552557924849, 0.00035446977765090878, 
    0.00022949038102293429, 0.00013304312179033916, 6.6977825850978091e-05, 
    3.2626540581764664e-05, 3.0749304523142136e-05, 6.1511825854988794e-05, 
    0.00012446233203963552, 0.00021856171629826241, 0.00034219834636959776, 
    0.00049324901256838727, 0.00066913659693977037, 0.00086690142263147149, 
    0.0010832820242741219, 0.0013148061574942984, 0.0015578680668283031, 
    0.0018088319737939332, 0.0020641337290285182, 0.0023203639385907578, 
    0.0025743483477056106, 0.0028232194097814701, 0.0030644536359234883, 
    0.0032958798955140724, 0.0035156623481313546, 0.0037222474201666625, 
    0.0039143176888331317, 0.0040907171959431513, 0.0042504057148608897, 
    0.0043924229770753746, 0.0045158627055889213, 0.0046198614641474612, 
    0.0047036202307667307, 0.0047663964124891184, 0.0048074999410803064, 
    0.0048262913511407535, 0.0048221587213897257, 0.0047945031324044436, 
    0.0047427373682818333, 0.0046662552219283978, 0.0045644291037423533, 
    0.0044366160025573502, 0.004282157837334947, 0.0041004078361505233, 
    0.0038907740721915137, 0.0036527799553403412, 0.0033861379733344755, 
    0.0030908149405629464, 0.0027670855699055167, 0.0024155792703311422, 
    0.0020373088911989478, 0.0016337003238149096, 0.001206602053772769, 
    0.00075833643821783493, 0.00029170193742395639, -0.00019000455000129572, 
    -0.0006829779735483849, -0.0011829233455161051, -0.001685093845907861, 
    -0.0021843768067771902, -0.002675362519867947, -0.0031524956233429219, 
    -0.0036101850948510837, -0.0040429381227601036, -0.0044454989520343159, 
    -0.0048129571433241968, -0.005140845859179349, -0.0054252098826181126, 
    -0.0056626635182842697, -0.0058504350684361345, -0.0059863659693727561, 
    -0.0060689449151841626, -0.0060972972468534585, -0.0060711811218495193, 
    -0.005990999584803724, -0.0058578040630835205, -0.0056732979346485373, 
    -0.0054398500502719164, -0.0051604719131409524, -0.004838820994916916, 
    -0.0044791779264454802, -0.0040863846286154238, -0.0036657889967399884, 
    -0.0032231632812185331, -0.0027646057221248307, -0.002296424860278467, 
    -0.0018250221749364418, -0.0013567669442682215, -0.00089787412468171678, 
    -0.00045427699935813388, -3.1545391541791973e-05, 0.00036518734802062854, 
    0.00073129238949817626, 0.0010626526481900093, 0.0013556854964601646, 
    0.00160734194214705, 0.0018151024699104546, 0.0019770002893122222, 
    0.0020916376751981876, 0.0021581819686195217, 0.0021763618203979721, 
    0.0021464670270565189, 0.002069310697256117, 0.001946194092873805, 
    0.0017788717687932951, 0.001569503705562701, 0.0013205867515930253, 
    0.0010348658885165416, 0.00071525361263299436, 0.00036471622897217906, 
    -1.3841736388700131e-05, -0.00041762714831330343, 
    -0.00084396930228819336, -0.0012902537781553087, -0.0017538152635963654, 
    -0.0022317912391444819, -0.0027209731697910339, -0.0032177029512731751, 
    -0.0037178268092760581, -0.0042168035704528324, -0.0047098423954292081, 
    -0.0051922104089442587, -0.0056594652717363737, -0.0061076751554755187, 
    -0.0065334798030052127, -0.0069341111915304805, -0.0073073569284574013, 
    -0.0076515170189222666, -0.0079653824630639726, -0.0082482577840960053, 
    -0.0084999254064510813, -0.0087206587153479745, -0.0089111581310963289, 
    -0.0090725253611506854, -0.0092061527952124571, -0.0093136478189594259, 
    -0.0093967334027152717, -0.0094571582518152321, -0.0094966192667380253, 
    -0.0095167231622613844, -0.0095189181828427179, -0.0095045139544292813, 
    -0.0094746926346088133, -0.0094305227824905604, -0.0093729886450976824, 
    -0.0093030533447918274, -0.0092216862538903356, -0.0091298924368196904, 
    -0.0090287735097051708, -0.0089195072835187572, -0.0088033970872222322, 
    -0.0086818397290719385, -0.0085563592282795371, -0.008428567246149354, 
    -0.0083001677221183727, -0.0081729756365718532, -0.0080489016690353243, 
    -0.0079298896136707382, -0.0078178613457691344, -0.0077146137026359958, 
    -0.0076217473511977192, -0.007540632416136523, -0.0074724155100953614, 
    -0.0074180800397592988, -0.0073785306120061206, -0.0073547437238760706, 
    -0.0073478783800935933, -0.0073593893464907641, -0.0073911003113901041, 
    -0.0074451902261417832, -0.0075241591455804998, -0.0076306795128837784, 
    -0.007767424549470785, -0.0079368043349133596, -0.0081407089435854944, 
    -0.0083802330686463221, -0.0086554833976594005, -0.0089654626741460033, 
    -0.009307991193642777, -0.009679793725006252, -0.01007656635021071, 
    -0.010493139734600171, -0.010923655737758942, -0.011361759589963126, 
    -0.01180082051682165, -0.012234134316861793, -0.012655114838566218, 
    -0.013057429131432092, -0.013435166453173756, -0.013782872117858072, 
    -0.014095623415637529, -0.014368998577652689, -0.014599103495204924, 
    -0.014782553674213215, -0.014916537628684773, -0.014998888482077153, 
    -0.015028214978450418, -0.015003975676566493, -0.014926497222526666, 
    -0.014796960962894908, -0.014617282018961224, -0.01438995088793776, 
    -0.014117874906735554, -0.013804263639943047, -0.013452438883772859, 
    -0.013065763361450681, -0.012647562939414511, -0.012201109498356785, 
    -0.011729582801452046, -0.011236114417110494, -0.010723825287952434, 
    -0.010195909110341437, -0.0096557039399366301, -0.0091067473309539952, 
    -0.0085527761170924831, -0.007997691304839941, -0.0074454205852792724, 
    -0.0068997543504990544, -0.0063641167237598554, -0.005841307536449048, 
    -0.0053332751235671593, -0.004840939490175747, -0.0043640713262001578, 
    -0.0039012758533517114, -0.0034501330098061075, -0.0030073349523828136, 
    -0.0025689076538621368, -0.0021304402193854399, -0.0016873649325708888, 
    -0.001235126839236727, -0.00076940585546760227, -0.00028627352020822575, 
    0.00021761247279687462, 0.00074495332551641332, 0.0012976243985958749, 
    0.0018765350045180272, 0.0024815624156329409, 0.0031113387696279997, 
    0.0037631543177398742, 0.0044328686663224221, 0.0051148275490645973, 
    0.0058018483154293459, 0.006485339081424589, 0.007155437058142187, 
    0.0078012864897989628, 0.0084115824526847325, 0.0089750153253803505, 
    0.0094809660414211308, 0.0099201532774795959, 0.010285237856439733, 
    0.010571302669266747, 0.010776146265640324, 0.010900464432913476, 
    0.010947549506931557, 0.010923189172708141, 0.010835113898938133, 
    0.010692454461634249, 0.01050515669008084, 0.010283181553228752, 
    0.010035741140581636, 0.0097705654538279389, 0.0094930186350359585, 
    0.0092055670583634022, 0.0089072402448859087, 0.0085935848189790092, 
    0.008256913816450483, 0.0078870223530399502, 0.0074718477863463112, 
    0.0069987713356764077, 0.006455797674613014, 0.0058327635718305624, 
    0.0051223213404212702, 0.0043206936495277029, 0.0034282128183059134, 
    0.0024492628871608936, 0.0013920328928988138, 0.00026765911162395569, 
    -0.0009103838331062337, -0.002127467459251145, -0.00336828856075903, 
    -0.0046180997178718285, -0.0058627895130982316, -0.0070900060352850208, 
    -0.0082885327562004472, -0.0094485963274417457, -0.010561381323024768,
  // Fqt-Na(4, 0-1999)
    1, 0.99757817015951877, 0.99036246758306068, 0.97849974693500841, 
    0.96222739002813229, 0.94186316263759917, 0.91779212783666553, 
    0.89045156574495665, 0.86031487635886272, 0.827875426831163, 
    0.79363119198592924, 0.75807085439117938, 0.72166185807225736, 
    0.68484071454866247, 0.64800565761879347, 0.61151161813727628, 
    0.57566734950226783, 0.54073447677491793, 0.50692814422214272, 
    0.47441898463717658, 0.44333606853561508, 0.41377055650048378, 
    0.38577977892102661, 0.35939150472501691, 0.33460823181167187, 
    0.31141132779649838, 0.28976493276906479, 0.26961954901742619, 
    0.25091526168499256, 0.23358458102162183, 0.21755490093464927, 
    0.20275057713657677, 0.1890946643394523, 0.17651032391989055, 
    0.164921941199069, 0.15425597741610034, 0.14444160456781727, 
    0.1354111527724923, 0.12710040727139629, 0.11944880632447163, 
    0.11239954412631969, 0.10589963467014887, 0.099899911490162724, 
    0.094355012360265833, 0.089223312367853164, 0.084466833254621787, 
    0.080051117196762112, 0.075945071125651922, 0.072120784120522377, 
    0.068553323202539762, 0.065220505662050982, 0.06210266865710172, 
    0.059182424023482033, 0.056444420144190002, 0.053875104730615769, 
    0.051462499993002869, 0.049195986942408801, 0.047066105705921762, 
    0.045064373736702967, 0.043183132036646157, 0.041415396703571035, 
    0.039754742185840387, 0.03819520049280728, 0.036731165006920627, 
    0.03535731217976739, 0.034068528697348624, 0.03285984401433132, 
    0.031726387099876574, 0.030663345181396916, 0.02966594331400178, 
    0.028729440969215283, 0.027849125957753369, 0.027020319979436935, 
    0.026238373260393962, 0.02549866736845724, 0.024796614673009958, 
    0.024127655326133046, 0.0234872674444194, 0.022870982943807981, 
    0.022274414554902006, 0.02169328972960867, 0.021123503125276614, 
    0.020561166566069537, 0.020002673181551276, 0.019444757636662161, 
    0.018884551805906192, 0.018319639529612925, 0.017748093763903593, 
    0.017168502268043912, 0.01657996819774905, 0.015982108943503385, 
    0.015375026167382804, 0.014759279506071563, 0.014135849725133431, 
    0.013506095448646603, 0.012871712241253072, 0.012234686702522214, 
    0.011597244654348389, 0.010961790343098339, 0.010330851079357556, 
    0.0097070084634121312, 0.0090928285230341827, 0.0084907954169252727, 
    0.0079032479358655226, 0.0073323281455339347, 0.0067799403183886374, 
    0.0062477277841468436, 0.0057370677135861366, 0.0052490797721933139, 
    0.0047846555811692643, 0.004344499900120642, 0.0039291796845050322, 
    0.0035391867008623948, 0.0031749822434852808, 0.0028370492701081463, 
    0.0025259207855389989, 0.002242195161707755, 0.0019865293973886288, 
    0.0017596247577890377, 0.0015622033454958965, 0.0013949759522332598, 
    0.0012586160270276459, 0.0011537302601378854, 0.0010808409897627167, 
    0.0010403599814791853, 0.0010325756930438241, 0.0010576346911232134, 
    0.0011155241478009838, 0.0012060514952140185, 0.001328820080342828, 
    0.0014831998774702563, 0.0016682996930002347, 0.0018829321079419166, 
    0.0021255829342280972, 0.0023943930455508997, 0.0026871458101904622, 
    0.0030012814075409218, 0.0033339187404576422, 0.0036818998460008442, 
    0.0040418451278892674, 0.0044102175376903021, 0.0047833920143772312, 
    0.0051577207887013631, 0.0055295996037021825, 0.0058955204181168168, 
    0.0062521135395659996, 0.0065961842070770367, 0.0069247312834474026, 
    0.0072349627322070703, 0.0075243034249982471, 0.0077904032139443071, 
    0.0080311307072308234, 0.0082445924052838206, 0.0084291341692298138, 
    0.0085833578456547422, 0.0087061405856500781, 0.0087966462278308965, 
    0.008854353852062043, 0.0088790689570837043, 0.0088709503388397972, 
    0.0088305273972004005, 0.0087587236655713406, 0.008656868769413309, 
    0.0085267047221421425, 0.008370377921040395, 0.0081904121144206112, 
    0.0079896653843882764, 0.0077712621171094108, 0.0075385227828920522, 
    0.0072948754924687092, 0.0070437821026655117, 0.0067886681403848117, 
    0.0065328637617120804, 0.0062795460410321711, 0.0060316945096741195, 
    0.0057920442294690736, 0.0055630519244314136, 0.00534686060421338, 
    0.0051452748208788953, 0.0049597411030386429, 0.0047913298553465319, 
    0.004640732968820057, 0.004508257204775999, 0.0043938363583628948, 
    0.0042970434406994001, 0.0042171249596168548, 0.0041530312091082964, 
    0.0041034643103093158, 0.0040669272107949159, 0.0040417810563064755, 
    0.00402629891925654, 0.0040187237969827108, 0.0040173221811666349, 
    0.0040204318887683659, 0.0040265050943648541, 0.0040341403734263119, 
    0.0040421105493571741, 0.0040493843705599096, 0.0040551307542835424, 
    0.0040587172111797758, 0.0040596956242164505, 0.0040577814209933529, 
    0.004052819423424588, 0.0040447540676598996, 0.0040335945638363332, 
    0.0040193829573478028, 0.0040021674435350629, 0.0039819832102527359, 
    0.0039588404414274718, 0.0039327261383144052, 0.0039036067503087665, 
    0.0038714506466078751, 0.0038362515280621389, 0.0037980590024910381, 
    0.0037570082872527195, 0.0037133519301595333, 0.0036674756597883979, 
    0.0036199147405163975, 0.0035713376348696681, 0.0035225329992403585, 
    0.0034743634251009959, 0.0034277161563009114, 0.0033834412173758227, 
    0.0033422883418876069, 0.0033048437893500576, 0.0032714729305653124, 
    0.0032422751530728688, 0.0032170507769633937, 0.003195287933971815, 
    0.0031761619107816361, 0.0031585646550657547, 0.0031411413609163312, 
    0.0031223484827038743, 0.0031005256816220906, 0.0030739711070339, 
    0.0030410235673550296, 0.0030001379081251722, 0.0029499553972965795, 
    0.0028893594380792562, 0.0028175137025204721, 0.0027338847753618943, 
    0.0026382425138224948, 0.0025306394599205204, 0.0024113812687883499, 
    0.002280976844530983, 0.0021400880764500365, 0.0019894667645708637, 
    0.0018299010795901473, 0.0016621617785697971, 0.0014869624783549057, 
    0.0013049236183534021, 0.0011165603751474365, 0.00092227959389177563, 
    0.00072238998158083336, 0.00051712810383251426, 0.00030669637205273646, 
    9.1315956764403939e-05, -0.00012871201477764722, -0.00035294084588964603, 
    -0.00058071867034640223, -0.00081113762424609684, -0.0010430009789442235, 
    -0.0012748169155422267, -0.0015048183546358075, -0.0017309974544770497, 
    -0.0019511564720264872, -0.0021629620135725793, -0.0023640035026802619, 
    -0.0025518473931941681, -0.002724079326945641, -0.0028783520904923769, 
    -0.0030124218279617837, -0.0031241816310391161, -0.0032116971447468138, 
    -0.0032732264268720535, -0.0033072442431826242, -0.0033124539570573565, 
    -0.0032877956466229497, -0.0032324535823358607, -0.0031458488559523066, 
    -0.0030276453429656466, -0.0028777467839089786, -0.0026963049993390395, 
    -0.0024837225996735017, -0.0022406653767479173, -0.0019680747252821076, 
    -0.0016671810607801556, -0.0013395129973214823, -0.00098691009299511738, 
    -0.00061152833724789342, -0.00021584959471730671, 0.0001973185875349682, 
    0.00062484087467675777, 0.0010632620790104374, 0.0015088203558233631, 
    0.0019574719008895458, 0.0024049222706531976, 0.002846675282692611, 
    0.0032780913506756082, 0.0036944600127095709, 0.0040910835596769815, 
    0.0044633666745665128, 0.0048069150001837585, 0.0051176319552408336, 
    0.0053918155210012251, 0.0056262439344779754, 0.0058182497582140716, 
    0.0059657741797109259, 0.0060674032972364723, 0.0061223770873744783, 
    0.0061305843576642295, 0.0060925390540408414, 0.0060093445961991393, 
    0.0058826493732293018, 0.0057145877466889287, 0.0055077252410895942, 
    0.005264993683592299, 0.0049896281928534783, 0.0046851052477353003, 
    0.0043550804925110561, 0.0040033191194566503, 0.0036336243863130313, 
    0.0032497594633261696, 0.0028553609945073423, 0.002453850443361875, 
    0.0020483488963011823, 0.0016415920889727834, 0.0012358756331284995, 
    0.00083300809647241598, 0.00043431217088649214, 4.0654314397361221e-05, 
    -0.00034747661166598532, -0.00072986127887225065, -0.0011064118807961577, 
    -0.0014770236673422015, -0.0018414352883160501, -0.0021991203125632203, 
    -0.0025492117425364252, -0.0028904617467176595, -0.0032212491569112772, 
    -0.003539613040793913, -0.0038433147343017171, -0.0041299147789060978, 
    -0.0043968634937684289, -0.0046416014396950317, -0.0048616556713012753, 
    -0.0050547374602848668, -0.0052188307152734566, -0.0053522682328119575, 
    -0.0054537869021274088, -0.0055225748720175013, -0.0055582908492153617, 
    -0.0055610681507539473, -0.0055315027488555338, -0.0054706269144339263, 
    -0.0053798719301503001, -0.0052610190736670408, -0.0051161368770126564, 
    -0.0049475140276943781, -0.0047575830532896775, -0.0045488399073132738, 
    -0.0043237676372997989, -0.0040847639563359817, -0.0038340784020837299, 
    -0.0035737596484096252, -0.003305614244736139, -0.0030311821151462878, 
    -0.0027517219377788185, -0.0024682089161191705, -0.0021813528920793346, 
    -0.0018916224175984471, -0.0015992840725081235, -0.0013044479610492669, 
    -0.0010071197353699768, -0.00070724727610137618, -0.0004047679281717563, 
    -9.9642243286095689e-05, 0.00020811691076599284, 0.00051842436297660718, 
    0.00083111020336825337, 0.0011459096574904443, 0.0014624590096225399, 
    0.0017802882915002327, 0.0020988176953786351, 0.0024173520316596486, 
    0.0027350765704816926, 0.0030510554928750914, 0.0033642344090016301, 
    0.0036734526981780811, 0.0039774541195604857, 0.0042749060173362871, 
    0.0045644182797804052, 0.004844563898608354, 0.0051139158924352768, 
    0.0053710767632853349, 0.0056147267244847972, 0.0058436626451267267, 
    0.006056835064989192, 0.0062533802260427897, 0.0064326459747983504, 
    0.0065942089205723855, 0.0067378864389202762, 0.0068637254347842522, 
    0.0069719928093495082, 0.007063142691090752, 0.0071377732455716091, 
    0.007196578683744773, 0.0072402978953573279, 0.007269661630172071, 
    0.007285348021254804, 0.007287945075302572, 0.0072779222166367476, 
    0.0072556154682706479, 0.0072212268565365733, 0.0071748233273942405, 
    0.0071163534125498621, 0.0070456599372305442, 0.006962499978711169, 
    0.0068665663989798511, 0.0067575156197104812, 0.0066350014105676638, 
    0.0064987174636997064, 0.0063484390805583213, 0.0061840689063852837, 
    0.0060056770278612698, 0.0058135400282822861, 0.005608169077641981, 
    0.0053903366550897532, 0.0051610880279942001, 0.004921743227488261, 
    0.0046738890968745913, 0.004419349572108505, 0.0041601437410439734, 
    0.0038984256393342662, 0.0036364108604695056, 0.0033763070056925994, 
    0.0031202409271291328, 0.0028702000784430258, 0.0026279822636463192, 
    0.0023951671132532741, 0.0021730948356745634, 0.001962868731339368, 
    0.0017653638780286234, 0.0015812487436400672, 0.0014110098460546464, 
    0.0012549780522370683, 0.0011133540605552847, 0.00098622513331278494, 
    0.00087358233781585734, 0.00077532276200234366, 0.00069124832153573564, 
    0.00062104954082680807, 0.00056428540410900611, 0.00052035052717328543, 
    0.00048844458453009641, 0.00046754294709590544, 0.00045638373166204073, 
    0.00045347381824707158, 0.00045711030751553744, 0.00046543091997854172, 
    0.00047647324402520417, 0.00048824335380161623, 0.00049879102583013908, 
    0.00050627708948389042, 0.00050904209942924503, 0.00050566229150184722, 
    0.00049499930505446247, 0.00047623244502582992, 0.0004488863618996234, 
    0.00041283660196656826, 0.00036830224383332114, 0.00031582376686336005, 
    0.00025622730212283872, 0.00019058051550203522, 0.000120138860952129, 
    4.6290995014149734e-05, -2.9494556839522327e-05, -0.00010572865256123267, 
    -0.00018095118478573941, -0.00025378579126152052, 
    -0.00032298525592384822, -0.00038747426707594129, 
    -0.00044638384193502903, -0.00049908349303434034, 
    -0.00054519796210450596, -0.00058462931728399826, 
    -0.00061755519502861684, -0.00064443250051724832, 
    -0.00066598470351214903, -0.0006831698437424912, -0.00069715282240437261, 
    -0.00070924556987458681, -0.00072085197718999505, 
    -0.00073339927886651086, -0.00074827785270379786, 
    -0.00076678206937648733, -0.00079007028557938385, 
    -0.00081913150543303317, -0.00085476560594933255, 
    -0.00089757277908660601, -0.00094795355823870827, -0.001006107471893194, 
    -0.0010720438114339168, -0.0011455880652203269, -0.0012263944670742224, 
    -0.0013139596712925384, -0.0014076483119681476, -0.0015067205675816076, 
    -0.0016103598692779023, -0.0017177050347417671, -0.0018278661620398846, 
    -0.0019399318269469621, -0.0020529666589567479, -0.0021660027181421766, 
    -0.0022780275757727851, -0.0023879787742832788, -0.0024947428861225559, 
    -0.002597158622663992, -0.0026940331714360708, -0.002784156644239599, 
    -0.0028663174632637114, -0.002939320630339054, -0.0030020009146520597, 
    -0.0030532356275591349, -0.0030919582251610605, -0.0031171628237199882, 
    -0.0031279192424182025, -0.0031233945139758747, -0.0031028901103294362, 
    -0.0030658844968918407, -0.0030120897802026311, -0.0029414993044412693, 
    -0.0028544212582285516, -0.002751502866021628, -0.0026337345351193676, 
    -0.0025024359993315458, -0.0023592246859415471, -0.002205965265819163, 
    -0.0020447014040341667, -0.0018775748304483033, -0.0017067307631400178, 
    -0.0015342220135959703, -0.0013619158419407454, -0.0011914049162683289, 
    -0.0010239276313767668, -0.00086030742129947994, -0.00070090368277411579, 
    -0.00054559053877212987, -0.00039375129344734478, 
    -0.00024430550818030068, -9.5747573765029279e-05, 5.378757809894368e-05, 
    0.00020644377768370417, 0.00036455600308132842, 0.00053054737705700945, 
    0.00070682278351090499, 0.00089566212080747771, 0.0010991112702140905, 
    0.001318883009991695, 0.0015562649407411221, 0.0018120449235421924, 
    0.0020864529451019498, 0.0023791216481093723, 0.0026890682504932947, 
    0.0030146974117906873, 0.0033538232194483038, 0.0037037080191326026, 
    0.0040611297014181416, 0.0044224642419887729, 0.0047837786183766145, 
    0.0051409472008263546, 0.0054897663843272385, 0.0058260753281548254, 
    0.006145871675541272, 0.0064454119047855137, 0.0067213043227083167, 
    0.0069705825579870935, 0.0071907583488613064, 0.0073798605765183619, 
    0.0075364490062501364, 0.0076596199663747019, 0.0077489843723917585, 
    0.00780463584769037, 0.0078271063524515856, 0.0078173171489384439, 
    0.0077765138528665349, 0.0077062127640779802, 0.0076081310381473626, 
    0.0074841335693093597, 0.0073361731211395043, 0.0071662437789572165, 
    0.0069763442786016979, 0.0067684493161350645, 0.0065444987021052873, 
    0.0063063960765979039, 0.006056023797855188, 0.0057952603745525738, 
    0.005526004702816445, 0.0052501987399608107, 0.0049698446890663389, 
    0.0046870145762062457, 0.0044038499432759119, 0.0041225559484148857, 
    0.0038453829320679481, 0.0035746062934561957, 0.003312494216515928, 
    0.0030612775055541539, 0.0028231125108700936, 0.0026000445127685999, 
    0.002393971510901669, 0.0022066091083918745, 0.0020394588610885057, 
    0.0018937807386853163, 0.0017705726659726835, 0.0016705516656519246, 
    0.0015941472428398188, 0.0015414918510189028, 0.00151241853542, 
    0.0015064620460432505, 0.0015228602065398109, 0.0015605609547702597, 
    0.0016182246159609319, 0.0016942334576929006, 0.0017867034699749101, 
    0.0018934958369302409, 0.0020122367511312324, 0.0021403460034244027, 
    0.0022750671040890503, 0.0024135059094000794, 0.0025526695979492687, 
    0.0026895107792331697, 0.0028209675457578297, 0.0029440167378647028, 
    0.003055714669155656, 0.0031532554591398917, 0.0032340173979374283, 
    0.0032956232100261199, 0.0033359976144348544, 0.0033534235039383124, 
    0.0033465947738491788, 0.0033146582837498234, 0.0032572455164150207, 
    0.0031744849522073429, 0.0030670001101575587, 0.0029358835285384919, 
    0.0027826595540763896, 0.0026092413334543379, 0.0024178720731324915, 
    0.0022110764196130463, 0.0019916012397983704, 0.0017623650601189893, 
    0.001526398869136426, 0.0012867915574103733, 0.0010466291585705689, 
    0.00080893624063053439, 0.00057661338556460489, 0.00035237435380739378, 
    0.00013868888548818981, -6.2272172950108054e-05, -0.00024868879732258627, 
    -0.00041912638192109612, -0.00057256183780415545, 
    -0.00070838902969149917, -0.00082640463507710742, 
    -0.00092677775773964983, -0.0010099952360170896, -0.0010768026694158435, 
    -0.0011281294731320638, -0.0011650171198990581, -0.0011885539617404318, 
    -0.0011998271755711313, -0.0011998898058080401, -0.0011897564127761426, 
    -0.0011704121041606434, -0.001142847090420924, -0.0011080931036596625, 
    -0.0010672718083778725, -0.0010216371038949293, -0.0009726160745244897, 
    -0.00092183848203870964, -0.00087114298961522829, 
    -0.00082257306458846332, -0.00077834261359023755, -0.0007407753979911659, 
    -0.00071222864645685677, -0.00069500442502983505, 
    -0.00069125596459548334, -0.00070289359585002753, 
    -0.00073150979759458877, -0.00077831057107641906, 
    -0.00084406896115425103, -0.00092908596549191598, -0.0010331818163864363, 
    -0.0011556892725444199, -0.0012954720000827786, -0.001450946723445735, 
    -0.0016201348557016927, -0.0018007196786997803, -0.0019901302929337126, 
    -0.0021856281545896278, -0.0023843996147437344, -0.0025836367911835174, 
    -0.0027806076633197165, -0.002972716883638146, -0.0031575417890641901, 
    -0.0033328731795674834, -0.003496720695228201, -0.0036473331136849959, 
    -0.0037831933431810567, -0.0039030237775873949, -0.004005782625113875, 
    -0.0040906549651866658, -0.0041570546483000207, -0.0042046075438395255, 
    -0.0042331418137504413, -0.0042426712308954052, -0.0042333737385383497, 
    -0.0042055707198913076, -0.0041597009051187418, -0.0040963083832705567, 
    -0.0040160235100036691, -0.0039195607663482486, -0.0038077195837291386, 
    -0.0036813896774560173, -0.0035415613911272009, -0.0033893385602852188, 
    -0.0032259522367805524, -0.0030527617809017228, -0.0028712666662726624, 
    -0.0026831069037264697, -0.0024900571314626333, -0.0022940193561735004, 
    -0.002097003333395677, -0.0019011055801275575, -0.0017084693705699549, 
    -0.0015212444875917375, -0.0013415340339532117, -0.0011713384257366071, 
    -0.0010125011781873668, -0.00086666231021118099, -0.00073522239650611408, 
    -0.00061932354647734706, -0.00051984574717019031, 
    -0.00043742783131123654, -0.00037249738120645617, 
    -0.00032531380329719236, -0.00029601317520993367, 
    -0.00028464892669515445, -0.00029121861282151791, 
    -0.00031568071466605939, -0.00035796366846262796, 
    -0.00041796108960142432, -0.00049551612610183274, 
    -0.00059039517977812627, -0.00070225477503053706, 
    -0.00083061101379908674, -0.00097480678674854125, -0.0011339971196784296, 
    -0.0013071399526836433, -0.001492995394577425, -0.0016901369241902817, 
    -0.0018969683974538801, -0.0021117492660450714, -0.0023326276975789606, 
    -0.0025576720364493522, -0.0027849092051603734, -0.0030123521122658388, 
    -0.0032380295934108108, -0.0034600040489957819, -0.0036763793806626269, 
    -0.0038853045871804297, -0.0040849574307792215, -0.004273537675534512, 
    -0.0044492464015861771, -0.0046102796215390833, -0.0047548237617998082, 
    -0.0048810602382437247, -0.0049871767385039258, -0.0050713854282665571, 
    -0.0051319477215473058, -0.0051672002809032141, -0.0051755893534872434, 
    -0.0051557068478095946, -0.0051063334286318282, -0.0050264823738831819, 
    -0.0049154519237836715, -0.0047728699393892347, -0.00459874060615379, 
    -0.004393478002154028, -0.0041579333357330507, -0.0038934038576930443, 
    -0.0036016248499774394, -0.0032847590583129525, -0.0029453632601750528, 
    -0.0025863593184112582, -0.002210994193521981, -0.0018228062952309848, 
    -0.0014255833035157527, -0.0010233174808870643, -0.00062015951222167459, 
    -0.00022035920450924607, 0.00017179794119233702, 0.0005520529092304027, 
    0.00091625409246206874, 0.0012604333218546025, 0.0015808853819732952, 
    0.0018742537152324709, 0.0021376080538845123, 0.0023685099519913672, 
    0.0025650671391542219, 0.0027259674416437321, 0.0028504841455561335, 
    0.0029384581993522393, 0.0029902639385448182, 0.0030067600635713078, 
    0.0029892354635634734, 0.0029393474075259944, 0.0028590642696822081, 
    0.0027506074464290582, 0.0026163886836575285, 0.0024589556440934861, 
    0.002280933576131973, 0.0020849682070173499, 0.0018736720530015166, 
    0.0016495783208109553, 0.0014150935373032911, 0.0011724653982037611, 
    0.00092375337280984206, 0.00067081341051579099, 0.00041529126635340822, 
    0.00015861834095959857, -9.7979639095888764e-05, -0.00035347569823931436, 
    -0.00060701857191887095, -0.00085791899941042133, -0.0011056217247708325, 
    -0.0013496820462843065, -0.0015897418851272831, -0.0018255069375391092, 
    -0.0020567308045743075, -0.0022831979536766917, -0.0025047206539606276, 
    -0.0027211352664381584, -0.0029323057900571795, -0.0031381343175858473, 
    -0.0033385641578888114, -0.0035335889235149089, -0.0037232548516933834, 
    -0.0039076579503511044, -0.004086930063375932, -0.004261225251040399, 
    -0.0044306932829602016, -0.0045954543346591889, -0.0047555640071132322, 
    -0.0049109824212326906, -0.0050615416092988667, -0.0052069168281958138, 
    -0.0053466022741789458, -0.0054799058402053985, -0.0056059469870548785, 
    -0.0057236801501805209, -0.0058319237765734611, -0.0059294009770083558, 
    -0.006014785421806901, -0.0060867482182950508, -0.0061440035045318437, 
    -0.0061853562195126758, -0.0062097446815541062, -0.0062162854844183199, 
    -0.0062043182131307096, -0.006173444062118158, -0.0061235667409552186, 
    -0.0060549224435140526, -0.0059681026179187295, -0.005864062097549516, 
    -0.0057441074070022384, -0.0056098694219172086, -0.0054632658409137745, 
    -0.0053064446832477401, -0.0051417304410418261, -0.0049715619309769823, 
    -0.0047984318610100711, -0.004624831485887112, -0.0044531904956821959, 
    -0.0042858251343265152, -0.0041248778855702533, -0.0039722642473001852, 
    -0.003829629929667404, -0.003698312183977666, -0.003579321827866903, 
    -0.0034733393808448585, -0.0033807252842776398, -0.0033015457840177937, 
    -0.0032356039573550512, -0.0031824767895697595, -0.003141549698021441, 
    -0.0031120411976019234, -0.003093029142824796, -0.0030834595717394437, 
    -0.0030821541699177246, -0.0030878118627674562, -0.0030990126828642551, 
    -0.0031142309282061386, -0.0031318629803442737, -0.0031502694166592403, 
    -0.0031678298135288342, -0.003183005732317569, -0.0031943972193642063, 
    -0.0032007923278016162, -0.0032011942985097513, -0.0031948336848611784, 
    -0.0031811657929441241, -0.0031598702328534548, -0.0031308461106607289, 
    -0.0030942081882361725, -0.0030502868236971336, -0.0029996071241641695, 
    -0.0029428654480319902, -0.0028808877863885827, -0.002814586202622143, 
    -0.0027449088851717405, -0.0026727931779486234, -0.002599128123300311, 
    -0.0025247279455545019, -0.002450316402751646, -0.0023765239981260351, 
    -0.0023038938834908174, -0.0022328943580510905, -0.0021639276361623554, 
    -0.0020973417170314442, -0.0020334388544857103, -0.0019724732029248737, 
    -0.0019146515534284509, -0.0018601326877383134, -0.0018090247770308921, 
    -0.0017613863349699975, -0.0017172342104369044, -0.0016765605960337114, 
    -0.0016393555635045472, -0.0016056364571228206, -0.0015754757427807518, 
    -0.0015490220651474085, -0.0015265125500393091, -0.0015082729069725077, 
    -0.0014947049985025124, -0.0014862631469178336, -0.0014834253603418918, 
    -0.0014866592337605586, -0.0014963912849286251, -0.0015129805815100954, 
    -0.0015366905129089331, -0.001567673907155195, -0.001605950041562195, 
    -0.0016513941911728341, -0.001703728383657874, -0.0017625175510395453, 
    -0.0018271710541315257, -0.0018969523988845351, -0.0019709925741452773, 
    -0.0020483093143192832, -0.0021278319506202702, -0.0022084252917932909, 
    -0.002288914377159701, -0.0023681050818171183, -0.0024447971879527717, 
    -0.0025177937465950206, -0.0025859076926656737, -0.0026479652644374996, 
    -0.0027028127423474064, -0.0027493262103626521, -0.0027864301916490346, 
    -0.002813121261128045, -0.0028284980587924943, -0.0028317930764952788, 
    -0.0028223964055463036, -0.0027998860535867992, -0.0027640425421375982, 
    -0.0027148533184230528, -0.0026525223171488315, -0.0025774583081933072, 
    -0.002490279410730328, -0.0023918070104904801, -0.0022830656119177703, 
    -0.0021652835622490161, -0.0020398932610993072, -0.0019085292093045545, 
    -0.0017730211858442084, -0.0016353807426063955, -0.0014977788791842171, 
    -0.0013625141479755257, -0.0012319590435618845, -0.0011085055233174591, 
    -0.00099448620509153224, -0.00089208624873464502, 
    -0.00080326555633774286, -0.00072967976217695046, 
    -0.00067262410752229405, -0.00063299138073353992, -0.0006112523672084163, 
    -0.00060745030468920967, -0.00062121014799779509, 
    -0.00065176288018259257, -0.00069798125259576925, 
    -0.00075842353738359545, -0.00083139412144239938, 
    -0.00091500096468548353, -0.0010072155515744954, -0.0011059217861376933, 
    -0.0012089528144322722, -0.0013141210523088592, -0.0014192314006015328, 
    -0.0015221013769633517, -0.0016205800293681025, -0.0017125901970490402, 
    -0.0017961726905668526, -0.0018695426295638063, -0.0019311409654336705, 
    -0.0019796745053818326, -0.0020141514267025158, -0.0020339053610778481, 
    -0.002038608968212677, -0.0020282963862507889, -0.0020033701943896857, 
    -0.001964612336615709, -0.0019131821222221547, -0.0018506047850268912, 
    -0.001778742875113472, -0.001699749536641561, -0.0016160071703317882, 
    -0.001530056249155882, -0.0014445154873961527, -0.0013619982769956704, 
    -0.0012850400401534915, -0.0012160220160507182, -0.0011571124389326312, 
    -0.0011102165804278245, -0.0010769383202882035, -0.0010585541254030124, 
    -0.0010560027451815132, -0.0010698804357703361, -0.0011004590125915834, 
    -0.0011476975492585766, -0.0012112711581868092, -0.0012905879190153082, 
    -0.0013848105019976216, -0.0014928602473476124, -0.0016134190629329525, 
    -0.0017449226505849391, -0.0018855505009886336, -0.0020332262786284323, 
    -0.0021856261284325367, -0.0023402048653574006, -0.0024942461555581266, 
    -0.0026449245609436304, -0.0027893771240666402, -0.0029247868391544182, 
    -0.0030484638088367796, -0.0031579172793031402, -0.0032509271604060654, 
    -0.0033255990697724364, -0.0033804117191316447, -0.0034142510818157131, 
    -0.0034264359950955995, -0.0034167220390189782, -0.0033852938330592524, 
    -0.0033327222398321812, -0.0032599162299100986, -0.0031680492634493193, 
    -0.0030584745270465031, -0.0029326396323031516, -0.0027919958357467971, 
    -0.0026379210571188918, -0.0024716438458679442, -0.0022941893057968326, 
    -0.002106340095760112, -0.0019086230233411965, -0.0017013262028129767, 
    -0.0014845334741300158, -0.001258193625584823, -0.0010221966480109649, 
    -0.00077646104777479876, -0.00052101600991429271, 
    -0.00025607012693719709, 1.7937866828673173e-05, 0.00030030905321596512, 
    0.0005900734100141371, 0.00088599105311593042, 0.0011865623915434315, 
    0.0014900519326853637, 0.0017945107108176537, 0.0020978091086999483, 
    0.0023976664989715834, 0.0026916780622239741, 0.0029773425728900457, 
    0.0032520875168262028, 0.0035133008891109199, 0.0037583583833711563, 
    0.0039846665403658332, 0.0041897063676388929, 0.0043710794341189621, 
    0.0045265579987255385, 0.0046541398180263635, 0.0047521015120901774, 
    0.0048190532141507104, 0.0048539910294545605, 0.0048563453146365822, 
    0.0048260158799043771, 0.0047633945648428936, 0.004669373655700311, 
    0.0045453381576418391, 0.004393136875443667, 0.0042150433546839965, 
    0.0040136951390331932, 0.0037920300924455252, 0.0035532041051388533, 
    0.0033005066641471205, 0.0030372729320199934, 0.0027668062944261875, 
    0.0024923172433694817, 0.0022168764898989053, 0.0019433980030726362, 
    0.0016746416146318484, 0.0014132300953876322, 0.0011616712770456811, 
    0.00092237836208474864, 0.00069767831930999552, 0.00048980884916849821, 
    0.00030089817027810549, 0.00013294021855274622, -1.2234285498124455e-05, 
    -0.00013298729243458939, -0.0002278998467750838, -0.00029579909117276478, 
    -0.00033577276583460122, -0.000347191876188196, -0.00032972261544224449, 
    -0.00028333694095815815, -0.0002083188311891167, -0.00010527071873416249, 
    2.487965755172168e-05, 0.00018088233014000663, 0.0003611625607020989, 
    0.00056382763319704344, 0.000786668047138314, 0.0010271675849977161, 
    0.0012825163701724162, 0.0015496126434369319, 0.0018250891185606838, 
    0.0021053355190700416, 0.002386528290026549, 0.0026646848934298722, 
    0.002935718075331131, 0.0031955053768588952, 0.0034399742421175623, 
    0.0036651934321406472, 0.0038674667730661072, 0.0040434269340689786, 
    0.0041901240882265328, 0.004305095993258237, 0.0043864279520423061, 
    0.0044327913547113828, 0.0044434680064994745, 0.0044183557178134525, 
    0.0043579630226005719, 0.0042633909105511498, 0.0041362987966494218, 
    0.0039788611553523649, 0.0037937041664784792, 0.0035838384345694089, 
    0.0033525811643291287, 0.0031034689278292373, 0.0028401680913356332, 
    0.0025663882919972226, 0.0022857941820355757, 0.0020019345345852766, 
    0.0017181678106548495, 0.0014376114464027664, 0.001163100577216421, 
    0.00089716259081612146, 0.00064201428922296838, 0.00039956182172173416, 
    0.00017141817356824805, -4.1070448820882299e-05, -0.00023680233125216701, 
    -0.00041488977586791938, -0.00057463378125227507, 
    -0.00071551013627014462, -0.00083715206463975565, 
    -0.00093934875119606846, -0.0010220441432100518, -0.0010853460369919412, 
    -0.0011295339472495807, -0.0011550647258997491, -0.0011625779139451484, 
    -0.0011528917275313738, -0.0011269953751862584, -0.0010860317303254961, 
    -0.0010312757190142404, -0.00096410744750591076, -0.00088597623806973831, 
    -0.00079836613672612002, -0.00070275105969891676, 
    -0.00060054975996859275, -0.00049307398824509178, 
    -0.00038148622670886902, -0.00026676173289220863, 
    -0.00014966329461699093, -3.0732629623920604e-05, 8.9705328576670249e-05, 
    0.00021151877998773125, 0.00033474622896425654, 0.00045955482490228627, 
    0.00058621911993059239, 0.00071507176228059548, 0.00084647557445474719, 
    0.0009807771507210968, 0.001118260221324047, 0.0012590968049005832, 
    0.0014032983389969847, 0.0015506757849583098, 0.001700810062766472, 
    0.0018530326256439064, 0.0020064297093886998, 0.0021598524940482709, 
    0.0023119464208213635, 0.0024611817054175926, 0.0026058928652794057, 
    0.0027443145226515495, 0.0028746164221782437, 0.00299492806135931, 
    0.0031033733223683503, 0.00319809689956134, 0.0032772953909685977, 
    0.0033392540702280402, 0.0033823903454489618, 0.0034052949400861479, 
    0.0034067874849389949, 0.0033859551770028446, 0.0033422003947867246, 
    0.0032752771944833592, 0.0031853185697371398, 0.0030728571501154093, 
    0.002938829676581294, 0.0027845751556668055, 0.0026118157480235155, 
    0.0024226368906053739, 0.0022194540235564893, 0.0020049663105386542, 
    0.0017821048389859255, 0.001553981246378838, 0.0013238204405434529, 
    0.0010948819308023432, 0.00087038734694551163, 0.00065342657235139211, 
    0.00044686171618226259, 0.00025322617136623734, 7.4623578533450672e-05, 
    -8.7338830417712279e-05, -0.00023160431857257197, 
    -0.00035766952953960446, -0.00046556743576585061, 
    -0.00055581899538050439, -0.00062938627724139998, 
    -0.00068762261372710357, -0.00073222506077431026, 
    -0.00076520083035001537, -0.00078882164349043595, -0.0008055631541644139, 
    -0.00081802684751920945, -0.00082883920122977725, 
    -0.00084054116959946998, -0.00085548462466989925, 
    -0.00087573461113700339, -0.00090300286843044038, 
    -0.00093860247551793956, -0.00098343017009676608, -0.0010379669821302586, 
    -0.0011023085973698539, -0.0011761895381801721, -0.0012590239888310806, 
    -0.0013499441695574844, -0.0014478364768316185, -0.0015513971132216377, 
    -0.0016591753726762064, -0.0017696330207625714, -0.0018812101028207685, 
    -0.0019923775410717274, -0.0021016989147251797, -0.0022078645014070777, 
    -0.0023097234097714486, -0.0024062911928150184, -0.0024967508626174244, 
    -0.0025804383659910448, -0.0026568297740493922, -0.0027255239452032916, 
    -0.0027862280762677386, -0.0028387512648845163, -0.0028830036600495362, 
    -0.0029190026784421943, -0.002946875776020888, -0.0029668755071532555, 
    -0.0029793976085826582, -0.0029849947422546006, -0.0029844005876632591, 
    -0.0029785472201585448, -0.0029685868393219822, -0.0029558950382109284, 
    -0.0029420693199140443, -0.0029289044604406864, -0.0029183520163346263, 
    -0.0029124714083580915, -0.0029133689186499907, -0.002923151817871626, 
    -0.002943866830561576, -0.0029774504055037421, -0.0030256755696242551, 
    -0.0030901162701081394, -0.0031720966692251207, -0.0032726625629756747, 
    -0.0033925350774646782, -0.0035320824964195975, -0.0036912851036439024, 
    -0.0038697103097770674, -0.0040665109350934581, -0.0042804428222546565, 
    -0.0045098986540698192, -0.0047529609581260547, -0.0050074615298379256, 
    -0.0052710399215693338, -0.0055411954448557569, -0.0058153234757619019, 
    -0.0060907419937158234, -0.0063647198788319911, -0.0066344964392622127, 
    -0.0068973188306741748, -0.007150479904373187, -0.0073913724227080502, 
    -0.0076175435980838256, -0.0078267660865442117, -0.0080170960532810562, 
    -0.0081869364015133509, -0.0083351014168310776, -0.0084608656554029243, 
    -0.0085640227934906839, -0.0086449133310253102, -0.0087044417752143704, 
    -0.0087440620804037118, -0.0087657274470625025, -0.0087718086080785119, 
    -0.0087649732565190201, -0.0087480521499093706, -0.0087238872207554916, 
    -0.008695194542912876, -0.0086644441990866086, -0.0086337506190993507, 
    -0.0086048204695397881, -0.0085789092964234388, -0.0085568226102323685, 
    -0.0085389336345474513, -0.0085252245274527513, -0.0085153459215068835, 
    -0.0085086820840833775, -0.0085044336754708533, -0.0085017038927462391, 
    -0.0084995870404794057, -0.0084972539764705257, -0.0084940294414454481, 
    -0.0084894575085250334, -0.0084833401936962177, -0.0084757590407426118, 
    -0.0084670699928750988, -0.0084578614185042804, -0.0084489002156373106, 
    -0.008441058996016753, -0.0084352421150407503, -0.0084323275758610376, 
    -0.0084331156162191223, -0.0084382715349088575, -0.0084482670985420432, 
    -0.0084632923401293126, -0.0084831606041321402, -0.0085072217408665059, 
    -0.0085343082907100628, -0.0085627259290793449, -0.008590299226075012, 
    -0.0086144747811676484, -0.0086324553204518741, -0.0086413596171881248, 
    -0.0086383798244336965, -0.00862091477771618, -0.0085866831987356073, 
    -0.0085337870072279259, -0.0084607553370916622, -0.0083665379787815682, 
    -0.0082504874450480565, -0.0081123085256127551, -0.0079520036772735576, 
    -0.0077698259083273484, -0.0075662153346507605, -0.0073417645674039083, 
    -0.0070971879365313842, -0.0068333192815560996, -0.0065511107275614076, 
    -0.006251650730168647, -0.0059361904163774369, -0.0056061645584131398, 
    -0.0052632199318712533, -0.0049092333525095396, -0.0045463186386754629, 
    -0.0041768350518972073, -0.0038033684250816562, -0.0034287018713903723, 
    -0.0030557552268247966, -0.0026875258719335723, -0.0023269973039203337, 
    -0.0019770561264329852, -0.0016404265365240862, -0.0013196022625655193, 
    -0.0010167976032940038, -0.0007339180041891131, -0.000472542623179582, 
    -0.00023392009680275633, -1.8969346562033276e-05, 0.00017171061991712799, 
    0.00033782053775971454, 0.00047935325287258091, 0.00059657714772596009, 
    0.00069000897845613749, 0.00076039029273744995, 0.00080865609478763167, 
    0.00083589830345935775, 0.00084334092464505859, 0.00083230835283835632, 
    0.00080420549419943474, 0.00076050169713301799, 0.00070271615879445213, 
    0.00063241670765698727, 0.00055120565357862496, 0.00046070453801411708, 
    0.0003625460005722039, 0.00025834302611601573, 0.00014968411606776683, 
    3.8087964718507922e-05, -7.5012245232456228e-05, -0.00018829537127627955, 
    -0.00030056375446763518, -0.00041073206638693542, 
    -0.00051780939361192933, -0.00062086110575698629, 
    -0.00071898172994247695, -0.00081128851482978076, 
    -0.00089692035486259466, -0.0009750644871919478, -0.0010450000249517071, 
    -0.0011061246378871563, -0.0011580061520664465, -0.0012004149188367989, 
    -0.0012333299150795697, -0.0012569541672215838, -0.0012716794297064822, 
    -0.0012780509485549433, -0.0012767206461432065, -0.0012683777040920438, 
    -0.0012536881596839609, -0.0012332426734302478, -0.0012075288728293238, 
    -0.0011769139336680861, -0.0011416560231089902, -0.0011019252722846891, 
    -0.0010578433753771239, -0.0010095134503058151, -0.00095705972827696295, 
    -0.00090066083858129833, -0.00084057326816434561, 
    -0.00077715168032664486, -0.00071085797419248727, 
    -0.00064226574315716443, -0.00057205578476720415, 
    -0.00050099132492198971, -0.00042989949340494968, 
    -0.00035962588064417024, -0.00029100720026189791, -0.0002248242373598645, 
    -0.00016178475714500153, -0.00010249893687621628, 
    -4.7474908230635271e-05, 2.8854188455923208e-06, 4.8288846544642609e-05, 
    8.8567868738528063e-05, 0.00012370389937726143, 0.00015387067178302695, 
    0.00017947255198789394, 0.00020117832435871962, 0.00021995307581279143, 
    0.00023705352812273343, 0.00025399800989938775, 0.00027251035184082471, 
    0.00029443980189851853, 0.00032167401887461529, 0.00035605223309477242, 
    0.00039928151176207339, 0.00045287091069936517, 0.00051808285618574329, 
    0.00059587934378291935, 0.00068689959078887088, 0.00079142774476187352, 
    0.00090938209443527191, 0.001040305322526274, 0.0011833758006307158, 
    0.0013374115443002983, 0.0015009071892073747, 0.0016720722780020705, 
    0.0018488916470161235, 0.0020291902365099806, 0.0022106999451434869, 
    0.0023911305129792077, 0.00256822727674977, 0.0027398361462387237, 
    0.0029039405216733202, 0.0030587136697272604, 0.0032025428094982137, 
    0.0033340549760521891, 0.003452127654228327, 0.0035558951887257116, 
    0.0036447458792487823, 0.0037183286991384111, 0.0037765479107911733, 
    0.0038195747264627897, 0.0038478267070775861, 0.0038619729136015546, 
    0.0038628908779874569, 0.0038516350924949561, 0.0038293910050250547, 
    0.0037974256356232508, 0.0037570419067660303, 0.0037095415857614339, 
    0.0036561951124081944, 0.0035981943206356551, 0.0035366172571633901, 
    0.0034723823925522654, 0.0034061912631965507, 0.0033384914801457832, 
    0.0032694472057087053, 0.0031989487842885131, 0.0031266414233987717, 
    0.003051992412546133, 0.0029743552081050754, 0.0028930493620201673, 
    0.002807382926000281, 0.0027166564018899549, 0.0026201339809446503, 
    0.002516996535468509, 0.0024063097235017469, 0.0022870064301262105, 
    0.0021578891113700339, 0.0020176429812192448, 0.0018648474834042116, 
    0.0016980202931850543, 0.0015156618839197397, 0.0013163247176791904, 
    0.0010986852265725733, 0.00086162522195439267, 0.00060430555985488551, 
    0.00032622302901411007, 2.7234700405763719e-05, -0.00029243230016424667, 
    -0.00063220874213484879, -0.00099120802294150258, -0.001368279226073013, 
    -0.0017620195954761787, -0.0021707974472971016, -0.0025927440220768513, 
    -0.0030257506018811328, -0.0034674491597636702, -0.0039152078663313959, 
    -0.0043661150952787548, -0.0048169794868499847, -0.0052643321803337801, 
    -0.0057044603431263812, -0.0061334248519028965, -0.0065471232946430306, 
    -0.0069413468258327261, -0.0073118564787453787, -0.0076544746342292296, 
    -0.0079651838687363353, -0.0082402354249170671, -0.0084762537319975663, 
    -0.008670328961533422, -0.0088201014783933079, -0.0089238077242323553, 
    -0.0089803133017339089, -0.0089891284508144265, -0.0089503978212983823, 
    -0.0088648986537346094, -0.008733995459800319, -0.0085595994220461716, 
    -0.0083441050346307818, -0.0080903247941191449, -0.0078014111847289624, 
    -0.0074807751891306437, -0.0071320093381303943, -0.0067588416415065109, 
    -0.0063651011741723178, -0.0059546988701701664, -0.0055316266270568019, 
    -0.0050999448316842617, -0.0046637652976307918, -0.0042272134566641341, 
    -0.003794385126366027, -0.003369272917524581, -0.0029557074537598089, 
    -0.0025572775087088061, -0.0021772723053529799, -0.0018186219040784253, 
    -0.0014838503192667945, -0.0011750702089868719, -0.00089398889966448361, 
    -0.00064196680910142518, -0.00042008365218346318, 
    -0.00022920690059251281, -7.0032970795381186e-05, 5.6906381823571797e-05, 
    0.00015129171490755179, 0.00021309366202777106, 0.00024267139729432046, 
    0.00024085949726569201, 0.00020901437182175512, 0.00014901695670743742, 
    6.3228168631383188e-05, -4.5600560323383284e-05, -0.00017443661500779936, 
    -0.00032007458619348042, -0.00047921181161159694, 
    -0.00064850241923307232, -0.00082455948731792971, -0.0010039522088279038, 
    -0.001183173646728639, -0.0013586110122117329, -0.0015265475326861969, 
    -0.0016831586513890377, -0.0018245624218968079, -0.0019469001554652272, 
    -0.0020464252050517405, -0.002119632688913047, -0.0021633904815188667, 
    -0.0021750819059359302, -0.0021527095377488958, -0.0020949898669720022, 
    -0.0020013904649982335, -0.0018721239958392705, -0.0017081479565380614, 
    -0.0015111338442527296, -0.0012834594909388942, -0.0010281800426400135, 
    -0.00074899769574776382, -0.0004502027237046288, -0.00013658831745946127, 
    0.00018664704996218463, 0.00051400846739783207, 0.00083982432433005356, 
    0.0011583455141526713, 0.0014638871316717623, 0.0017509447896851746, 
    0.00201431094261379, 0.0022492233306383798, 0.0024514593897219036, 
    0.0026174335996744296, 0.0027442781832848753, 0.0028298630726583049, 
    0.0028728147135798341, 0.0028725017808658147, 0.0028290045998017352, 
    0.0027430854369614472, 0.002616144671077061, 0.0024501781393673899, 
    0.0022477356313609469, 0.0020118899616045137, 0.0017461602044066234, 
    0.0014544648461019057, 0.0011410556285720011, 0.00081043942370974051, 
    0.00046732083428050754, 0.00011653183910307686, -0.00023702724623032953, 
    -0.00058844623009364949, -0.00093288308606158811, -0.0012656351577231806, 
    -0.0015822291280939657, -0.001878524529496962, -0.0021508225800275964, 
    -0.0023959932637768193, -0.0026115955226512118, -0.0027960032417120705, 
    -0.0029485172058621835, -0.0030694230737701596, -0.0031600082266869259, 
    -0.0032225301013591445, -0.0032601202116328471, -0.0032766585334512727, 
    -0.0032765896259758262, -0.0032647434863887505, -0.0032461484789460472, 
    -0.0032258354676330172, -0.0032086836266315851, -0.0031992716868075402, 
    -0.0032017929980389295, -0.0032199504425931983, -0.0032569215258124776, 
    -0.0033153089298514904, -0.0033970977011849651, -0.0035036428088155596, 
    -0.0036356472013569581, -0.0037931703505973613, -0.00397560694969268, 
    -0.0041817168914401615, -0.0044096590641229203, -0.0046570371226221713, 
    -0.0049209621813386352, -0.0051981500095280323, -0.0054850312175990486, 
    -0.0057778831520615848, -0.0060729601043705986, -0.0063666513349032033, 
    -0.0066556084232525566, -0.0069368737240004582, -0.0072079453169359483, 
    -0.0074668228103800752, -0.0077120117869317936, -0.0079424747751050476, 
    -0.0081576077535092106, -0.0083571860523513567, -0.0085413256373320038, 
    -0.0087104420863243076, -0.0088652155070202028, -0.0090065427908634435, 
    -0.0091354927941959124, -0.009253242786880984, -0.0093610481720557085, 
    -0.0094601655441548058, -0.009551796325653384, -0.0096370552429751212, 
    -0.0097168927740334966, -0.0097920646887133863, -0.0098631024754078245, 
    -0.0099302926013061857, -0.0099936944560447983, -0.010053152190620673, 
    -0.010108315527650999, -0.010158649513726843, -0.010203453835355708, 
    -0.010241900598250756, -0.010273051912023436, -0.010295875858919151, 
    -0.010309288282457887, -0.01031217195603657, -0.010303415666877841, 
    -0.01028194438465754, -0.010246784296514357, -0.010197132920091915, 
    -0.010132427695204612, -0.010052414321463504, -0.0099571908526777109, 
    -0.0098472024256309933, -0.0097232279720394256, -0.0095863111073801761, 
    -0.0094377250635410952, -0.0092789108448129223, -0.009111445113535897, 
    -0.0089370162231049554, -0.0087573878950448995, -0.0085743686730211394, 
    -0.0083897790549994737, -0.0082053509871734664, -0.0080226783401159598, 
    -0.0078431385775499813, -0.0076678221228029565, -0.0074974917839986588, 
    -0.0073325796783632637, -0.0071731773368095622, -0.007019103989118855, 
    -0.0068699697520149729, -0.0067252440446277373, -0.0065843673092809765, 
    -0.0064468011872243292, -0.0063120721912437085, -0.0061797785631810499, 
    -0.0060495455067290978, -0.0059209506596295553, -0.0057934684818647377, 
    -0.0056663554479067547, -0.0055386005628493299, -0.005408867821624949, 
    -0.0052755091051528381, -0.0051365877263291381, -0.0049899740671361728, 
    -0.0048334393277283463, -0.0046647927098399074, -0.0044819915046098602, 
    -0.0042832760094168379, -0.0040672802186039079, -0.003833097676223726, 
    -0.0035803473083038167, -0.0033091795023665492, -0.0030202653001683969, 
    -0.0027147241939758354, -0.0023940523201674106, -0.0020600021020286815, 
    -0.0017144714793878137, -0.0013593957916143956, -0.00099665783441715817, 
    -0.00062806157285771706, -0.00025531136080767262, 0.00011994642816819828, 
    0.00049610908110175791, 0.00087154226631614177, 0.0012445422818545275, 
    0.0016132838262801175, 0.0019758133748787993, 0.0023300367891175779, 
    0.0026737178679537132, 0.0030045511976522694, 0.0033201987160917366, 
    0.0036184058910510705, 0.0038970680799544359, 0.0041543112272008249, 
    0.004388607886164974, 0.0045988817095474121, 0.004784584337978133, 
    0.0049458290630948146, 0.0050834712998025014, 0.0051991917136382012, 
    0.0052954967465293976, 0.00537557948961592, 0.0054430080727766476, 
    0.0055011754931902036, 0.00555269593670154, 0.0055988690066994971, 
    0.005639437158337186, 0.0056725945604279111, 0.0056952816692221759, 
    0.0057035968727201011, 0.0056932259632846809, 0.0056598483305965574, 
    0.0055995181911258499, 0.0055088966579999168, 0.0053854811644442075, 
    0.0052276306129224867, 0.0050346474873932279, 0.0048066575412489716, 
    0.0045446228983321733, 0.004250258966001081, 0.0039260055084987628, 
    0.0035750080511283227, 0.0032010495562493193, 0.0028084571236676051, 
    0.0024019949363604529, 0.0019867280109374811, 0.0015678541796861347, 
    0.001150533380246921, 0.0007397055830980372, 0.00033989550191180855, 
    -4.4950868491225424e-05, -0.00041160708060765556, 
    -0.00075764332997579681, -0.001081460472724992, -0.0013822265655770189, 
    -0.0016597707807184604, -0.0019144068017272378, -0.0021467211836905396, 
    -0.0023574100116369465, -0.0025470281501843903, -0.0027158981388518857, 
    -0.0028640001097639534, -0.0029909090358237922, -0.0030957876699355125, 
    -0.0031774043812737704, -0.0032341293703434301, -0.003264041386338051, 
    -0.0032649649831825132, -0.0032345863463385245, -0.0031705241601648962, 
    -0.0030704330715635932, -0.0029320719379318165, -0.0027534295908516657, 
    -0.0025328144558949659, -0.0022689501589174665, -0.0019610577854030169, 
    -0.0016088858599663152, -0.0012127240549996816, -0.00077341418197731889, 
    -0.00029232179615637207, 0.00022862946117526757, 0.00078698973948865822, 
    0.0013797541659949714, 0.0020033222754559758, 0.0026535139060247519, 
    0.0033255542978653462, 0.0040140846649932335, 0.0047132872555515626, 
    0.0054169251081142853, 0.0061184973617545539, 0.0068114556131756276, 
    0.0074894163568419818, 0.0081464010338037074, 0.0087770526392312361, 
    0.0093768352972620067, 0.0099421313968909159, 0.010470223244534168, 
    0.010959202125750918, 0.011407818373227968, 0.01181524476275372, 
    0.01218087683298563, 0.012504160271717052, 0.012784313820583006, 
    0.013020267163829398, 0.013210524174109603, 0.013353228548703484, 
    0.013446433605419, 0.01348849024810298, 0.013478451704162347, 
    0.01341661726400601, 0.013304847946909427, 0.013146812935068647, 
    0.012948132552795737, 0.012716252593888939, 0.012460259925561625, 
    0.012190491394248592, 0.011918107703712839, 0.011654553093617546, 
    0.011410963972818527, 0.011197659217855061, 0.011023654045837198, 
    0.010896302555674165, 0.010821088774124916, 0.010801580525128704, 
    0.010839493275016552, 0.010934863127453148, 0.011086191335018545, 
    0.011290639707746068, 0.01154421681386387, 0.011841798541577827, 
    0.012177379448521427, 0.012544061080940321, 0.012934055481950601, 
    0.013338601375684008, 0.013747784912453405, 0.014150396971100893, 
    0.014533802619122327, 0.014884114349904219, 0.015186366221876567, 
    0.015424905369374671, 0.015583991885637442, 0.015648374866298938, 
    0.01560395816991612, 0.015438419061265111, 0.015141757982584322, 
    0.014706615233556012, 0.014128453390013385, 0.013405538911713718, 
    0.012538687963738323, 0.011531093604708649, 0.010388105780091162, 
    0.0091171215812570275, 0.0077278460586299265, 0.0062324992365505056, 
    0.0046458911813602316, 0.0029854461262074803, 0.0012708401865238977, 
    -0.00047668052498866229, -0.0022350061650645544, -0.0039823279357876773, 
    -0.0056980509126820051, -0.0073638491586766504, -0.008964390396501435, 
    -0.010488073203007922, -0.011927286078769113, -0.013278428304263739, 
    -0.014541937832184144, -0.015721850342932397, -0.016825198413148643, 
    -0.01786159566981934, -0.018842284912042456, -0.019779440728412812, 
    -0.020685330277757614, -0.021571338084710911, -0.022446939376162069, 
    -0.023318779660560739, -0.024190053135333268, -0.025059843721441349, 
    -0.025922964787365055, -0.026770451377716446, -0.027590002500718167, 
    -0.028367239446743353, -0.029086928259038101, -0.029733815187922435, 
    -0.030293714954195083, -0.03075460607203425, -0.031106408865280585, 
    -0.031341788445253281, -0.031456244990441688,
  // Fqt-Na(5, 0-1999)
    1, 0.9965599533218914, 0.98633114227439644, 0.96958230314595195, 
    0.94674512482704054, 0.91839180889223337, 0.88520647900824689, 
    0.8479528115856575, 0.80744031621606804, 0.76449156840708066, 
    0.71991233685957268, 0.6744660322565792, 0.62885338662664247, 
    0.58369774740673297, 0.53953588366007521, 0.49681387808914196, 
    0.45588739857488086, 0.41702553441409773, 0.38041727375099371, 
    0.34617981761175881, 0.31436791687765514, 0.284983600438872, 
    0.25798576187548927, 0.23329920735627649, 0.21082293222230861, 
    0.19043743734665006, 0.17201104372636189, 0.1554051885035522, 
    0.14047873764141566, 0.12709140254455079, 0.11510635233120306, 
    0.1043921363428789, 0.094824038333605434, 0.086284960298451813, 
    0.078665941887143473, 0.071866390850303857, 0.065794101900841784, 
    0.060365118731880198, 0.055503475151018937, 0.05114087286677612, 
    0.047216288500892219, 0.043675562848348393, 0.040470947072414838, 
    0.037560645867381059, 0.034908328195078289, 0.032482632949416758, 
    0.030256669746918142, 0.028207515918353042, 0.026315725388558309, 
    0.024564850933387512, 0.022940986773443462, 0.02143235043967421, 
    0.020028901310768902, 0.018722010810583608, 0.017504188664676405, 
    0.016368862684788224, 0.015310220606611958, 0.014323104369539432, 
    0.013402941547609388, 0.012545723501776872, 0.011747981563657171, 
    0.011006779437550055, 0.01031968654260795, 0.0096847309799695681, 
    0.0091003258560021383, 0.0085651730771212718, 0.008078128411298199, 
    0.0076380609643246925, 0.0072436801119566251, 0.0068933743838192167, 
    0.0065850678324588605, 0.0063161069499981471, 0.0060831928039950366, 
    0.0058823684463705722, 0.0057090687963676128, 0.0055582168223604631, 
    0.0054243758313213802, 0.0053019352380704963, 0.0051853204822515497, 
    0.0050692125759659668, 0.0049487490781419188, 0.0048197083987463517, 
    0.0046786489314104623, 0.0045229996842730495, 0.0043510981627964389, 
    0.0041621748660575627, 0.0039562933221902862, 0.0037342561137334207, 
    0.0034974831227859815, 0.0032478730166665584, 0.0029876790028064782, 
    0.0027193748546249542, 0.0024455413794231265, 0.002168762030696349, 
    0.0018915242616729399, 0.0016161358774598312, 0.0013446588095645704, 
    0.0010788545245808032, 0.00082014567881965521, 0.00056959998293112132, 
    0.0003279291307348256, 9.549341429120631e-05, -0.00012767733395283598, 
    -0.00034185442482577856, -0.00054757211827370427, -0.0007455829555355906, 
    -0.000936802262411684, -0.0011222434934712458, -0.0013029439408167615, 
    -0.0014798749081516445, -0.0016538429435434185, -0.0018253873241434327, 
    -0.001994674339360061, -0.0021614123351596294, -0.0023247821142558561, 
    -0.0024834110319226664, -0.0026353791674091731, -0.0027782821675796216, 
    -0.0029093236631618775, -0.0030254427352701665, -0.0031234646719801125, 
    -0.003200259598852465, -0.0032529053654542332, -0.0032788322745894139, 
    -0.0032759575437030439, -0.0032427886816972095, -0.0031784870760141653, 
    -0.0030829043662007867, -0.0029565780848190412, -0.00280069506944972, 
    -0.0026170367660135322, -0.0024079011736341154, -0.0021760237673952017, 
    -0.0019244895488533405, -0.0016566442555574585, -0.001376012796097539, 
    -0.0010862092324722453, -0.00079085997033495365, -0.00049353618336918945, 
    -0.00019768716236216591, 9.3404518213000942e-05, 0.00037666622986269339, 
    0.00064926139592294335, 0.00090861005721042825, 0.0011524006283761741, 
    0.0013785967638423439, 0.0015854425104762338, 0.0017714568541037114, 
    0.0019354301440475817, 0.0020764142289237085, 0.0021937113979146198, 
    0.0022868552483668041, 0.0023556130502949786, 0.0023999880906037576, 
    0.0024202466511723062, 0.0024169522945023149, 0.0023910088996683611, 
    0.0023436973335506459, 0.0022766854755895999, 0.0021920138836110351, 
    0.0020920579778730191, 0.0019794641908234146, 0.0018570816671741085, 
    0.001727885047526744, 0.0015949000619526132, 0.0014611261133510663, 
    0.0013294633355625347, 0.0012026354269550276, 0.0010831255859523338, 
    0.00097311140304946308, 0.00087441907208565795, 0.000788495379543589, 
    0.0007163868757939537, 0.00065873338162604966, 0.00061576693745714578, 
    0.00058730775075658995, 0.00057277543938806291, 0.00057119848469155965, 
    0.00058123953989738407, 0.00060123228871527623, 0.00062922807996433606, 
    0.00066306653774874248, 0.00070044877377939635, 0.00073904405190635953, 
    0.00077659391999803274, 0.00081103699843422907, 0.00084062198581158606, 
    0.0008640021296652075, 0.00088031227024204419, 0.00088920225530523145, 
    0.00089083574448451546, 0.0008858455322773998, 0.00087526259357683289, 
    0.00086041417314993449, 0.00084281667414960661, 0.00082406800034161428, 
    0.00080574052629506557, 0.00078929987450875743, 0.00077601891452396292, 
    0.0007669159310098718, 0.00076270799242509442, 0.00076378117458817004, 
    0.00077018110280583773, 0.00078162271520250718, 0.00079751323150558263, 
    0.00081699167806045228, 0.00083898691413261813, 0.00086227148042547345, 
    0.00088552884968647278, 0.0009074186585945823, 0.00092663699973632627, 
    0.00094197026206512316, 0.00095234838194273395, 0.00095688413235303811, 
    0.00095490826790531238, 0.00094599786702073739, 0.00092999355252290508, 
    0.00090700837458870614, 0.00087741491504141631, 0.00084182427272026946, 
    0.00080104286544336624, 0.00075600892006364015, 0.00070772223114676117, 
    0.00065716131894427124, 0.00060519556543509013, 0.000552501163634773, 
    0.0004994872167616573, 0.00044623057727805862, 0.00039243975108881957, 
    0.00033744353044129981, 0.00028020944715926037, 0.00021940014344280637, 
    0.00015345107805200478, 8.0674237066875008e-05, -6.3381114652748824e-07, 
    -9.2072142342031617e-05, -0.00019503364310040062, -0.0003106092833669691, 
    -0.00043952026035740213, -0.00058206488594049932, 
    -0.00073808593459977374, -0.00090696470225508211, -0.0010876361860924471, 
    -0.0012786265225224504, -0.0014781149985995999, -0.0016840061001513825, 
    -0.0018940199223698496, -0.002105778163410918, -0.0023168860428623064, 
    -0.0025250035369176818, -0.0027279021683117282, -0.002923516066379632, 
    -0.0031099762939181615, -0.003285644786935269, -0.0034491384726669711, 
    -0.0035993468071586756, -0.0037354384051754542, -0.0038568570691986017, 
    -0.0039633084978089863, -0.0040547363463709048, -0.0041312882252072932, 
    -0.0041932877558846712, -0.0042412005325726948, -0.0042756182790458222, 
    -0.0042972403568941062, -0.004306860640742283, -0.0043053450837789616, 
    -0.0042935978397993799, -0.0042725139868919643, -0.0042429119944689267, 
    -0.0042054707814515296, -0.0041606560230010746, -0.0041086661565549361, 
    -0.0040493905186121818, -0.0039823949681079005, -0.0039069277933826297, 
    -0.0038219611399806035, -0.0037262520013652592, -0.0036184325918287895, 
    -0.0034971112888779353, -0.0033609921769672574, -0.0032089940275244764, 
    -0.0030403636753292191, -0.0028547779300764002, -0.0026524268797423734, 
    -0.0024340707068485996, -0.0022010691009723389, -0.001955374401440287, 
    -0.0016995036236320915, -0.0014364735500908962, -0.0011697228222593303, 
    -0.00090300991739918502, -0.00064029646674387364, 
    -0.00038562161920763715, -0.00014297719576859217, 8.3810384690549678e-05, 
    0.00029119201383139373, 0.00047598150300053813, 0.00063542212920543678, 
    0.00076723123020133342, 0.00086962458056445962, 0.00094132075938743124, 
    0.00098153189516654083, 0.0009899449171703093, 0.00096669524187455874, 
    0.0009123341158999473, 0.00082779226460402775, 0.00071434591412294207, 
    0.00057358530941091078, 0.0004073763702162127, 0.00021783375717060932, 
    7.2727734843492808e-06, -0.00022184219865454326, -0.00046695920063231255, 
    -0.00072550659486964367, -0.00099495234081184349, -0.0012728526356286403, 
    -0.0015568831096603507, -0.0018448486227123034, -0.0021346756107297978, 
    -0.0024243938787699257, -0.0027121172339087231, -0.0029960252441245099, 
    -0.0032743637202140284, -0.0035454612721317236, -0.0038077473370558318, 
    -0.0040597896508717873, -0.0043003056916780446, -0.0045281793619401205, 
    -0.0047424363023736808, -0.0049422037684030947, -0.0051266408824132597, 
    -0.0052948557177857581, -0.0054458296359556502, -0.005578348262645025, 
    -0.0056909748203180528, -0.0057820569958551594, -0.0058497851319691792, 
    -0.0058922843374497923, -0.0059077362703136025, -0.0058945129350661098, 
    -0.0058513072279160333, -0.0057772480444241072, -0.0056719910816555768, 
    -0.0055357828622520002, -0.005369481887551414, -0.0051745642173876023, 
    -0.0049530812782544037, -0.0047076051008881244, -0.0044411381380402796, 
    -0.0041570156091651073, -0.0038587858452961712, -0.0035500931852558023, 
    -0.0032345517456610243, -0.0029156450912109226, -0.0025966329315190379, 
    -0.0022804834545377098, -0.0019698170882194062, -0.0016668600087848501, 
    -0.0013734108631496787, -0.0010908096044731572, -0.00081992012419346175, 
    -0.00056112629114141339, -0.00031434623818600474, 
    -7.9065078872720762e-05, 0.00014560802447596263, 0.00036087388338437297, 
    0.00056816245352597078, 0.00076905300979336676, 0.00096519661936812957, 
    0.0011582522752101691, 0.0013498358922643422, 0.0015414852206854994, 
    0.0017346388415028491, 0.0019306281012766205, 0.0021306833042835003, 
    0.0023359341998844788, 0.0025474184715200874, 0.0027660676134920151, 
    0.0029926840289923162, 0.0032279000513520638, 0.0034721176678140027, 
    0.0037254442996174173, 0.0039876205264370076, 0.0042579589495129128, 
    0.0045352988389806169, 0.0048179941780565044, 0.0051039280034832196, 
    0.0053905683716357093, 0.0056750455984372165, 0.0059542566949586564, 
    0.0062249746754747927, 0.0064839675506693766, 0.0067281143141998453, 
    0.0069545145158703492, 0.0071605914200298772, 0.0073441730315113862, 
    0.0075035585839213952, 0.0076375549579648571, 0.0077454860197756466, 
    0.0078271752945602343, 0.0078828994115451648, 0.0079133325004700807, 
    0.0079194705607164798, 0.0079025579091358926, 0.0078640128665412312, 
    0.0078053599768764005, 0.007728172742593865, 0.007634017929829701, 
    0.0075244214892493111, 0.0074008396897897715, 0.0072646481578923644, 
    0.0071171444902706459, 0.0069595676969188922, 0.0067931275221538891, 
    0.0066190518112015668, 0.0064386203348788841, 0.0062531991022339358, 
    0.0060642465435163471, 0.0058733024850943158, 0.0056819429544326897, 
    0.0054917195731065396, 0.0053040773338655922, 0.0051202717908066138, 
    0.0049412863824090519, 0.0047677660774669934, 0.0045999692874210112, 
    0.0044377484187352913, 0.0042805500651325141, 0.0041274446245855943, 
    0.0039771602619216228, 0.0038281325329998202, 0.003678551075425739, 
    0.00352640865641108, 0.0033695542987373906, 0.0032057586749415605, 
    0.0030327945305534802, 0.002848545725550444, 0.0026511375242674919, 
    0.0024390788370589498, 0.0022114103208244907, 0.0019678278956416378, 
    0.0017087692820847732, 0.0014354436433576725, 0.0011498028080173424, 
    0.00085445264667592246, 0.00055251399089925764, 0.00024744711841095468, 
    -5.7141279671727075e-05, -0.00035769108289970418, 
    -0.00065085752617906659, -0.00093364847682583991, -0.0012035287386733063, 
    -0.001458500935861093, -0.001697166655131322, -0.0019187707954881345, 
    -0.0021232182021618359, -0.002311048344923496, -0.0024833571108895842, 
    -0.0026416729457666242, -0.002787788964460366, -0.0029235848028034248, 
    -0.0030508277936796887, -0.0031710052282968031, -0.0032851734491931234, 
    -0.0033938415117701292, -0.0034968980477224107, -0.0035935814269288705, 
    -0.0036824978064890481, -0.0037616853185467869, -0.0038287269611228429, 
    -0.003880899922968336, -0.0039153603155365488, -0.0039293389941747877, 
    -0.0039203367150609592, -0.0038863124853276932, -0.0038258379624932569, 
    -0.0037382210130343335, -0.003623584467272832, -0.0034829005552195797, 
    -0.0033179757815887979, -0.0031313987092653145, -0.0029264551975314757, 
    -0.002707023289467445, -0.0024774482599495338, -0.0022424229761555605, 
    -0.0020068615382132439, -0.0017757849690538574, -0.001554213712854018, 
    -0.0013470608605910637, -0.00115903490357455, -0.00099454406875525408, 
    -0.00085758697909198134, -0.00075165877213213643, 
    -0.00067964922216919249, -0.00064374808044273752, 
    -0.00064536296141360716, -0.00068503959454210427, 
    -0.00076239861433807072, -0.00087608840008657988, -0.0010237770690213731, 
    -0.0012021670071365642, -0.0014070661164926079, -0.0016334890340282487, 
    -0.0018758036288830278, -0.0021278934395799207, -0.0023833405630215672, 
    -0.0026356036728008422, -0.002878207938934515, -0.0031049243026690016, 
    -0.0033099479663438935, -0.0034880722519641744, -0.0036348469818095414, 
    -0.0037467214598353085, -0.0038211527895940416, -0.0038566800134725893, 
    -0.0038529433280664557, -0.0038106599812321889, -0.003731548729458026, 
    -0.0036182187845002658, -0.0034740355028100825, -0.0033029681652302243, 
    -0.0031094432720775423, -0.0028982065417153427, -0.0026741996817239602, 
    -0.0024424527368564373, -0.0022079914325744982, -0.0019757629037749072, 
    -0.001750556665480821, -0.0015369343272401013, -0.0013391477675976497, 
    -0.001161062986881328, -0.0010060785164144079, -0.00087705338153729853, 
    -0.00077622719265561129, -0.00070515431478588761, 
    -0.00066463916292943033, -0.00065469991532148973, 
    -0.00067454989089759157, -0.00072261025728347626, 
    -0.00079655233196827856, -0.00089335964297714314, -0.0010094202353714541, 
    -0.0011406347597750768, -0.0012825398637189463, -0.0014304477298356672, 
    -0.0015795856907283774, -0.0017252443596483971, -0.0018629163609950759, 
    -0.0019884263288521701, -0.0020980386906727681, -0.0021885381599605343, 
    -0.0022572798394732058, -0.0023022064175341975, -0.002321828754662289, 
    -0.0023151798359980144, -0.0022817417247325473, -0.0022213739647296477, 
    -0.0021342325344419814, -0.0020207089720796225, -0.0018813786106242625, 
    -0.0017169679318418786, -0.0015283374929624738, -0.001316471643257878, 
    -0.0010824803128268827, -0.00082760688595783253, -0.00055324326952488746, 
    -0.00026094554169377496, 4.7547444328792344e-05, 0.00037028928124309207, 
    0.00070510931630746523, 0.0010495950287303744, 0.0014010803486632201, 
    0.0017566441730084855, 0.0021131136384073112, 0.0024670762540675729, 
    0.0028149038335809201, 0.0031527809228076753, 0.0034767535492335228, 
    0.0037827833182952678, 0.0040668244203081547, 0.004324903259114817, 
    0.0045532129054283322, 0.0047482160150707359, 0.0049067446151524466, 
    0.0050261042327444574, 0.0051041727893319424, 0.0051394806599908962, 
    0.0051312863919981879, 0.0050796243654147484, 0.0049853280720282044, 
    0.0048500359886246699, 0.0046761612282218657, 0.0044668438704146291, 
    0.0042258681674106728, 0.0039575577260879185, 0.0036666452178765407, 
    0.0033581171301805633, 0.0030370496344547409, 0.0027084380310138383, 
    0.0023770447925385569, 0.0020472602909679658, 0.0017230026883780032, 
    0.0014076410514791164, 0.0011039697694025076, 0.0008142069721109803, 
    0.00054003023631665076, 0.0002826338845548788, 4.2804963796723872e-05, 
    -0.00017899483866374785, -0.00038254910681091101, -0.0005678096936868281, 
    -0.00073483336796710888, -0.00088372839438123759, -0.0010146207685453536, 
    -0.0011276321745178838, -0.0012228765309903783, -0.0013004659392981551, 
    -0.0013605334923901932, -0.0014032620269642285, -0.0014289201689077686, 
    -0.0014378819842292513, -0.001430656517828949, -0.0014079000110444519, 
    -0.0013704165418469733, -0.0013191515590732002, -0.0012551845398417953, 
    -0.0011797129994568704, -0.0010940372988971154, -0.00099954255893896365, 
    -0.00089767967446098269, -0.00078994699010572508, 
    -0.00067787702755437861, -0.00056302772012266659, 
    -0.00044696493827765587, -0.00033126046579756382, 
    -0.00021747367038639942, -0.00010713597573548623, 
    -1.7292188156013363e-06, 9.7346112126304063e-05, 0.00018881254581857665, 
    0.00027156041306687694, 0.00034470506342665352, 0.00040763950122078515, 
    0.00046009357376269991, 0.00050218400892346042, 0.00053447054424108969, 
    0.00055798116942973948, 0.00057423059116558557, 0.00058520181220180032, 
    0.00059330191862027649, 0.00060128555576699364, 0.00061214871059613409, 
    0.00062900472084461952, 0.00065494839270546616, 0.00069291208757572538, 
    0.00074553025614046008, 0.00081501468305278011, 0.00090304562461067904, 
    0.0010106839553810601, 0.0011383070566003334, 0.0012855741138734693, 
    0.0014514198209971763, 0.0016340830549532097, 0.0018311674805483388, 
    0.0020397371169925947, 0.002256446836833547, 0.0024776900762120677, 
    0.0026997624270919088, 0.002919025968859265, 0.0031320532434006838, 
    0.0033357407320474455, 0.0035273893526023802, 0.0037047371794994405, 
    0.0038659557736186829, 0.0040096045712347478, 0.0041345577810171039, 
    0.0042399134602502482, 0.0043248881825417723, 0.0043887181489326611, 
    0.0044305702706698268, 0.0044494785218110134, 0.004444313512857, 
    0.0044138001683563686, 0.0043565768929490828, 0.0042712852367232197, 
    0.0041566892423182547, 0.0040118046474348808, 0.0038360375631776161, 
    0.0036293199698197247, 0.0033922367057983259, 0.0031261340776306897, 
    0.0028331815347257604, 0.0025164007128225412, 0.0021796349917907873, 
    0.0018274757574385002, 0.0014651453727305846, 0.0010983382514251187, 
    0.00073303962814698787, 0.0003753166274832303, 3.111958086683932e-05, 
    -0.00029391004258624945, -0.00059459053775071287, 
    -0.00086631897096670226, -0.0011051494246142306, -0.0013078399996665009, 
    -0.0014718631468536422, -0.0015953982793159027, -0.0016773057735711488, 
    -0.0017171015109201122, -0.0017149292596963161, -0.001671527299952051, 
    -0.0015882112491531267, -0.0014668506279914507, -0.0013098457498561884, 
    -0.0011200981168841646, -0.00090096788284368609, -0.00065620915019553271, 
    -0.00038988415600213423, -0.00010626416759944822, 0.00019029117781216997, 
    0.00049545937933839551, 0.00080507942609786868, 0.0011152670932100734, 
    0.0014225175872100708, 0.0017237789151162029, 0.0020165061534623092, 
    0.0022986853820904075, 0.0025688254757197859, 0.0028259245974256008, 
    0.0030694096772431716, 0.0032990617457435813, 0.0035149374393263783, 
    0.0037172895158453043, 0.0039064909965421763, 0.0040829693061541893, 
    0.0042471482858073457, 0.0043993894948713775, 0.0045399543990163379, 
    0.0046689641120724419, 0.0047863766555315893, 0.0048919718767555954, 
    0.0049853484116666371, 0.0050659255879105334, 0.0051329428428916806, 
    0.0051854699378773685, 0.0052224132865311855, 0.0052425377893861452, 
    0.0052445086516702171, 0.0052269434692501591, 0.00518848683490848, 
    0.0051278919943471574, 0.0050441052871579364, 0.0049363508868697659, 
    0.0048042037132165795, 0.0046476470686600624, 0.0044671146469636028, 
    0.0042635189082164534, 0.0040382683125463493, 0.0037932625527051229, 
    0.0035308837183859829, 0.003253956824510385, 0.0029657009608985009, 
    0.0026696593949347893, 0.0023696153421687177, 0.0020694950834679328, 
    0.0017732755899989173, 0.0014848956628801878, 0.0012081727634683792, 
    0.00094673149966233248, 0.00070394520604019238, 0.00048287285589339188, 
    0.00028620911328117898, 0.00011623133304246986, -2.5250055594534825e-05, 
    -0.0001369314589336893, -0.00021805190750323248, -0.00026842042824371816, 
    -0.00028842978047972223, -0.00027906106059376551, 
    -0.00024188223226517201, -0.00017902228546778475, 
    -9.3142411180507391e-05, 1.2613577846582835e-05, 0.00013469285243550646, 
    0.00026922283881301791, 0.00041211978099679866, 0.00055921045195175237, 
    0.0007063617463046166, 0.00084960910586003187, 0.00098527475381755803, 
    0.0011100743000290313, 0.0012212072092338292, 0.001316427946570024, 
    0.0013940978320532114, 0.0014532213351837093, 0.0014934591529694122, 
    0.0015151257677917685, 0.0015191637404183285, 0.0015071025461968156, 
    0.001480996262643131, 0.0014433444565644404, 0.001396993564997485, 
    0.0013450200878072091, 0.0012906034546637931, 0.0012369050472144181, 
    0.0011869400483141448, 0.0011434742949789139, 0.0011089453967989484, 
    0.0010854142687983317, 0.0010745396153436604, 0.0010775771437192484, 
    0.00109539598456489, 0.0011285040645706477, 0.0011770676150947533, 
    0.0012409405516451109, 0.0013196885498793017, 0.0014126088591455354, 
    0.0015187569283766828, 0.0016369649696674562, 0.0017658690969827365, 
    0.0019039321297258957, 0.0020494596469682633, 0.0022006268246791845, 
    0.0023554975677837612, 0.0025120478991575617, 0.0026681926474028052, 
    0.0028218182295590049, 0.0029708147008116101, 0.0031131141246665971, 
    0.0032467297563067085, 0.0033697968884594401, 0.0034806152990321348, 
    0.0035776860539631105, 0.0036597503503530741, 0.0037258140430709527, 
    0.0037751721658218478, 0.0038074124734648936, 0.003822414645445465, 
    0.0038203260790193256, 0.0038015455527563792, 0.0037666863304364842, 
    0.0037165453824897195, 0.0036520713661314774, 0.0035743312967482853, 
    0.0034844863447819501, 0.003383757185698796, 0.0032733990866313629, 
    0.0031546734614860939, 0.0030288194427177118, 0.0028970245586134201, 
    0.002760399768575136, 0.002619951574407451, 0.0024765564162010836, 
    0.0023309411262903211, 0.0021836647520103317, 0.0020351083294892279, 
    0.0018854857530777079, 0.0017348656512748931, 0.0015832173456791442, 
    0.0014304813177100058, 0.0012766499073215091, 0.001121864008157389, 
    0.00096649992899492537, 0.00081125300670770802, 0.00065718102770977855, 
    0.00050572148452150581, 0.00035865449425747341, 0.00021801788463821255, 
    8.5982914383331169e-05, -3.5295420484683063e-05, -0.0001438426071794013, 
    -0.00023800547835991451, -0.00031656527271310035, 
    -0.00037880782451276285, -0.0004245562218664578, -0.00045416401511998747, 
    -0.0004684983631224565, -0.00046888325663066487, -0.00045704162756857473, 
    -0.00043501760782586299, -0.00040509027686360354, 
    -0.00036967232932780237, -0.0003312144713459354, -0.00029210167400059266, 
    -0.00025456635917952912, -0.00022061961079558427, 
    -0.00019199691055509231, -0.00017014329169927692, 
    -0.00015621474711054054, -0.00015110413308686357, 
    -0.00015547587997266144, -0.0001698076719876861, -0.00019441837361585084, 
    -0.00022949281037668273, -0.0002750898826329065, -0.0003311374034195468, 
    -0.00039742223158195417, -0.00047356816231388515, 
    -0.00055902978262381358, -0.00065308225226991148, 
    -0.00075482443563922898, -0.00086319188889681588, 
    -0.00097697975850112757, -0.0010948664018184092, -0.0012154503916803568, 
    -0.0013372871534900626, -0.001458930631383369, -0.0015789784795757478, 
    -0.0016961144453337821, -0.0018091486555854757, -0.001917050265433263, 
    -0.0020189752295075489, -0.0021142790221084311, -0.002202520718036784, 
    -0.002283446802279326, -0.0023569659175428689, -0.0024231110941931437, 
    -0.002481980989329917, -0.0025336981139084847, -0.0025783607050485621, 
    -0.0026160069320216349, -0.0026466078444683846, -0.0026700696972929479, 
    -0.0026862572663342043, -0.0026950242318487896, -0.0026962479228912436, 
    -0.0026898568382339896, -0.0026758531659377615, -0.0026543249053884699, 
    -0.0026254428232908296, -0.0025894412391972771, -0.0025465903258694153, 
    -0.0024971452538475178, -0.0024412909998011651, -0.0023790767380647269, 
    -0.0023103608338069419, -0.0022347739131479455, -0.0021517133370214641, 
    -0.0020603907034076603, -0.0019599105900053393, -0.0018493956621286767, 
    -0.0017281270588882232, -0.0015956749217752113, -0.001452010877921735, 
    -0.0012975709430886261, -0.0011332949515126111, -0.0009606194609546564, 
    -0.00078144466738712967, -0.00059808210423296546, 
    -0.00041317265264732936, -0.00022958971366642282, 
    -5.0324353184118915e-05, 0.00012162502464097284, 0.00028337097639681314, 
    0.00043222961559604117, 0.00056580560088791653, 0.0006820491429537362, 
    0.0007792980964255546, 0.00085631434440237094, 0.00091230483255843068, 
    0.00094694870825676126, 0.00096041323434924869, 0.0009533611286634407, 
    0.00092693796159279331, 0.00088273521251468906, 0.00082273795211240241, 
    0.00074923779651797954, 0.00066474380565924611, 0.00057187842113620897, 
    0.00047327461753323422, 0.00037147805350020666, 0.00026886393809981847, 
    0.00016757662227411517, 6.947511550578981e-05, -2.3884749438082587e-05, 
    -0.00011126088767147478, -0.000191707781686084, -0.000264565151112188, 
    -0.0003294216157133941, -0.00038609293924684159, -0.00043459403043487235, 
    -0.00047511892532244395, -0.00050801320762838137, 
    -0.00053375188826382193, -0.00055291379387686392, 
    -0.00056615390849879248, -0.00057418332813326711, -0.0005777587073036751, 
    -0.00057767805638653811, -0.00057478824940774946, 
    -0.00056999002871595305, -0.000564237795702015, -0.0005585242507126669, 
    -0.00055385489134217834, -0.00055120620050802516, 
    -0.00055147759996991932, -0.00055543786638109576, 
    -0.00056367353544605771, -0.00057653492806820472, 
    -0.00059409947118612425, -0.00061613499644371092, -0.0006420794667414525, 
    -0.00067103447549053197, -0.00070176966862532165, -0.0007327450443750719, 
    -0.00076213748661022658, -0.00078789453309141143, 
    -0.00080778289879820649, -0.00081946932945064664, -0.0008206000711814429, 
    -0.00080889175094210565, -0.00078221989930831067, 
    -0.00073870251485082781, -0.00067677728961388196, 
    -0.00059527144055406022, -0.00049346100468893744, 
    -0.00037113240708056461, -0.00022863749060362041, 
    -6.6939515463148203e-05, 0.00011234094193882072, 0.00030691441598681719, 
    0.00051382768924895794, 0.00072950709205259765, 0.00094983575235394716, 
    0.0011702740717531765, 0.0013860055097895136, 0.001592122620367324, 
    0.001783826967105485, 0.001956643808788355, 0.0021066354252177633, 
    0.0022305924712702706, 0.0023261925820470784, 0.0023921018287793544, 
    0.002428019441548513, 0.0024346537784845582, 0.0024136322631489473, 
    0.0023673652967315714, 0.0022988668530497768, 0.0022115531381982066, 
    0.0021090419457363402, 0.0019949536655175419, 0.0018727402190296901, 
    0.0017455396118610208, 0.0016160720791699196, 0.0014865774106651284, 
    0.0013587868317035605, 0.0012339465311841059, 0.001112861908022897, 
    0.00099597560443034612, 0.00088344693077478469, 0.00077523611039859597, 
    0.00067116885354693624, 0.00057097939044403452, 0.00047433066256915809, 
    0.00038082501067536543, 0.00029000449078639585, 0.00020136012565016595, 
    0.00011436305660293775, 2.8501695888396932e-05, -5.6659775152582124e-05, 
    -0.00014142451048747707, -0.00022591101417517029, 
    -0.00031002705461773508, -0.000393452658771352, -0.00047563453727242355, 
    -0.0005557850370925487, -0.00063288331498716145, -0.00070568514727885161, 
    -0.00077273783083576641, -0.00083239581996626252, -0.0008828510106667839, 
    -0.00092216025996667318, -0.000948280843935655, -0.00095911776289326831, 
    -0.00095256195128933397, -0.00092655049237059639, 
    -0.00087912634255805282, -0.00080851145870468224, 
    -0.00071318891704355732, -0.00059198592960733572, 
    -0.00044414927770240146, -0.00026941911134742511, -6.807169620780013e-05, 
    0.00015904920450520257, 0.00041052882768659023, 0.00068440409973176527, 
    0.00097820826012244826, 0.0012890372699418606, 0.0016136336065761224, 
    0.0019484918568732081, 0.0022899586161329302, 0.0026343359206519347, 
    0.0029779638280878649, 0.0033172817031799184, 0.0036488721259856642, 
    0.0039694928392263237, 0.0042761102388354753, 0.0045659413064648791, 
    0.0048365132178797895, 0.0050857299646241624, 0.0053119424417004081, 
    0.0055140144035507165, 0.0056913830857475613, 0.0058440939142989498, 
    0.0059728247070817324, 0.0060788669116687557, 0.0061640938382895322, 
    0.0062308788838236926, 0.0062819987220162762, 0.0063204978747330096, 
    0.0063495355363756365, 0.0063722240232062712, 0.0063914729948171501, 
    0.0064098410916764896, 0.0064294227946391702, 0.0064517622677426048, 
    0.0064778123133228758, 0.006507935546478944, 0.0065419435467089782, 
    0.006579172035589183, 0.0066185787989997864, 0.0066588545681471592, 
    0.0066985225359296324, 0.0067360381565564056, 0.0067698652559637267, 
    0.0067985268320169016, 0.0068206367786065453, 0.0068349199204732411, 
    0.0068401999135443, 0.006835401332633266, 0.0068195270122243723, 
    0.006791655998070645, 0.0067509414191575558, 0.0066966217445085831, 
    0.0066280451124312474, 0.0065446937375262951, 0.0064462071450398853, 
    0.0063324083385319588, 0.0062032997562561087, 0.0060590583355169631, 
    0.0059000082507796479, 0.0057265820241685214, 0.0055392746166011177, 
    0.0053386016985046717, 0.005125058709184613, 0.0048991031401920725, 
    0.0046611441468550176, 0.0044115647514246254, 0.004150750570956022, 
    0.0038791379692712491, 0.0035972699781963886, 0.0033058468267758256, 
    0.0030057748635374799, 0.0026982069493681807, 0.0023845731807651204, 
    0.0020666083602094462, 0.0017463646656498768, 0.0014262119356727573, 
    0.0011088257748722895, 0.00079715130326902704, 0.00049435046583858099, 
    0.00020372777511105676, -7.1352084359104883e-05, -0.00032757038239653421, 
    -0.0005617576645995365, -0.00077099037220411133, -0.00095270102198914805, 
    -0.0011047666458689862, -0.001225599724885424, -0.0013142229933673657, 
    -0.0013703367164580654, -0.0013943568227272681, -0.0013874350755476955, 
    -0.0013514457583461833, -0.0012889399758287674, -0.0012030833784197463, 
    -0.0010975679632742005, -0.00097651460551060915, -0.00084437678318937054, 
    -0.00070582805796227911, -0.0005656648417413935, -0.00042870477546170691, 
    -0.00029967533371956403, -0.00018310529491876229, 
    -8.3202440773360296e-05, -3.7288371456711865e-06, 5.2123489132695666e-05, 
    8.1867383289607526e-05, 8.3839822659526812e-05, 5.7298118796583037e-05, 
    2.4963828697318474e-06, -7.9279816084228865e-05, -0.00018571437468749698, 
    -0.00031351988062341485, -0.00045852248966619426, 
    -0.00061578847015347077, -0.00077978888008744043, 
    -0.00094459161041753341, -0.0011040715572243108, -0.0012521338361234022, 
    -0.0013829501965925296, -0.0014911799350291605, -0.0015721849822338547, 
    -0.0016222156561459743, -0.0016385694691961122, -0.0016197087962819725, 
    -0.001565335809379685, -0.0014764144003287193, -0.0013551462716351393, 
    -0.0012049050600026919, -0.0010301238564489866, -0.00083615690131103135, 
    -0.00062910956074200479, -0.00041565667103414625, 
    -0.00020283903293262881, 2.152779718676373e-06, 0.00019219658815927308, 
    0.00036045876418148797, 0.00050061708592029808, 0.00060706937716438979, 
    0.0006751279421281848, 0.0007011625266449494, 0.00068272152352400557, 
    0.00061859298384517455, 0.00050881277219281358, 0.00035462361063712917, 
    0.00015838908661552095, -7.6534638921353496e-05, -0.00034595856493079875, 
    -0.00064503613953026623, -0.00096844906710537358, -0.0013105900418575005, 
    -0.001665729704810147, -0.0020281578016213926, -0.0023922939375065479, 
    -0.0027527636214295576, -0.0031044562260911868, -0.0034425625809705812, 
    -0.0037626031997841799, -0.0040604759516899907, -0.0043324987243234386, 
    -0.0045754594452267761, -0.0047866700842580821, -0.0049640079109171441, 
    -0.0051059475321090604, -0.0052115917000464876, -0.0052806863997178193, 
    -0.0053136251572694993, -0.0053114594797324969, -0.0052758855591229972, 
    -0.005209217194820058, -0.0051143241820561991, -0.0049945516004769666, 
    -0.0048536024173170267, -0.0046954108276930561, -0.0045239949144068462, 
    -0.0043433269193322872, -0.0041572068942800668, -0.0039691599869176464, 
    -0.0037823522333650102, -0.0035995298615842603, -0.0034229752277795292, 
    -0.0032544836873957287, -0.0030953652685269386, -0.0029464478229075533, 
    -0.0028080918664109391, -0.0026802168048605688, -0.0025623157562495043, 
    -0.0024534708862551441, -0.0023523733590033427, -0.0022573584290761879, 
    -0.0021664559083552199, -0.0020774579093392987, -0.0019880024663985613, 
    -0.0018956650976173404, -0.0017980531160831671, -0.0016928997085893847, 
    -0.0015781673807312205, -0.0014521423664701479, -0.0013135433281621354, 
    -0.0011616097586380383, -0.00099618087363583484, -0.00081775985664659723, 
    -0.00062754217391946339, -0.00042741752623787579, 
    -0.00021994392835664265, -8.2789434520066409e-06, 0.00020391723723156248, 
    0.00041261049543463418, 0.0006135479802379482, 0.00080242610087914311, 
    0.00097506292059515128, 0.0011275623859941701, 0.0012564737883226837, 
    0.0013589332161218462, 0.0014327906530331755, 0.0014767179406958548, 
    0.0014902951627145603, 0.001474063103781047, 0.0014295313654669188, 
    0.001359143190150797, 0.001266189522840193, 0.001154678693258462, 
    0.0010291636144518443, 0.00089455124654608394, 0.00075590841667586884, 
    0.00061826069773460689, 0.00048640564940822731, 0.00036474762395483795, 
    0.00025716315003183464, 0.0001668757215180328, 9.6377422329773694e-05, 
    4.7356858842971254e-05, 2.064695454411933e-05, 1.6177264983238884e-05, 
    3.2954380422338579e-05, 6.9031663433847406e-05, 0.00012154062529125975, 
    0.00018674783924212907, 0.00026018851665946414, 0.00033684999600719324, 
    0.00041139121041423464, 0.000478394639353562, 0.00053262931441329289, 
    0.00056929899040747444, 0.00058426867604947225, 0.00057424809566042779, 
    0.00053692089659861976, 0.00047102620501866246, 0.00037637838941365119, 
    0.00025384034567277444, 0.00010525056360711452, -6.6673176774388534e-05, 
    -0.00025847237437508219, -0.00046611128417484084, 
    -0.00068516655619357911, -0.00091103470946961394, -0.0011391454251860954, 
    -0.0013651588446166518, -0.0015851511645028175, -0.0017957600957301313, 
    -0.0019943016284016588, -0.0021788261837911512, -0.0023481470374980286, 
    -0.0025018143309909393, -0.0026400441020837601, -0.0027636194490578527, 
    -0.002873755213657272, -0.002971942173546641, -0.0030597893911590971, 
    -0.003138867485349423, -0.0032105590444199083, -0.0032759478372287078, 
    -0.0033357290692370336, -0.0033901661314975854, -0.0034390869292289261, 
    -0.0034819258293094825, -0.0035178105305461393, -0.003545680595721266, 
    -0.0035644101468302368, -0.0035729303582941064, -0.0035703075118719788, 
    -0.0035557872110583109, -0.0035287792641561472, -0.0034888106785797134, 
    -0.0034354330632110734, -0.0033681365064671251, -0.0032862825590798117, 
    -0.0031890884891478412, -0.0030756618778796556, -0.0029451003329369228, 
    -0.0027966534480867002, -0.0026298901655348299, -0.0024449055526590052, 
    -0.00224249484449784, -0.0020242905573444824, -0.0017928523532221229, 
    -0.0015516507755098138, -0.00130498729783227, -0.0010577986267041263, 
    -0.00081541313827265577, -0.00058324053784867842, 
    -0.00036644078265123825, -0.00016960715057192966, 3.5138023214937664e-06, 
    0.00015023294817595846, 0.00026904187051821825, 0.0003596374235246252, 
    0.00042286514499606856, 0.00046057819277039167, 0.00047544256593045145, 
    0.00047072336157793912, 0.000450043325296215, 0.00041717104198452852, 
    0.00037581513932583076, 0.0003294743895401019, 0.00028132252732581927, 
    0.00023414494301844432, 0.00019029923198862666, 0.00015172236856252002, 
    0.00011995588880069254, 9.6173563028919727e-05, 8.1227326913582264e-05, 
    7.5682932846648815e-05, 7.9851806774136678e-05, 9.3825187404532936e-05, 
    0.00011748768182030372, 0.00015051814626414368, 0.00019236742251451798, 
    0.00024222699951111765, 0.00029898229979800634, 0.00036114985907097978, 
    0.00042684621101745447, 0.00049374279544359329, 0.00055907307014993089, 
    0.0006196536013859332, 0.00067192994984183445, 0.00071207117140375544, 
    0.00073607481228648523, 0.00073991276641379854, 0.00071969521269580803, 
    0.00067185798315067414, 0.00059335546410473809, 0.00048184569634512734, 
    0.00033584405939788621, 0.00015484250778489302, -6.0615826967025946e-05, 
    -0.00030892245970547399, -0.00058744392855793106, 
    -0.00089259396357508421, -0.001219969203766006, -0.0015644894007461256, 
    -0.001920587050467592, -0.0022823785401096808, -0.0026438620308604039, 
    -0.0029990920618395657, -0.0033423398184285569, -0.0036682359807191679, 
    -0.0039718769743365264, -0.0042489350148106819, -0.0044957410158811776, 
    -0.0047093826225006142, -0.0048877990850874223, -0.005029854593259925, 
    -0.0051353971225247845, -0.005205277537047419, -0.0052413471409003768, 
    -0.0052464314298097843, -0.0052242795688061637, -0.0051794838978655965, 
    -0.0051173699347297468, -0.0050438356089732659, -0.0049651578457736113, 
    -0.004887770447037738, -0.0048180237011327849, -0.0047619421913061019, 
    -0.0047249805514479977, -0.0047118248046435088, -0.0047262071993830878, 
    -0.0047707773623707197, -0.0048470032795989966, -0.0049551043479388575, 
    -0.0050940067149747173, -0.0052613207015325689, -0.0054533794443183932, 
    -0.0056653003370107707, -0.0058911200619162834, -0.0061239950415977081, 
    -0.0063564727995417984, -0.0065807868127680481, -0.0067891706350000037, 
    -0.0069741578811935521, -0.0071288266413897725, -0.0072470001027548081, 
    -0.0073234023635159497, -0.007353770359842123, -0.0073349389261982431, 
    -0.0072648731169665595, -0.0071426670112462211, -0.0069684958723691846, 
    -0.0067435263901179689, -0.0064698053184918322, -0.0061501147521371919, 
    -0.0057878496426860479, -0.005386896944698529, -0.0049515343605112932, 
    -0.0044863328469091903, -0.0039960791058671723, -0.0034856910986952681, 
    -0.0029601625226451812, -0.0024245098946224118, -0.0018837540043371783, 
    -0.0013429085487419124, -0.0008069760632658414, -0.0002809173048796892, 
    0.00023038580031506666, 0.00072220786163978198, 0.0011900600983603296, 
    0.0016297890553158916, 0.0020376749268982961, 0.0024105460796901698, 
    0.0027458979618099483, 0.0030419987116811994, 0.0032979999887703957, 
    0.0035140140627389063, 0.0036911533286140201, 0.0038315348549322796, 
    0.0039382256153501572, 0.0040151313519740184, 0.0040668530885336115, 
    0.0040984846042601553, 0.0041154170500186018, 0.0041231204024517465, 
    0.0041269634532100892, 0.0041320453218388715, 0.0041430478572934111, 
    0.0041641368235041882, 0.0041988644191070616, 0.0042501117339334288, 
    0.0043200513157742471, 0.0044101181662674939, 0.0045210214742454, 
    0.0046527460476633283, 0.0048046164195682502, 0.0049753400223208561, 
    0.0051630848775567808, 0.0053655659757881309, 0.0055801135249239414, 
    0.0058037571213521745, 0.0060332807977955391, 0.0062652690428931894, 
    0.0064961294438875602, 0.0067221243156552002, 0.0069393929516820491, 
    0.0071439830888956803, 0.0073318967794297864, 0.0074991629055683566, 
    0.0076419068459705648, 0.0077564440623412584, 0.0078393510637804493, 
    0.007887549854384588, 0.0078984144552248989, 0.0078698772939670997, 
    0.0078005874808654355, 0.0076900838348157256, 0.007538956973685086, 
    0.0073489632471964057, 0.0071230729750013161, 0.0068653915760095979, 
    0.00658101862370075, 0.0062758237565096152, 0.0059562400705335042, 
    0.0056290544123746645, 0.0053012225711200353, 0.0049796960306249553, 
    0.0046712580114990293, 0.0043823616299901464, 0.0041189324079958494, 
    0.0038862071793365331, 0.0036885398577037464, 0.0035292424906824961, 
    0.0034104591437998958, 0.0033330783601693186, 0.0032967195598473695, 
    0.0032997937958273212, 0.0033396051600342817, 0.0034125159035173686, 
    0.0035141542699240391, 0.0036396040820846918, 0.0037836096866223049, 
    0.0039407447836003291, 0.0041055748316293208, 0.0042727880365302263, 
    0.0044373170831174952, 0.004594440308416878, 0.0047398574262657936, 
    0.0048697887533892779, 0.0049810301442671286, 0.0050710436226016446, 
    0.0051380098043675758, 0.0051808733775031476, 0.0051993317603524457, 
    0.0051938255302121502, 0.0051654457653068251, 0.0051158458109580116, 
    0.0050470957754712113, 0.0049615643513919059, 0.004861738454051405, 
    0.0047501048453105696, 0.0046290392653991295, 0.0045007615614883877, 
    0.0043673429247603965, 0.0042307514351868974, 0.004092910574782907, 
    0.0039557713425948209, 0.0038213651993433012, 0.0036918482764731319, 
    0.0035695114958058743, 0.0034567737497805144, 0.0033561590842256994, 
    0.0032702530273755154, 0.0032016054527348129, 0.003152614107463978, 
    0.0031253514188309384, 0.0031213504827472044, 0.0031413529509190432, 
    0.0031850801569741315, 0.0032509867149692999, 0.0033361158179749228, 
    0.0034360451595290046, 0.0035449318635664478, 0.0036556831294328584, 
    0.0037602018636767455, 0.0038497336580396078, 0.0039152445162613193, 
    0.0039478518369309608, 0.0039392506222545179, 0.0038821460101190501, 
    0.003770615651012272, 0.0036004411831249239, 0.0033693669553402123, 
    0.003077252786188625, 0.0027261420781256223, 0.0023202139470892783, 
    0.001865592364102799, 0.0013700807553292552, 0.00084279691654311846, 
    0.00029377652426314639, -0.00026644099489253582, -0.00082717552230192532, 
    -0.0013779268978558585, -0.001908622912284929, -0.002409802374873162, 
    -0.0028727760846056897, -0.0032897207983050873, -0.0036537778556172597, 
    -0.0039591218065924251, -0.0042010028577575895, -0.0043758111642478352, 
    -0.0044810877748211742, -0.0045155377167770058, -0.0044790168160635628, 
    -0.0043725075049120743, -0.0041980803496223951, -0.0039588620403726111, 
    -0.0036589599254009588, -0.0033033620236742026, -0.0028977898702146386, 
    -0.0024485113832757597, -0.0019621598241289367, -0.0014455493716228449, 
    -0.00090552652282169309, -0.00034882752427230012, 0.00021805826200871494, 
    0.00078899090458472087, 0.0013582646519462874, 0.0019206844312660998, 
    0.0024716155603273287, 0.003007054121066801, 0.0035237292759951735, 
    0.0040191959813557993, 0.0044919709232369032, 0.0049416082013359836, 
    0.005368734315195565, 0.0057749990761054035, 0.0061629314610721388, 
    0.0065357403090272742, 0.0068970257430732507, 0.0072505178589097469, 
    0.0075998028393854701, 0.0079480944428124041, 0.0082980833306316917, 
    0.0086518359140648048, 0.0090107210751540767, 0.0093753766160414569, 
    0.0097456780874875856, 0.010120699178707346, 0.010498664684234037, 
    0.010876919830001736, 0.011251911910373934, 0.011619211183014665, 
    0.011973594450931492, 0.012309180226980543, 0.012619635353210231, 
    0.012898423141169658, 0.013139050210145326, 0.0133353614526552, 
    0.01348176686772585, 0.013573473862147132, 0.01360667511281502, 
    0.013578692363124893, 0.013488095554316751, 0.013334763242997099, 
    0.013119873732547267, 0.012845816373572344, 0.012516008846906134, 
    0.012134675124459364, 0.0117065899924381, 0.011236785768490831, 
    0.010730330643488094, 0.010192077048609055, 0.0096264483161785947, 
    0.0090372321793982524, 0.0084274700209053827, 0.0077993329063669658, 
    0.0071541284578133246, 0.0064923556551754373, 0.005813829306019782, 
    0.0051179173211092655, 0.0044037879598085618, 0.0036707196846163886, 
    0.0029183739070515282, 0.0021470616001201259, 0.0013579043637216553, 
    0.00055296213567226265, -0.00026475022556932923, -0.0010912503279911726, 
    -0.0019216514595008789, -0.0027502230258955357, -0.0035705051882186354, 
    -0.0043754170265402903, -0.0051574425031703222, -0.0059088102164155431, 
    -0.0066217592328934585, -0.0072887776515522503, -0.0079028690743301634, 
    -0.0084578289121905337, -0.0089484503142833703, -0.0093706812304346614, 
    -0.0097217667687933759, -0.010000241893619746, -0.010205920060447838, 
    -0.010339773903874257, -0.010403803454563409, -0.010400825396583824, 
    -0.010334294396780094, -0.010208091196665889, -0.010026366867047788, 
    -0.0097933889710561627, -0.0095134266035534817, -0.0091906994337711424, 
    -0.0088293460053160688, -0.0084334225942340156, -0.0080069298496936014, 
    -0.0075538466489549413, -0.0070781399702606928, -0.006583777410670056, 
    -0.0060747027428383529, -0.0055548516510004666, -0.0050280983300093045, 
    -0.0044982760211766792, -0.003969163675425132, -0.0034444934387377097, 
    -0.0029279728633684163, -0.0024232685027670954, -0.0019339815538311328, 
    -0.0014635985583718852, -0.0010153594661664056, -0.0005921187552401252, 
    -0.00019618762085670308, 0.00017082832020737172, 0.00050811741460210437, 
    0.00081568843406123169, 0.0010942974086060003, 0.001345258184334192, 
    0.0015701960611751867, 0.0017707389449055848, 0.001948210568064775, 
    0.0021033917982434315, 0.0022363316218360764, 0.0023462655342268361, 
    0.0024316390739280271, 0.0024901897960757646, 0.0025191530530524952, 
    0.0025154870743294461, 0.0024761158349352096, 0.0023982155673221753, 
    0.0022794391467617714, 0.0021181247888774541, 0.0019134581344047356, 
    0.001665542840572212, 0.0013754457660731475, 0.0010451941290983138, 
    0.00067773722924766044, 0.00027688592302091831, -0.00015275058366438031, 
    -0.00060583441662499544, -0.0010763904144742995, -0.0015579104680914927, 
    -0.0020435241259483669, -0.0025262048900800103, -0.0029990381356408565, 
    -0.0034554904835114139, -0.0038896771211723163, -0.0042966229625236718, 
    -0.0046724440062976486, -0.0050144420335517248, -0.0053211308889406679, 
    -0.0055921865992597693, -0.0058282853739222151, -0.0060309323338682552, 
    -0.0062022029675823515, -0.0063444994188833871, -0.0064602726578564945, 
    -0.0065517921859465636, -0.0066209312690883142, -0.0066690403399634057, 
    -0.0066968240887509923, -0.0067043401171245987, -0.0066910080217725239, 
    -0.0066556204348196075, -0.0065964430557924484, -0.0065113007010339057, 
    -0.0063977684523612108, -0.0062533900455307642, -0.0060759732094150792, 
    -0.0058639667210667766, -0.0056168242128488196, -0.0053353592395303639, 
    -0.0050220794064264242, -0.0046813390871470574, -0.0043194358236993587, 
    -0.0039444896527822603, -0.0035661950317013671, -0.0031953890615844995, 
    -0.0028435190570972675, -0.0025220084354963977, -0.0022416451782140728, 
    -0.0020119751728175242, -0.0018408698292888769, -0.0017341912634780948, 
    -0.0016957651299364294, -0.0017275645141819193, -0.0018301506570400296, 
    -0.0020031916343582895, -0.0022458691090477831, -0.002557013998981067, 
    -0.0029349577403634097, -0.0033771767284685172, -0.0038799078775265958, 
    -0.0044378153237563433, -0.0050438169122602305, -0.0056890630047791643, 
    -0.0063630843227024721, -0.007054091895657635, -0.0077493550549464271, 
    -0.0084356555589369872, -0.0090997269072345521, -0.0097286733187150684, 
    -0.010310361137991697, -0.010833764888182034, -0.011289364094514717, 
    -0.011669480516844589, -0.011968543904709937, -0.012183315694859063, 
    -0.012312911908906526, -0.01235877105238037, -0.012324496356434792, 
    -0.01221558063380433, -0.012039108655582914, -0.011803441657774829, 
    -0.011517819573391536, -0.01119198949062853, -0.010835796473972533, 
    -0.010458756763410043, -0.010069611973325229, -0.0096759337099653966, 
    -0.0092837787375828901, -0.0088974658408690482, -0.0085194889988817, 
    -0.0081505492188303236, -0.0077898068590737009, -0.0074351291327078026, 
    -0.0070835655556828626, -0.0067316775635986566, -0.0063759442314650951, 
    -0.0060130349072257663, -0.0056400231495535042, -0.0052544771073780618, 
    -0.0048544995868378907, -0.0044387429608302963, -0.0040063656493616092, 
    -0.0035571089097282439, -0.0030913383931838803, -0.0026102404855901482, 
    -0.0021159550067261484, -0.0016117509145835893, -0.0011021354120251646, 
    -0.00059288629328401138, -9.1012878790459959e-05, 0.00039538402352612786, 
    0.00085740265511794194, 0.001285747051337978, 0.0016711564943571356, 
    0.0020049405820656147, 0.0022795309180170878, 0.0024889105187383131, 
    0.0026290125234970313, 0.0026979817045905061, 0.002696272181859965, 
    0.0026266299185693166, 0.0024939169110197667, 0.0023048397369999384, 
    0.0020675576861623707, 0.0017912957410382096, 0.0014858607856020199, 
    0.0011612357285865384, 0.00082712789047854158, 0.00049254073941628295, 
    0.00016539983565961355, -0.00014777918573786043, -0.00044196855663421408, 
    -0.00071360695891111488, -0.00096025728967599733, -0.001180060693764168, 
    -0.001371228223089882, -0.0015314564323905704, -0.0016575970947544393, 
    -0.0017456202722853096, -0.0017908663629566, -0.001788501486252424, 
    -0.0017341876079562343, -0.001624786112802703, -0.0014590701943747759, 
    -0.0012383266308391102, -0.00096672518134406312, -0.00065146998453680127, 
    -0.00030257230192253675, 6.7569209292513621e-05, 0.00044503246653384264, 
    0.00081519819310303426, 0.0011637829145901416, 0.001477664058385064, 
    0.0017456113814928334, 0.0019586588697185232, 0.0021103537681886075, 
    0.002196821224385961, 0.0022166574412007768, 0.0021709507061823939, 
    0.002063073705522298, 0.0018985500284197229, 0.0016847423489321314, 
    0.001430454680265196, 0.0011455445617939543, 0.00084030497213276952, 
    0.00052494276012711514, 0.00020904820661625132, -9.8753716630018383e-05, 
    -0.00039112132292740782, -0.00066215754323278603, 
    -0.00090734260851400893, -0.0011235180750976564, -0.0013087854507798716, 
    -0.0014623871801613913, -0.0015847005055129888, -0.0016772073817775206, 
    -0.0017425833690033364, -0.0017846262201628199, -0.0018077694839148646, 
    -0.0018165607790236109, -0.0018146485852957891, -0.0018037823853959659, 
    -0.0017827225143802754, -0.0017468456330510464, -0.0016879719443629064, 
    -0.0015952012143561249, -0.0014560703706836299, -0.0012583253636050395, 
    -0.00099175034880113859, -0.00064985829285142422, 
    -0.00023150132268245872, 0.0002582946686328553, 0.00080793290238373753, 
    0.0013997149365360209, 0.0020107717831059396, 0.0026148116577844778, 
    0.0031842836755485997, 0.0036926370626910671, 0.004117213579926185, 
    0.004441335531093534, 0.004655833582553023, 0.0047597729780485837, 
    0.004759943646777379, 0.0046697921952209807, 0.0045079552155162959, 
    0.0042969156903066132, 0.0040616866902773189, 0.0038287668876511157, 
    0.0036249072941104601, 0.0034753706461120104, 0.0034023465892352276, 
    0.0034232367402194401, 0.003548934523107645, 0.0037836647841262916, 
    0.0041243797047809047, 0.0045623027389385517, 0.0050825937798804951, 
    0.005667028425276755, 0.0062940844269204991,
  // Fqt-Na(6, 0-1999)
    1, 0.99525514200276555, 0.98118345865806333, 0.95826197249951617, 
    0.92725015280821366, 0.88914136643478581, 0.84510217195588988, 
    0.79640533442726058, 0.7443624430501119, 0.69026140116349077, 
    0.63531290417668107, 0.58060855147365653, 0.52709180469108974, 
    0.47554167684725823, 0.42656795033076378, 0.38061607008016901, 
    0.33797942376950707, 0.29881669941117411, 0.26317208751700505, 
    0.23099651924544262, 0.20216840491364976, 0.17651284361453751, 
    0.15381861301812955, 0.13385258810941031, 0.11637153789108087, 
    0.1011313757662415, 0.087894119975661697, 0.076432853935906944, 
    0.066535017818098952, 0.058004367235986273, 0.050661901130126211, 
    0.044346024548025186, 0.038912186978035244, 0.034232152845768936, 
    0.030193052678729817, 0.026696302510363788, 0.023656464258557258, 
    0.021000097268087891, 0.018664619638260351, 0.016597219535317863, 
    0.014753793918420891, 0.013097950037149123, 0.011600028341108423, 
    0.010236181120547042, 0.0089874812713434584, 0.0078390704433615819, 
    0.0067793637161826948, 0.0057993051296101848, 0.0048917076472989778, 
    0.004050669433042847, 0.0032711028009851594, 0.0025483735755924843, 
    0.0018780519384820889, 0.0012557833028370446, 0.00067725591915545995, 
    0.00013824576149541241, -0.00036527460204755901, -0.00083700034587513102, 
    -0.0012801601614883167, -0.0016973922751314515, -0.0020906687259973134, 
    -0.0024612656174989147, -0.0028097862523695401, -0.0031362252606148533, 
    -0.0034400724442465191, -0.0037204177941450958, -0.0039760889717422674, 
    -0.0042057754423930156, -0.004408194169637219, -0.0045822615301920316, 
    -0.0047272787773026299, -0.0048430935112285575, -0.0049302192103070986, 
    -0.0049898711375860961, -0.0050239116879113943, -0.0050347217964491278, 
    -0.0050249930025340088, -0.004997492633095334, -0.0049548225654002442, 
    -0.004899207637744098, -0.0048323422387746284, -0.0047553156649760269, 
    -0.0046686164149376966, -0.004572219069641662, -0.0044657342696331863, 
    -0.004348603016201969, -0.0042203063393001349, -0.0040805696065497471, 
    -0.0039295401698712356, -0.0037679209629917091, -0.0035970459124058537, 
    -0.0034189006685147851, -0.0032360920957028713, -0.003051767152280315, 
    -0.0028694999523468075, -0.0026931359634355259, -0.0025266171388279336, 
    -0.0023737869535100137, -0.0022382063358321754, -0.0021229778275645233, 
    -0.0020305999872787606, -0.0019628700041209269, -0.0019208150244079472, 
    -0.0019046680695001834, -0.0019138738971227805, -0.0019471143461838288, 
    -0.0020023596671055917, -0.0020769203865764999, -0.0021675140878508188, 
    -0.0022703328358441416, -0.002381121027117222, -0.0024952669818029492, 
    -0.0026079067448042084, -0.0027140675596133714, -0.0028088230809589026, 
    -0.0028874958652835695, -0.0029458661254801043, -0.0029804004438136154, 
    -0.0029884518402980126, -0.0029684236591668292, -0.0029198678080791921, 
    -0.002843504110243636, -0.0027411614886325127, -0.0026156422430639653, 
    -0.0024705178027259315, -0.00230987369070968, -0.0021380141126543426, 
    -0.0019591646766754811, -0.0017771973837995155, -0.0015954095377886622, 
    -0.0014163832507710665, -0.0012419357650883815, -0.0010731532162010339, 
    -0.0009104889993652121, -0.00075389929838398477, -0.00060300868604365974, 
    -0.00045725884263097345, -0.00031603831484728587, 
    -0.00017879349437473679, -4.5094980193350503e-05, 8.5316581585928933e-05, 
    0.00021251311421656774, 0.00033637484337497876, 0.00045659939465145271, 
    0.00057271387772098235, 0.00068409403482521118, 0.00078999406087561252, 
    0.00088957469392184616, 0.00098194708099300196, 0.0010662134732907004, 
    0.0011415065414647316, 0.0012070138550423926, 0.0012619894321030444, 
    0.0013057441604447492, 0.0013376388849169591, 0.0013570687679244782, 
    0.0013634772852469728, 0.0013563778356957133, 0.0013353889868197748, 
    0.0013002599735492627, 0.0012508929913670199, 0.0011873335289457332, 
    0.0011097577945739332, 0.0010184408007302872, 0.00091374378907783287, 
    0.00079611039793178772, 0.00066609757163861951, 0.00052440560051251095, 
    0.00037193890158424139, 0.00020983917832651054, 3.952840337644047e-05, 
    -0.00013726988070252288, -0.00031853152080500539, 
    -0.00050194885735687039, -0.00068499022668811436, 
    -0.00086498715578519443, -0.0010392453555654294, -0.001205172714316316, 
    -0.0013604067666248413, -0.0015029195007473643, -0.0016311163171724239, 
    -0.0017438872287825896, -0.0018406470025634611, -0.0019213330552795007, 
    -0.001986390011865723, -0.002036715201969427, -0.002073592628651779, 
    -0.0020986154188945109, -0.0021135969243157087, -0.0021204812717672988, 
    -0.0021212636481066651, -0.002117913860805727, -0.002112298668310854, 
    -0.002106124382583919, -0.0021008700427885929, -0.0020977418309703947, 
    -0.0020976348079409825, -0.002101094971214113, -0.0021083045336922394, 
    -0.0021190610130823063, -0.0021327663896326234, -0.0021484242629405304, 
    -0.0021646509698647468, -0.0021797029105996586, -0.0021915283149565317, 
    -0.0021978373348341294, -0.0021961904674384631, -0.0021841058258672743, 
    -0.0021591679766756553, -0.0021191364983205573, -0.0020620420525054662, 
    -0.0019862645594348736, -0.0018905786334708422, -0.0017741832845940522, 
    -0.0016366968665413714, -0.0014781331509384306, -0.001298862755328491, 
    -0.0010995641619749308, -0.00088118565492987882, -0.00064491300269313347, 
    -0.00039215490860222148, -0.00012456055701879173, 0.00015595145953740654, 
    0.00044714431957000128, 0.00074640338610733521, 0.0010506866659800627, 
    0.0013564841883282829, 0.0016598060570771891, 0.0019561937528546815, 
    0.0022407819748132803, 0.0025083974825475365, 0.0027537004086735342, 
    0.0029713605075218437, 0.0031562619420643437, 0.0033037112587304984, 
    0.0034096496728671238, 0.0034708426218899883, 0.0034850478253767802, 
    0.0034511433752594748, 0.0033692141965297904, 0.0032405861205618467, 
    0.0030678066362178347, 0.0028545604468012443, 0.0026055321155312597, 
    0.0023262115737032246, 0.0020226639605782793, 0.0017012755138863407, 
    0.0013684918271734499, 0.0010305754134686206, 0.00069339387108995065, 
    0.00036224924363247556, 4.1758617439069412e-05, -0.00026422395324417273, 
    -0.00055264464792290405, -0.0008212601681583478, -0.0010686299708113317, 
    -0.0012940975659128039, -0.0014977600253547041, -0.0016804239925417856, 
    -0.001843537569598459, -0.0019891137489312337, -0.0021196308404406012, 
    -0.0022379180729640942, -0.0023470431190093489, -0.0024501815618544467, 
    -0.0025504724814898556, -0.0026508597653996774, -0.0027539117975453479, 
    -0.0028616405862830489, -0.00297532689366824, -0.0030953984641701564, 
    -0.0032213453625931951, -0.0033517337259487251, -0.0034842807566660152, 
    -0.0036160188302186039, -0.0037435038114565383, -0.0038630738256736773, 
    -0.0039711165246550904, -0.0040643365861967465, -0.0041399789223838532, 
    -0.0041960204486071401, -0.0042312851424789744, -0.004245485605543344, 
    -0.0042391808425117352, -0.0042136593651990722, -0.0041707490300726307, 
    -0.0041125732516349104, -0.0040412754995986519, -0.0039587474755586822, 
    -0.0038663779734697604, -0.0037648674557598173, -0.0036541389002305983, 
    -0.0035333517048436935, -0.0034010353824737941, -0.0032553280449071137, 
    -0.0030942886647750728, -0.0029162566400536085, -0.0027201998903269133, 
    -0.0025060361831789808, -0.002274867238199202, -0.0020291132679275863, 
    -0.0017725332022651124, -0.0015101364501581196, -0.0012479889880849925, 
    -0.00099292578448222199, -0.00075221193882164729, 
    -0.00053317249336235937, -0.00034281325845869425, 
    -0.00018746833692542418, -7.2504296692798417e-05, 
    -2.0839421347213665e-06, 2.0977358447929554e-05, -4.7308506482243083e-06, 
    -7.9252782457747608e-05, -0.00020136867997714143, 
    -0.00036875265979088281, -0.00057815126616617715, -0.0008255460879075568, 
    -0.0011062868490279106, -0.0014151813941603315, -0.0017465384645122687, 
    -0.0020941985832825176, -0.0024515565589622178, -0.0028116256430947644, 
    -0.003167134725644033, -0.0035106887931696923, -0.0038349651696188364, 
    -0.0041329450962344265, -0.0043981514486491884, -0.0046248749950874267, 
    -0.0048083788510710733, -0.0049450595608035632, -0.0050325608737775678, 
    -0.0050698388430258194, -0.0050571725457223384, -0.0049961236092292381, 
    -0.0048894453801964612, -0.0047409496589776983, -0.0045553329796284093, 
    -0.0043379692783964072, -0.0040946733531729285, -0.0038314480557243773, 
    -0.0035542292511356851, -0.0032686426664795903, -0.0029797801076815451, 
    -0.0026920228621487288, -0.002408913516801451, -0.0021330814855405147, 
    -0.0018662466740216848, -0.0016092944781810404, -0.001362415617308802, 
    -0.0011253004167467268, -0.00089735242700246412, -0.00067789978725670474, 
    -0.00046638168274213744, -0.00026248999036595111, 
    -6.6255434355477999e-05, 0.00012194013177112067, 0.00030141773243589872, 
    0.00047130086983229768, 0.00063065492560966804, 0.0007786412110434716, 
    0.00091465993379144755, 0.0010384676890654574, 0.0011502572414686147, 
    0.0012506867335697865, 0.0013408507632924143, 0.0014222109288605969, 
    0.0014964799778853753, 0.0015654914070147327, 0.0016310641466306154, 
    0.0016948887237429478, 0.0017584373595049046, 0.0018229186952089774, 
    0.0018892530279930992, 0.0019580852032344475, 0.002029799115333374, 
    0.0021045450749648362, 0.0021822610914017655, 0.0022626803800026738, 
    0.0023453339648249875, 0.0024295351381050695, 0.0025143535319817564, 
    0.0025985881896539087, 0.0026807444962069953, 0.0027590209788906288, 
    0.002831325096906619, 0.002895309657841392, 0.0029484573905279362, 
    0.0029882006550312396, 0.0030120863655437686, 0.003017967020260207, 
    0.0030042176030312898, 0.0029699333987408616, 0.0029151042314264435, 
    0.0028407412633741675, 0.002748943512337656, 0.0026428918883501171, 
    0.0025267609451341032, 0.0024055542064730568, 0.0022848570545602517, 
    0.0021705221763446136, 0.0020683186306947408, 0.0019835559859609406, 
    0.0019207315230016487, 0.001883214624804482, 0.0018730090783725341, 
    0.0018906098369593973, 0.0019349682254226051, 0.0020035552492360712, 
    0.0020925392754979023, 0.0021970313034427699, 0.0023113959884101215, 
    0.0024295955691576452, 0.0025455488695534374, 0.0026534815589830266, 
    0.0027482476010868562, 0.0028256056368798094, 0.0028824285720588459, 
    0.0029168400079266012, 0.002928260748222067, 0.0029173613959619462, 
    0.0028859288345530034, 0.0028366475523002653, 0.0027728319220425529, 
    0.002698138985931413, 0.0026162926696284092, 0.0025308453866967409, 
    0.0024449902188976957, 0.0023614298664649197, 0.0022822962909226346, 
    0.0022091244622332879, 0.0021428657172495287, 0.0020839432340424156, 
    0.0020323401641024019, 0.0019877113188216467, 0.0019495100007589929, 
    0.0019171253102690912, 0.0018900080538213509, 0.0018677822145246313, 
    0.0018503185520504085, 0.0018377522137050383, 0.0018304521864494334, 
    0.0018289285896556811, 0.0018337052769499056, 0.0018451725011684348, 
    0.0018634352450159941, 0.0018881880213470915, 0.0019186187109734316, 
    0.0019533654649666627, 0.0019905112421277692, 0.0020276486744120244, 
    0.0020619860406284741, 0.0020904943606525851, 0.0021100721311695515, 
    0.0021176989494074965, 0.0021105606031028177, 0.0020861385624622564, 
    0.0020422787866443818, 0.0019772407917493157, 0.0018897414632088703, 
    0.0017789881613400641, 0.0016447125553671399, 0.0014871872603457851, 
    0.0013072330880046926, 0.001106214256244498, 0.00088602445565408923, 
    0.00064906474260343532, 0.00039822325494076724, 0.00013684558885941299, 
    -0.00013130686747637383, -0.00040211506807504461, 
    -0.00067118237616117088, -0.00093394142221513393, -0.0011857700134366, 
    -0.0014221281255121893, -0.001638692178209968, -0.0018314909336971873, 
    -0.0019970333773729333, -0.002132409871399326, -0.0022353831524921505, 
    -0.0023044464705444336, -0.0023388553944966198, -0.0023386358863642723, 
    -0.0023045619513563107, -0.0022381142543922623, -0.0021414165056683936, 
    -0.0020171564272543669, -0.0018684924085573061, -0.0016989449980318932, 
    -0.0015122859952057259, -0.0013124210071953088, -0.0011032773967476323, 
    -0.00088870007471279571, -0.00067235136243782494, 
    -0.00045761045894544264, -0.00024748751611895466, 
    -4.4520916082570438e-05, 0.00014930657011358886, 0.0003326378947416756, 
    0.00050478001704088913, 0.00066569619270729133, 0.00081595928455933226, 
    0.00095666168116359648, 0.0010892852976834443, 0.0012155481516049566, 
    0.0013372194555061516, 0.0014559371748167739, 0.001573034426575358, 
    0.0016893926810466202, 0.0018053285594402291, 0.0019205240415401895, 
    0.0020340082717123205, 0.002144171987344139, 0.0022488418324549827, 
    0.0023453842019216945, 0.0024308487831523622, 0.0025021405412334074, 
    0.0025562085624950088, 0.0025902463366062585, 0.0026018797822683756, 
    0.0025893402823166886, 0.0025515923477920678, 0.0024884276866359275, 
    0.0024004959496874557, 0.0022892837818526924, 0.0021570430867096377, 
    0.0020066653982362768, 0.0018415279750524137, 0.001665309737831122, 
    0.001481814866093706, 0.0012947961773317885, 0.001107801266762478, 
    0.00092402769099876375, 0.00074620443814865244, 0.0005764891642841424, 
    0.00041640640662325175, 0.0002668208798100812, 0.00012794819683026483, 
    -6.0720365213954783e-07, -0.00011979637881211175, 
    -0.00023105506681937759, -0.00033623532691131469, -0.0004375320215049819, 
    -0.00053739599432098782, -0.00063843737157919119, 
    -0.00074331731398395696, -0.0008546228592239861, -0.0009747314620308803, 
    -0.0011056708287177474, -0.0012489780145076585, -0.0014055612094059301, 
    -0.001575585119001404, -0.0017583716934367769, -0.0019523431625036922, 
    -0.0021550026116727351, -0.0023629587881027823, -0.0025719943770103186, 
    -0.0027771762491395069, -0.0029730092691264598, -0.0031536331482475612, 
    -0.0033130616201593214, -0.0034454498761813785, -0.0035453759984555269, 
    -0.0036081224297562506, -0.0036299344971605263, -0.0036082405231533336, 
    -0.0035418134443378621, -0.0034308543661956932, -0.003277009420981687, 
    -0.0030832998575778684, -0.0028539840058282367, -0.0025943505900991089, 
    -0.0023104693543268013, -0.0020089103823673861, -0.0016964572523290387, 
    -0.0013798273931557455, -0.0010654255711470919, -0.00075913439110924076, 
    -0.00046615609108113028, -0.00019090143312079622, 6.3073575387342885e-05, 
    0.00029309433368327771, 0.00049735780585786278, 0.00067491166190327019, 
    0.00082560666082261299, 0.00095003926174133245, 0.0010494842060706448, 
    0.0011258006323970494, 0.0011813303319528508, 0.0012187763135525595, 
    0.0012410705569459726, 0.0012512353476010494, 0.0012522530835809328, 
    0.0012469314701628346, 0.0012377872330318639, 0.0012269265120080474, 
    0.0012159453322982546, 0.0012058401614535338, 0.0011969388173859346, 
    0.0011888798087342231, 0.0011806255607963263, 0.0011705455583138373, 
    0.0011565419426552536, 0.0011362307890308997, 0.0011071359666178578, 
    0.0010668819836264531, 0.0010133620467537097, 0.00094485227881566385, 
    0.00086008799691550441, 0.00075827821877320423, 0.0006390824845885169, 
    0.00050257700349863002, 0.00034920523541846001, 0.00017973993010636643, 
    -4.7445612322889893e-06, -0.00020288951320093389, 
    -0.00041306325242294059, -0.00063336960613333726, 
    -0.00086165290929613044, -0.001095504828806848, -0.0013322646510562602, 
    -0.0015690291068614082, -0.0018026611373528015, -0.0020298173144195596, 
    -0.0022469967161750024, -0.0024506338032745222, -0.0026372230778203623, 
    -0.0028034905651892657, -0.0029465804164792082, -0.0030642243864460565, 
    -0.0031548840120799917, -0.0032178208446196101, -0.0032531165563079909, 
    -0.0032616206753481318, -0.0032448573596407966, -0.0032048867634089551, 
    -0.0031441504638345598, -0.0030653030765760317, -0.0029710447952856476, 
    -0.0028639719838103057, -0.0027464513682457208, -0.0026205301470347822, 
    -0.0024878885722066034, -0.0023498338659950551, -0.0022073306000605086, 
    -0.0020610546953433034, -0.0019114698011450425, -0.0017589164007698486, 
    -0.0016036930065995883, -0.0014461320206458942, -0.0012866682596110455, 
    -0.0011258906417793875, -0.00096458042855496727, -0.00080373953939328875, 
    -0.0006446121646529893, -0.00048869067933201985, -0.00033771944660041648, 
    -0.00019367907442765343, -5.8763484857845638e-05, 6.4674316807062813e-05, 
    0.00017418422761462764, 0.00026730328816675482, 0.00034165077808086459, 
    0.00039502792262747724, 0.00042552531104546939, 0.00043163342604563823, 
    0.00041234801645450669, 0.00036726501788503067, 0.00029665681602899992, 
    0.00020152569531222298, 8.3621771933121839e-05, -5.456995711098343e-05, 
    -0.00020988641893361431, -0.00037856717964434748, 
    -0.00055637881489317871, -0.00073877764399182008, 
    -0.00092110313856404299, -0.001098794865065857, -0.0012676169106558023, 
    -0.0014238866335328803, -0.0015646756981759096, -0.0016879824309496763, 
    -0.0017928355855117094, -0.0018793449825043032, -0.0019486744521149549, 
    -0.0020029504749355725, -0.0020451172065954035, -0.002078727440848996, 
    -0.0021077119536126185, -0.0021361223506919523, -0.0021678667085239171, 
    -0.0022064755699308936, -0.0022549005812316212, -0.0023153746617450141, 
    -0.0023893310576479742, -0.0024774007012912319, -0.0025794484037644167, 
    -0.002694662126784441, -0.0028216530058233886, -0.0029585439491574108, 
    -0.0031030556048075777, -0.0032525659427958663, -0.0034041576587912521, 
    -0.0035546653276423016, -0.0037007243401089864, -0.003838837288708436, 
    -0.0039654675778961366, -0.0040771698680240063, -0.0041707508677752215, 
    -0.0042434578338936043, -0.0042931602786498747, -0.0043185206495599451, 
    -0.0043191121010887849, -0.0042954668518566247, -0.0042490515698172457, 
    -0.004182160358687334, -0.0040977382969607954, -0.0039991626280247265, 
    -0.0038899975937587137, -0.003773756804371876, -0.0036536860737920525, 
    -0.0035325996555631389, -0.0034127685311433681, -0.0032958783519657598, 
    -0.0031830505896940182, -0.0030749164782707524, -0.0029717278716488334, 
    -0.00287349200309124, -0.0027801114139045964, -0.0026915166351117762, 
    -0.0026077840995586349, -0.0025292337535838109, -0.0024564934650265764, 
    -0.0023905215036126724, -0.0023325713577562082, -0.0022841055858034785, 
    -0.0022466537125358397, -0.0022216336653380748, -0.0022101695893067402, 
    -0.0022129215731169845, -0.0022299532537126687, -0.0022606401937387429, 
    -0.0023036310056101569, -0.0023568485572653141, -0.0024175320275540845, 
    -0.0024823164660352894, -0.0025473361672253107, -0.0026083419978114391, 
    -0.0026608460321578663, -0.0027002797374433502, -0.0027221714066791632, 
    -0.0027223562549147529, -0.0026971837519174794, -0.0026437398476974027, 
    -0.0025600552655840937, -0.0024452913831084916, -0.0022998860045201938, 
    -0.0021256433173030141, -0.0019257473933832242, -0.0017046970694275291, 
    -0.0014681481682569948, -0.0012226746827864283, -0.00097545389294659518, 
    -0.00073388555345773807, -0.00050518747199071652, 
    -0.00029598204443314941, -0.00011191888178685848, 4.2627940455501557e-05, 
    0.0001647830869895114, 0.00025326340703661111, 0.00030836107270509639, 
    0.00033181015491699637, 0.00032655521255497223, 0.00029645739947487589, 
    0.00024596736982333508, 0.00017979063739953131, 0.00010257881413601889, 
    1.8658963359535654e-05, -6.8176109176251568e-05, -0.00015481964837136912, 
    -0.00023893299981666974, -0.00031895393850500219, 
    -0.00039404202650757353, -0.00046396451048869394, 
    -0.00052893674457910869, -0.0005894343812116186, -0.00064599127854791569, 
    -0.00069901802066621368, -0.0007486296842871583, -0.00079453780961439842, 
    -0.0008359718689473774, -0.00087166405808127142, -0.00089989625135113204, 
    -0.00091859220751403154, -0.00092546782762818237, 
    -0.00091820938847967856, -0.00089468115360289476, 
    -0.00085313605087510968, -0.00079241042668550497, 
    -0.00071209442306366714, -0.00061265032508486339, 
    -0.00049548665840700801, -0.00036296070637889842, 
    -0.00021833607356072204, -6.5671252537983691e-05, 9.0335455502542133e-05, 
    0.00024452691391129398, 0.000391499931319426, 0.00052581485923275959, 
    0.00064220830575287507, 0.00073579418090686318, 0.00080225819069957823, 
    0.00083804556677931049, 0.00084053319408696641, 0.00080817373189338935, 
    0.0007406103353541861, 0.00063872906363855318, 0.00050465074911583614, 
    0.00034165848344211045, 0.00015406092622840487, -5.3004126545421327e-05, 
    -0.00027380444730638269, -0.00050227747575409343, 
    -0.00073229191257871337, -0.00095789713528777619, -0.0011735400331955932, 
    -0.0013742315647535933, -0.0015556635349105847, -0.0017142738227955766, 
    -0.0018472615461435108, -0.0019525632305943709, -0.0020287926297197592, 
    -0.0020751720810297664, -0.0020914465067648088, -0.0020778096331041285, 
    -0.0020348318118132004, -0.0019634127604763905, -0.0018647406382275315, 
    -0.0017402680885212868, -0.0015916940796970674, -0.001420957616909654, 
    -0.001230228254744458, -0.001021904983085293, -0.00079860890649886514, 
    -0.0005631797368853852, -0.00031866397939084361, -6.8321874069423704e-05, 
    0.00018437397992580065, 0.00043573548005821977, 0.00068184400691606161, 
    0.00091855597375570296, 0.001141525605501311, 0.0013462601718059104, 
    0.0015282241545757386, 0.0016829878891205954, 0.0018064203034444228, 
    0.001894899476124535, 0.0019455334644210187, 0.0019563451846607875, 
    0.0019264272181987703, 0.0018560242717094405, 0.0017465509154917223, 
    0.0016005318701455442, 0.0014214796707640647, 0.0012136979145170009, 
    0.00098204041565889836, 0.00073164512031958834, 0.00046765873478889707, 
    0.00019498619952820865, -8.1903465917855436e-05, -0.00035910079532350963, 
    -0.00063330674165143659, -0.00090180167582648357, -0.0011623723181466913, 
    -0.0014132255123412954, -0.0016528907540441253, -0.0018801628194976879, 
    -0.0020940603317095648, -0.0022938097511600143, -0.0024788402313832419, 
    -0.0026487772226615486, -0.0028034294246840853, -0.0029427549619729307, 
    -0.0030668126354522246, -0.0031757146104596087, -0.0032695650613488014, 
    -0.0033484066522053257, -0.0034121591776030366, -0.0034605651628952256, 
    -0.0034931368901209604, -0.0035091130882857085, -0.0035074360005208022, 
    -0.0034867625273156165, -0.0034455132641370042, -0.0033819675681301658, 
    -0.0032943907062958381, -0.0031812047988097917, -0.0030411662036264582, 
    -0.0028735439111904695, -0.0026782823860980205, -0.0024561199388020288, 
    -0.0022086778360901915, -0.0019384843726372499, -0.0016489627367282937, 
    -0.0013443721957129033, -0.0010297051703304059, -0.00071055380496628129, 
    -0.00039292006132494257, -8.3010731081168375e-05, 0.00021303962361288132, 
    0.00048945727216930229, 0.00074113245367440743, 0.0009638978251411322, 
    0.0011547348227542932, 0.0013119097165354779, 0.0014350252674392762, 
    0.0015249977817322282, 0.0015839801585100194, 0.0016152324901633592, 
    0.0016229571662828457, 0.0016121093992163716, 0.0015881824401282997, 
    0.0015570000144460795, 0.0015245095885499046, 0.001496589814318539, 
    0.0014788726439327812, 0.0014765886633742128, 0.0014944177062867817, 
    0.0015363510041557712, 0.001605557275769717, 0.0017042596285724784, 
    0.0018336187809330556, 0.0019936319965149349, 0.0021830737872539788, 
    0.0023994618781823405, 0.0026391081538815787, 0.0028972181039896563, 
    0.003168067379209953, 0.003445233054223484, 0.0037218628674991917, 
    0.0039909534116734247, 0.0042456109867204956, 0.0044792815187209949, 
    0.0046859410249428185, 0.0048602500708937579, 0.0049976838980706033, 
    0.0050946395826454282, 0.0051485390169001381, 0.0051578962006483594, 
    0.0051223680018815188, 0.0050427659885025795, 0.004921013924785088, 
    0.0047600549395237605, 0.0045637024928452006, 0.0043364321126103996, 
    0.0040831467380705007, 0.003808920013371981, 0.0035187423946840104, 
    0.0032172967698869521, 0.0029087714908545806, 0.0025967334032191568, 
    0.0022840532320553054, 0.0019728991170580613, 0.0016647623404722088, 
    0.0013605471617694925, 0.001060676772029297, 0.00076522271768521342, 
    0.0004740449555957538, 0.00018692567544164985, -9.6297725775980943e-05, 
    -0.00037561114676962058, -0.00065070787157323724, 
    -0.00092088886341741148, -0.0011849747911203122, -0.0014412369121630472, 
    -0.0016873655603794797, -0.0019204725066114831, -0.0021371612067464089, 
    -0.0023336500233823547, -0.0025059699848943916, -0.0026502097524556279, 
    -0.0027628129565908295, -0.0028408744441951145, -0.0028824331698066117, 
    -0.0028867387810693123, -0.0028544458841455508, -0.0027877521505179238, 
    -0.0026904301883170691, -0.0025677630124382191, -0.002426370859026996, 
    -0.0022739215774135449, -0.0021187493108381535, -0.0019693807992089002, 
    -0.0018340038047049375, -0.0017199094739771294, -0.001632970264362754, 
    -0.0015771754074887965, -0.0015543156620114935, -0.001563809469085286, 
    -0.0016027293204448536, -0.0016660048202068963, -0.0017468096377569371, 
    -0.0018370795234335584, -0.0019281339488062068, -0.0020113170137457856, 
    -0.0020786066376711427, -0.0021231351397658503, -0.0021395579457121469, 
    -0.0021242630036767841, -0.002075427328748821, -0.0019929384031098503, 
    -0.0018782520410529878, -0.0017342065727255092, -0.0015648119421250936, 
    -0.0013750248474606267, -0.001170501475588541, -0.00095733096616054062, 
    -0.00074174968968968686, -0.00052985176240586047, 
    -0.00032731908806763182, -0.00013918866754303067, 3.0341219453744781e-05, 
    0.00017803754956295751, 0.00030171348100134412, 0.00040025995077180924, 
    0.00047363531426500923, 0.00052282154878352527, 0.00054972124311857234, 
    0.00055702267787842105, 0.00054801512682348846, 0.00052636621221691842, 
    0.00049586988219907759, 0.0004602007055273295, 0.00042267812238421573, 
    0.00038608056519551519, 0.00035250985919578221, 0.00032334034055776111, 
    0.00029923135700627741, 0.00028021343012459037, 0.00026583225693214036, 
    0.00025532871330178822, 0.00024783649892239914, 0.00024258344426618367, 
    0.00023905730036130726, 0.00023712235261424242, 0.00023706441340935936, 
    0.00023955988672952415, 0.0002455596119316216, 0.00025611712282787844, 
    0.00027219696067884116, 0.00029448400390353339, 0.00032322088825143187, 
    0.00035810404704111117, 0.00039821981179715587, 0.00044204219794704701, 
    0.00048746285770877112, 0.00053186405338719197, 0.0005722239100639469, 
    0.00060524321953575534, 0.00062750001333823906, 0.00063561319236626738, 
    0.00062642361851292727, 0.00059716613734992949, 0.00054563642763726041, 
    0.00047032197716146042, 0.00037051331743386603, 0.00024636058867825029, 
    9.8901801082045188e-05, -6.9944338369003342e-05, -0.00025740429460361568, 
    -0.00045990002478184618, -0.00067312011971442059, 
    -0.00089211635036258929, -0.001111436770950085, -0.0013253092102689379, 
    -0.0015278742525668934, -0.0017134641224060426, -0.0018769232433417256, 
    -0.0020139306078071828, -0.0021213028843683392, -0.0021972333109544959, 
    -0.0022414250925433875, -0.0022550949459774782, -0.0022408547194710982, 
    -0.0022024561284173733, -0.0021444495048658172, -0.0020717818777152681, 
    -0.0019893737536329781, -0.0019017231326594274, -0.0018125696714698448, 
    -0.0017246560700184535, -0.0016395924897733749, -0.0015578355066845221, 
    -0.0014787612633360345, -0.00140082350095355, -0.0013217651654263353, 
    -0.0012388725123265152, -0.0011492295730193369, -0.0010499802177189052, 
    -0.00093854202983985596, -0.00081278952901740103, 
    -0.00067119575264256272, -0.00051291164738308801, 
    -0.00033778620808312855, -0.00014633276103817811, 6.0366755623077358e-05, 
    0.00028079447493341801, 0.00051314707217577343, 0.00075548938003994703, 
    0.0010058920376287274, 0.0012625345359034523, 0.0015237732107888601, 
    0.0017881804841081146, 0.0020545462692047006, 0.0023218393111126591, 
    0.002589158241959575, 0.0028556500950603272, 0.0031203958227945298, 
    0.003382299233721334, 0.0036399473990260558, 0.0038915016979936064, 
    0.0041346279954883403, 0.0043664713155122927, 0.0045837206934931599, 
    0.0047827216069997918, 0.0049596749950718503, 0.0051108480604423476, 
    0.0052328175680807316, 0.0053226923114946994, 0.0053782953562267529, 
    0.0053982921757838214, 0.0053822684868385408, 0.0053307320986569397, 
    0.0052450742457141909, 0.00512749801246063, 0.004980923261881892, 
    0.0048088806947652702, 0.0046154085488785508, 0.0044049448938537402, 
    0.0041822099510959374, 0.0039520781865067973, 0.0037194374271591309, 
    0.0034890293879177941, 0.0032652877160096209, 0.0030521784862760364, 
    0.0028530613240596234, 0.0026705823732579496, 0.0025066155637179159, 
    0.0023622499084892212, 0.0022378429628182616, 0.0021331149824073106, 
    0.0020473058368686158, 0.0019793504866817318, 0.0019280890946942425, 
    0.0018924398395735926, 0.0018715513371351665, 0.0018648839490204934, 
    0.0018722126383386517, 0.0018935674019786453, 0.0019290911651303473, 
    0.0019788836923427745, 0.0020428171168801507, 0.0021203888811453988, 
    0.0022106086021974895, 0.0023119546731421472, 0.0024223933147830105, 
    0.0025394706633502431, 0.002660447045517161, 0.0027824678340958617, 
    0.002902755319895688, 0.0030187732494565771, 0.0031283798257372652, 
    0.0032299281286309492, 0.0033223240659222783, 0.0034050088574837331, 
    0.0034779091206860939, 0.0035413182209750034, 0.0035957346430317222, 
    0.0036416708304882351, 0.0036794373282580312, 0.0037089461738666171, 
    0.0037295541974540726, 0.0037399802480282502, 0.0037383000826748426, 
    0.0037220521652930588, 0.0036884038795822341, 0.0036343960588831568, 
    0.0035572032124296131, 0.0034544120620631216, 0.0033242643188554593, 
    0.0031658437481559844, 0.002979212316443638, 0.0027654555458560097, 
    0.0025266464431149818, 0.0022657533936698464, 0.0019864729308468518, 
    0.0016930331297800899, 0.0013899536512626059, 0.0010818167232349025, 
    0.00077303299427420593, 0.00046762463237017048, 0.00016903573681185317, 
    -0.00012002381809569072, -0.00039767839221179326, 
    -0.00066292512824550707, -0.00091560616031843172, -0.0011563197300707819, 
    -0.0013862741340446765, -0.0016071062677411444, -0.0018206804431109504, 
    -0.0020288715188062061, -0.0022333656917249947, -0.0024354656568208017, 
    -0.0026359230835435931, -0.0028347935665074008, -0.003031316939372052, 
    -0.003223849812415375, -0.0034098280613025752, -0.0035858086021482143, 
    -0.0037475713419317675, -0.0038903036936960237, -0.0040088536327589058, 
    -0.0040980231674671063, -0.0041529052146065939, -0.0041692005460968835, 
    -0.0041435044932783497, -0.0040735381337261289, -0.0039582835751450184, 
    -0.003798057488486108, -0.0035945071621000481, -0.0033505407442234424, 
    -0.0030702306060470205, -0.0027586732511196469, -0.0024218365026417396, 
    -0.0020663805460404876, -0.0016994818481225141, -0.0013286420958550714, 
    -0.00096149834221392438, -0.00060565974424400218, 
    -0.00026852344813797909, 4.2884286532753475e-05, 0.00032208858433512558, 
    0.00056332598273149833, 0.00076171546352535107, 0.00091341238683124765, 
    0.0010157490433668696, 0.0010673429663046058, 0.0010681661129358065, 
    0.0010195954266865458, 0.00092440731219175934, 0.00078673068507566072, 
    0.00061194178120960716, 0.00040648302775514076, 0.00017764707606061003, 
    -6.6707947462882669e-05, -0.00031846742849635999, 
    -0.00056959580360310051, -0.00081247613419296828, -0.0010402264046604857, 
    -0.0012469679778038601, -0.0014280298991645899, -0.0015800296447831834, 
    -0.0017008872432271544, -0.0017897287569143053, -0.0018467276145815424, 
    -0.0018729144830622246, -0.001869959073384159, -0.0018399805931240646, 
    -0.0017853673685560337, -0.0017086241253099009, -0.0016122364452502832, 
    -0.0014985754585444223, -0.0013698286345434822, -0.0012279721730916477, 
    -0.0010747968632730317, -0.00091196749176348537, -0.00074111780713103292, 
    -0.00056393821048156484, -0.00038224549206072064, 
    -0.00019801398655918995, -1.3371755467182984e-05, 0.00016945876376697923, 
    0.00034823453490278006, 0.00052080493371930319, 0.00068522699124992398, 
    0.00083988514665876127, 0.00098359156155572642, 0.0011156363609344379, 
    0.0012358006191747761, 0.0013443186473147829, 0.0014417796429657377, 
    0.0015289958875155756, 0.0016068446065063424, 0.0016761100380254372, 
    0.0017373445584636608, 0.0017907721567007255, 0.001836210072573377, 
    0.0018730571961886495, 0.0019003016555195216, 0.0019165526303894483, 
    0.0019201113762133859, 0.0019090470232983455, 0.001881307729094571, 
    0.0018348508931214013, 0.0017677919926624599, 0.0016785514574853074, 
    0.0015659965239838015, 0.0014295347090553276, 0.0012692003419687119, 
    0.0010856786888204604, 0.00088032931210680915, 0.00065516242679348709, 
    0.00041277876271737215, 0.0001562503595759823, -0.00011104598832277978, 
    -0.00038562644891119828, -0.00066410503824485933, 
    -0.00094337371132915059, -0.0012206876249222802, -0.0014936979839211355, 
    -0.0017604003365429906, -0.0020190564200795948, -0.0022681257333040973, 
    -0.0025062385089480205, -0.0027321934211120024, -0.0029450301441730146, 
    -0.0031441007753066096, -0.0033291949054340439, -0.0035006667201276142, 
    -0.0036595741370954167, -0.0038077696797819828, -0.0039479314408639972, 
    -0.0040835017174433198, -0.004218505862317124, -0.0043572677333120705, 
    -0.0045040547031970045, -0.0046626738863471831, -0.0048360793005258612, 
    -0.0050260304685634987, -0.005232850174877699, -0.0054553076626969298, 
    -0.0056906442090842065, -0.0059347240354629335, -0.0061822925646686034, 
    -0.0064273280349769991, -0.0066634356973827163, -0.0068842661224383268, 
    -0.0070839471384714974, -0.0072574846398381137, -0.0074011222384206881, 
    -0.007512617659336196, -0.0075914212610465118, -0.0076387220321508693, 
    -0.0076573584936844002, -0.0076515651247977805, -0.0076265859996426004, 
    -0.0075881873058023606, -0.0075421172832077265, -0.0074935756409063971, 
    -0.007446772411034067, -0.0074046194269458149, -0.0073685915494117495, 
    -0.0073387429554637434, -0.0073138899711227678, -0.0072919027390280257, 
    -0.0072700792543893477, -0.00724554000979186, -0.0072155993335103761, 
    -0.0071781034306734135, -0.0071316601639362827, -0.0070757895427189911, 
    -0.0070109475696900139, -0.0069384433029096235, -0.0068602479410970378, 
    -0.0067787048377674648, -0.0066961867397908629, -0.00661471421049987, 
    -0.0065356273277883672, -0.0064593426043506293, -0.0063852911676121459, 
    -0.0063120225798320006, -0.0062374410660855492, -0.0061591278796732799, 
    -0.0060746688754229911, -0.0059819565299858869, -0.0058794159844775254, 
    -0.0057661735975472906, -0.0056421239951551195, -0.00550791312769642, 
    -0.0053648320628109248, -0.0052146341101035835, -0.0050593035345185581, 
    -0.0049007866493563368, -0.004740774714706888, -0.0045805296774638279, 
    -0.0044208033003622551, -0.0042618641782345111, -0.0041036041901460155, 
    -0.0039457115386402498, -0.0037878513076343694, -0.0036298300252489749, 
    -0.0034717060321864291, -0.0033138263525943038, -0.0031568158864207969, 
    -0.0030015182387675204, -0.0028489165583206492, -0.0027000659327339515, 
    -0.0025560094611259301, -0.0024177182040678886, -0.0022860242081731304, 
    -0.002161584881535485, -0.002044843911306285, -0.0019360241357695045, 
    -0.0018351199159801603, -0.0017419228039594421, -0.0016560247677864957, 
    -0.0015768429298076661, -0.0015036189395654129, -0.0014354081617626536, 
    -0.0013710591617227949, -0.0013091994383468255, -0.0012482252142275571, 
    -0.0011863197810614966, -0.0011215066216450997, -0.0010517413245431225, 
    -0.00097502001036038513, -0.00088951844344555171, 
    -0.00079371478096575837, -0.00068651115529471166, 
    -0.00056733714963094132, -0.00043623302512554114, 
    -0.00029389457868740068, -0.00014171365192825836, 1.823772516072286e-05, 
    0.00018323473437071973, 0.00034997185682097639, 0.00051466049240154262, 
    0.00067314764189058184, 0.00082104621257045188, 0.00095386986401944885, 
    0.0010671420870113756, 0.0011564964030092724, 0.0012177659044234816, 
    0.0012470562539321664, 0.001240842066712725, 0.0011960755390701943, 
    0.0011103886742568072, 0.000982320570104125, 0.00081160548781477801, 
    0.00059944100034326885, 0.00034871148529024855, 6.4094649205170742e-05, 
    -0.00024796711033140979, -0.00057944031232986279, 
    -0.00092102537033507859, -0.0012626244863412493, -0.0015938916499773433, 
    -0.0019048579060830602, -0.0021865732802624164, -0.0024316617442683274, 
    -0.0026347546347357913, -0.0027927329194101826, -0.0029047150182422194, 
    -0.0029718661592539738, -0.0029970385023816533, -0.0029843586482173022, 
    -0.002938799053059122, -0.002865808274280404, -0.0027709652947994902, 
    -0.0026596766258673238, -0.0025368427996211021, -0.0024065256684393486, 
    -0.0022716586747833578, -0.0021338718041616941, -0.0019935003523504973, 
    -0.001849749539123733, -0.0017010081994898254, -0.0015452463224440273, 
    -0.0013804660618640758, -0.0012051422127940874, -0.0010186216802963331, 
    -0.00082142490485653038, -0.00061543355710948406, -0.0004039175367583892, 
    -0.00019141678184702568, 1.6496960785509053e-05, 0.00021356002801416803, 
    0.00039320946833793961, 0.00054898587275601296, 0.00067495307078402019, 
    0.0007660807621185789, 0.00081859858574777355, 0.00083028772431177622, 
    0.00080068975767767477, 0.00073120516398003893, 0.00062507553163785321, 
    0.00048725586225826015, 0.00032416162176781812, 0.00014333326952816814, 
    -4.6955361138412056e-05, -0.00023812197789006064, -0.0004216848038648831, 
    -0.00058964801617477215, -0.0007348803175299183, -0.00085141722558136569, 
    -0.00093470307986761713, -0.00098175807880174822, 
    -0.00099121479528967594, -0.00096326745742077321, 
    -0.00089951852072472221, -0.00080274938240547811, 
    -0.00067666085591903242, -0.00052559921728460835, 
    -0.00035428085882344531, -0.00016753520809794427, 2.9925366559569139e-05, 
    0.00023371881899766835, 0.00043996688955365835, 0.00064546953411648571, 
    0.00084779812369370456, 0.0010454043203921223, 0.0012376281545968472, 
    0.0014246628180312835, 0.0016074720676372278, 0.0017876261175250486, 
    0.001967099584531029, 0.0021480358521201197, 0.0023324984247504793, 
    0.0025222170029459709, 0.0027183650675422629, 0.0029213675408575395, 
    0.0031307580431796525, 0.003345085147753485, 0.003561872481279284, 
    0.0037776338952940744, 0.0039879572142169977, 0.0041876421592195968, 
    0.0043709203825328955, 0.004531693644980469, 0.0046637876683152408, 
    0.0047611615702056586, 0.0048180720179987211, 0.004829170476833111, 
    0.0047895856889778946, 0.0046950118454701832, 0.0045419019003879232, 
    0.0043277190153226657, 0.0040512363794112036, 0.0037128510766538804, 
    0.0033147607644905606, 0.002861031767130132, 0.0023574978728619859, 
    0.0018115707734885182, 0.0012319889645238575, 0.00062854913527220875, 
    1.1838110735930155e-05, -0.00060707693121479236, -0.0012169662550898046, 
    -0.0018067745051684747, -0.0023659549492658291, -0.0028847822445633611, 
    -0.0033546196655210299, -0.003768151198255203, -0.0041195353444014766, 
    -0.0044045265343357143, -0.0046205466427002807, -0.0047667434189651468, 
    -0.0048440288972711196, -0.0048550696000485456, -0.0048042576902509286, 
    -0.0046975902959624219, -0.004542507046771933, -0.0043476431213989109, 
    -0.0041225249511420677, -0.0038772508063993757, -0.0036220988440680154, 
    -0.0033671666286615039, -0.0031220093257623414, -0.002895303937996033, 
    -0.0026945763461534728, -0.002525988466834001, -0.0023941698862375003, 
    -0.0023021316444241159, -0.0022512199674156325, -0.0022411259824505819, 
    -0.0022699723537681245, -0.0023344367844087559, -0.0024299399988813512, 
    -0.0025508457074838791, -0.0026907097937465662, -0.0028425729606315294, 
    -0.0029992925339566412, -0.0031538664299647096, -0.0032997804258047083, 
    -0.0034312910845523464, -0.0035436378748588417, -0.0036331809216123166, 
    -0.0036973985668349403, -0.0037348012824676259, -0.0037447347539754129, 
    -0.0037271423341280066, -0.003682284159098631, -0.0036105033906104356, 
    -0.003512035510140424, -0.0033869121329551241, -0.0032349314311761242, 
    -0.003055729185368086, -0.0028489107956136944, -0.0026142367457453494, 
    -0.0023518165525576312, -0.0020623083038167882, -0.0017470944853199906, 
    -0.0014084047002750498, -0.0010493871824079324, -0.00067407313417008874, 
    -0.0002872195435554099, 0.00010597242483275553, 0.00050024925086415489, 
    0.00089075254367106886, 0.0012734712288927246, 0.0016455602055192821, 
    0.0020055552191357816, 0.0023533403920418978, 0.0026899699768989501, 
    0.0030172959080394142, 0.0033375491681161187, 0.0036529097617150758, 
    0.0039650870478878542, 0.0042749946168057652, 0.0045825158375801221, 
    0.0048863449656375221, 0.0051839384805504466, 0.0054715143329464849, 
    0.0057441549238909685, 0.0059959464974307028, 0.0062202021929324142, 
    0.0064097294707325019, 0.0065571880855302377, 0.0066553933723705648, 
    0.0066976923618226056, 0.0066782944640001634, 0.0065925075851703298, 
    0.0064369751570022898, 0.0062098113700800265, 0.0059106683531633432, 
    0.0055407985715848424, 0.0051030267421366231, 0.0046017473971688427, 
    0.0040428921366706073, 0.0034338397147039698, 0.0027832959196112251, 
    0.0021010399869143574, 0.0013975908727232376, 0.00068379124121526066, 
    -2.9586519446801447e-05, -0.0007322577282678212, -0.0014147331622953914, 
    -0.0020685338167096218, -0.0026863237283314867, -0.0032619258652532958, 
    -0.003790226396001586, -0.0042670436237159885, -0.0046889855569099206, 
    -0.0050532928310628149, -0.0053577750815853352, -0.0056007752647287516, 
    -0.0057812554194713282, -0.0058989144233340552, -0.0059543254180694028, 
    -0.0059490814510039566, -0.0058858319027940108, -0.0057682166531899401, 
    -0.0056007139128305015, -0.0053883727783411266, -0.005136514368279871, 
    -0.0048504769961718441, -0.0045353945584216786, -0.0041960752108191066, 
    -0.0038369399088889799, -0.0034620136154860206, -0.0030749196664161976, 
    -0.0026788365601920416, -0.0022764325552594535, -0.0018697222425938128, 
    -0.0014599363268644604, -0.0010473581660385754, -0.00063119462590726543, 
    -0.0002095208178285306, 0.00022070613101252327, 0.00066350034847426314, 
    0.0011235730845405776, 0.0016059471017368758, 0.0021154552389076428, 
    0.0026561571343425485, 0.0032307610382556308, 0.0038401197937689767, 
    0.0044828822336206407, 0.0051553191332191694, 0.0058513878461165913, 
    0.0065629409381756905, 0.0072800461508242646, 0.007991425532815899, 
    0.0086849282963265724, 0.0093480393813308877, 0.0099684280230853441, 
    0.01053448899693547, 0.011035883771232465, 0.011464004788719182, 
    0.011812382222065518, 0.012076946771058283, 0.012256157879050315, 
    0.012350957985236848, 0.012364598101439882, 0.012302318434112782, 
    0.012170939460475882, 0.011978448332435596, 0.011733541765979781, 
    0.011445255465530466, 0.011122666811964574, 0.010774693045236471, 
    0.01040997341287824, 0.010036772484168819, 0.0096629210962451834, 
    0.0092957486872145695, 0.0089419849082279079, 0.0086076416015092704, 
    0.0082978648244311087, 0.008016765873182995, 0.0077672303030489635, 
    0.0075508057334253047, 0.0073675508118263037, 0.007216028895597938, 
    0.0070933254103843508, 0.006995151225317223, 0.0069160403393502485, 
    0.0068495929425610377, 0.0067887499447522801, 0.0067260843583257816, 
    0.0066540396916000607, 0.0065651507749504706, 0.0064521596464503185, 
    0.0063081195110102524, 0.0061264857463287185, 0.0059012283266319651, 
    0.0056269535979239964, 0.005299091590258237, 0.0049140649341504385, 
    0.0044694154908290545, 0.0039640020572602524, 0.0033981007594987298, 
    0.0027735489600835845, 0.0020939038762246352, 0.0013645450632447827, 
    0.00059280830199697496, -0.00021196761576389612, -0.0010385451787281001, 
    -0.001874112729585156, -0.0027047590996120796, -0.0035161955642938518, 
    -0.004294553590325375, -0.0050271808984790499, -0.0057032922778409711, 
    -0.0063144625115303145, -0.0068548039695121498, -0.0073208968375893056, 
    -0.0077114655282242758, -0.0080269124321364054, -0.0082687356144407892, 
    -0.0084389389027531465, -0.0085395525577187555, -0.0085722553664822482, 
    -0.0085381610266632366, -0.0084377588105318119, -0.008271038787686421, 
    -0.0080377248135102986, -0.0077376422417482016, -0.0073711149736542057, 
    -0.0069394022152115108, -0.0064451095445834748, -0.0058924912347517976, 
    -0.0052876870956126325, -0.0046387528117782699, -0.0039555709934534361, 
    -0.0032495697612255946, -0.0025333838694272439, -0.0018204053757849589, 
    -0.0011243445912016425, -0.00045871576957907739, 0.00016360099931356256, 
    0.00073080503793919991, 0.001232546871323862, 0.0016601963085859427, 
    0.0020070042370492831, 0.0022681884492017717, 0.0024408532611460906, 
    0.0025238723533574105, 0.0025176576828587313, 0.0024239489382345803, 
    0.0022455835461825465, 0.0019863022817320618, 0.0016506063058856816, 
    0.0012436532760274372, 0.00077123298351449354, 0.00023981234192823339, 
    -0.0003434080644192924, -0.0009703855598048438, -0.0016321520671329307, 
    -0.0023186992359295693, -0.0030189280363085718, -0.0037205987504182977, 
    -0.0044103937967557953, -0.0050740665544698757, -0.0056967253397932184, 
    -0.0062632608013234699, -0.0067588860340985326, -0.0071697962672416619, 
    -0.0074837901871884901, -0.0076909640007560356, -0.0077843004754755384, 
    -0.007760164653731659, -0.0076187392073665452, -0.0073642600133416863, 
    -0.0070051758699979979, -0.0065540899348167135, -0.0060274731494745874, 
    -0.0054451158232609069, -0.0048292415401140461, -0.0042032587707323561, 
    -0.0035903889142650039, -0.0030122156215258403, -0.0024875057805276444, 
    -0.0020315018786055705, -0.0016558257940987573, -0.0013687626142301088, 
    -0.0011756479648311069, -0.0010790168716156197, -0.0010783145135714052, 
    -0.001169422372289456, -0.001344301659190467, -0.0015911158428604227, 
    -0.0018949051265370466, -0.0022387092044414752, -0.0026048846245271765, 
    -0.0029763484208050221, -0.0033375172083820823, -0.0036748217796139732, 
    -0.0039769521137676704, -0.0042348049970950541, -0.0044414698569382356, 
    -0.0045921428358646019, -0.0046841351867583543, -0.0047167778724423754, 
    -0.0046912841247606293, -0.0046105082746867891, -0.004478611104821611, 
    -0.004300768367594931, -0.0040828649709197459, -0.0038313997794530712, 
    -0.0035533531663504651, -0.0032561782916677561, -0.0029476554864714716, 
    -0.0026357058559037831, -0.0023279824973451661, -0.0020314188722495557, 
    -0.0017516177146530828, -0.0014923012401298497, -0.0012549356352163756, 
    -0.0010384513167744519, -0.00083934262941062592, -0.00065196956173963589, 
    -0.00046906245224848976, -0.00028239452393959022, 
    -8.3488426653444234e-05, 0.00013573161246967935, 0.00038238571977594296, 
    0.00066225292633484748, 0.00097952015724079287, 0.0013366711897358429, 
    0.00173441881693954, 0.0021716473829467941, 0.0026452810792159014, 
    0.0031502633856051272, 0.0036795836100968564, 0.0042244765473203778, 
    0.004774830195340544, 0.0053196643811868321, 0.0058476393671421144, 
    0.0063475663851424819, 0.0068088270602942487, 0.0072218625047546434, 
    0.0075785464765577449, 0.0078726399489877311, 0.0081001158310088292, 
    0.008259391084993491, 0.0083514776187829202, 0.0083799484047914971, 
    0.0083507117134614759, 0.00827169087322795, 0.008152333115001853, 
    0.0080031193742356004, 0.0078350927975394027, 0.0076594472272771058, 
    0.0074872161027839425, 0.0073291153427607033, 0.0071954402367806324, 
    0.0070959691293492758, 0.0070398333971528719, 0.0070352704825318649, 
    0.007089382083347244, 0.0072078291957127002, 0.0073946089003748446, 
    0.0076518540588539465, 0.0079798259065034984, 0.0083769427416648667, 
    0.0088399618598674779, 0.0093641157710672562, 0.0099434083658658974, 
    0.010570732822487819, 0.011238003465794358, 0.011936200637831764, 
    0.012655424946245693, 0.013384921502241003, 0.014113194499961989, 
    0.014828262414490116, 0.015518039230318567, 0.016170799501366115, 
    0.016775613680827677, 0.017322983559269055, 0.017805370989230154, 
    0.018217563213753139, 0.018557050124430843, 0.018824435991839545, 
    0.019023536870849973, 0.019161462794978792, 0.019248509309962893, 
    0.019297809491816777, 0.01932484935166957, 0.019346877476511842, 
    0.019382246215844404, 0.019449522125325983, 0.0195665281055563, 
    0.019749004425042904, 0.020009342490553972, 0.020355256969312771, 
    0.020788842890004391, 0.021305913076951764, 0.021895945903310357, 
    0.022542529823800513, 0.023224257758943691, 0.023915940590012539, 
    0.024589820001021112, 0.025216848553245037, 0.025767885632577772, 
    0.026214531090965248, 0.026530212451272954, 0.026691093766774792, 
    0.026676934535265737, 0.026472126692317105, 0.026066575112106558, 
    0.025456536352859081, 0.024645515787921408, 0.023644806293343999, 
    0.022473947050530116, 0.02116066917527467, 0.019740117132393389, 
    0.018253722016100378, 0.016747117940193981, 0.015267544340684364, 
    0.013861006444702364, 0.012569283947732948, 0.011427012991727516, 
    0.010459213935575145, 0.0096792204711308016, 0.0090873351006012688, 
    0.0086706200974861168, 0.0084030913796589307, 0.0082474067482921562, 
    0.0081572000939527187, 0.0080802715186417528, 0.0079623588307905762, 
    0.0077512811023223386, 0.0074009245749372199, 0.0068756181213229005, 
    0.0061532245127120973, 0.0052281742676659557, 0.0041129681617652928, 
    0.0028378732945958359, 0.0014488260221955313, 3.4201921840035926e-06, 
    -0.0014344250910503197, -0.0028013728812624414, -0.0040406554867100323, 
    -0.0051064455482983315, -0.0059669542082998548, -0.0066039284461092435, 
    -0.0070123392697914308, -0.0071982561048545401, -0.0071761757006036341, 
    -0.0069692106111981468,
  // Fqt-Na(7, 0-1999)
    1, 0.99388955835474724, 0.97581639143519294, 0.94653265328365088, 
    0.90722500109081805, 0.8594247419217107, 0.80489762203258208, 
    0.74552546291263466, 0.68319144741561499, 0.61967901993816554, 
    0.55659144711334962, 0.4952957284439311, 0.43689141914204466, 
    0.38220233354492078, 0.33178721788909848, 0.28596460264046386, 
    0.24484677459161244, 0.20837822957893259, 0.17637469572141343, 
    0.14855988295202482, 0.12459797543247829, 0.10412087616369443, 
    0.086749890444285757, 0.072112079401519522, 0.05985187937394134, 
    0.049638697239728115, 0.041171274438875416, 0.034179585226673567, 
    0.028424935433487904, 0.023698866377678405, 0.019821305054491811, 
    0.016638296086510122, 0.014019561076422561, 0.011855983471525625, 
    0.010057128034648635, 0.0085488254199887117, 0.0072708725284001746, 
    0.0061748941355030647, 0.0052223971304028753, 0.0043830715968713185, 
    0.0036333223825218731, 0.0029550425854330724, 0.0023345803518361715, 
    0.0017618694815430148, 0.0012296830303476925, 0.00073296798823543853, 
    0.00026825990664793925, -0.00016684388139221072, -0.0005741317568937357, 
    -0.00095515500299898557, -0.001311495253763683, -0.0016449222847335814, 
    -0.0019574383133881407, -0.0022512200945550183, -0.002528478273607367, 
    -0.0027912863180332937, -0.0030414084848555353, -0.003280172403640555, 
    -0.003508426430493847, -0.0037265763220278212, -0.0039347125232103994, 
    -0.0041327830991422692, -0.0043207911586826582, -0.0044989484717195974, 
    -0.0046677888894136139, -0.0048281679989737886, -0.0049812014049141172, 
    -0.0051281041111929373, -0.0052699964232784582, -0.0054076977781384429, 
    -0.0055415511745251335, -0.005671302337928159, -0.0057960496495346441, 
    -0.0059142405861009346, -0.0060237122255255206, -0.0061217490592586571, 
    -0.0062051497702873453, -0.0062703028214775918, -0.0063132718375706071, 
    -0.0063299143098065579, -0.0063160272872826205, -0.0062675529755421714, 
    -0.0061808103922483997, -0.0060527698487924022, -0.005881333813614437, 
    -0.005665608457836863, -0.0054061289445610332, -0.0051050381760527237, 
    -0.0047661858368737257, -0.0043951315487976714, -0.0039990632613537839, 
    -0.0035866087704021091, -0.0031675658413754756, -0.0027525590529085993, 
    -0.0023526440728381844, -0.0019788743550649248, -0.0016418618422558184, 
    -0.0013513454167402722, -0.0011158003384703515, -0.00094210718705413019, 
    -0.00083529784475809533, -0.00079840793055683331, 
    -0.00083242378580606583, -0.00093632955193948366, -0.0011072352619386639, 
    -0.0013405607843702742, -0.0016302580542344944, -0.0019690335921543128, 
    -0.0023485616736672408, -0.0027596711321517193, -0.003192514635023091, 
    -0.0036367189944403926, -0.0040815363441465587, -0.0045160310751483617, 
    -0.0049292829359643409, -0.005310657920876323, -0.0056501115085974768, 
    -0.005938540527885036, -0.006168134557800747, -0.0063327204438790472, 
    -0.0064280376343640267, -0.0064519152113058495, -0.0064043217204671817, 
    -0.0062872624380844594, -0.0061045274461522803, -0.0058613446707646549, 
    -0.0055639575179499698, -0.005219213734571136, -0.0048342107243482127, 
    -0.0044160385456338954, -0.0039716382544668499, -0.003507773232095778, 
    -0.0030310716752740365, -0.0025481268082464632, -0.0020655916890158247, 
    -0.0015902660120019588, -0.0011291365641345604, -0.00068935142328098095, 
    -0.00027814384092606035, 9.7306235631945941e-05, 0.00043007300770856529, 
    0.0007137057145131737, 0.00094248939544464342, 0.0011116999801946044, 
    0.0012178409288510525, 0.0012588345643311815, 0.0012341582074453217, 
    0.0011448870806562291, 0.00099366585033693229, 0.0007846042623146811, 
    0.00052310746494085912, 0.00021567090612043877, -0.00013035430034695386, 
    -0.00050701598129248193, -0.00090601202981974789, -0.0013189469801872706, 
    -0.0017375621592839617, -0.0021539494290826974, -0.0025607265805511026, 
    -0.0029511907871174921, -0.0033194481223390187, -0.0036605320373372567, 
    -0.0039704886343506027, -0.0042464388917747417, -0.0044865693639545203, 
    -0.0046900731491315009, -0.004857032185393551, -0.0049882751185638292, 
    -0.0050851973937317881, -0.005149576532268987, -0.0051833655684957874, 
    -0.0051885058910762149, -0.0051667806382068148, -0.0051197252858228223, 
    -0.0050486299612678923, -0.0049546208434512193, -0.0048388068193661541, 
    -0.0047024656643229364, -0.004547232476290743, -0.0043752465715738639, 
    -0.0041892341916680764, -0.0039924874054498918, -0.0037887496942943196, 
    -0.0035819971532531155, -0.0033761701029412735, -0.0031748725631615365, 
    -0.0029810998254676153, -0.0027970350651668908, -0.0026239391205654132, 
    -0.002462146587238387, -0.0023111672890714328, -0.0021698682093865031, 
    -0.0020366992093092517, -0.001909946938387766, -0.0017879551620536374, 
    -0.0016693087430891648, -0.001552945691600268, -0.0014381917977930327, 
    -0.0013247274747493192, -0.0012124886162568757, -0.0011015414923523921, 
    -0.00099195415843086041, -0.00088370392024597578, 
    -0.00077663648370434658, -0.00067048646695268656, 
    -0.00056496572531725662, -0.00045987670297107459, 
    -0.00035524385899595671, -0.00025142273106075236, -0.0001491542753579338, 
    -4.9561733204422356e-05, 4.5931606737413164e-05, 0.00013574500741021545, 
    0.00021833381807321136, 0.00029240604507999306, 0.0003571336898799922, 
    0.00041233245511205639, 0.00045858604570320341, 0.00049729401891982308, 
    0.00053062586054164625, 0.00056141012462125931, 0.00059293503625120945, 
    0.00062871085160836108, 0.00067220964680520781, 0.00072660372668243106, 
    0.00079455326212213404, 0.00087804368687915914, 0.00097829440121882053, 
    0.0010957390294095799, 0.0012300610688993276, 0.00138026458209064, 
    0.001544754660074083, 0.0017213958127529527, 0.001907539459932092, 
    0.0020999999105107466, 0.0022949982764904416, 0.0024880875850537493, 
    0.0026740856597276272, 0.0028470558473216948, 0.0030003716889795166, 
    0.0031268856443707757, 0.0032192156325629956, 0.0032701360978737606, 
    0.0032730428724951086, 0.0032224406784907987, 0.0031144072926339635, 
    0.0029469699958414464, 0.0027203609713977121, 0.002437118150657374, 
    0.0021020298411481586, 0.0017219439225707033, 0.0013054496915635315, 
    0.00086247718891712625, 0.00040383110164727805, -5.931342760483562e-05, 
    -0.00051592378603129957, -0.00095559664528154908, -0.0013689938886493737, 
    -0.0017481736562512534, -0.0020867999704757599, -0.002380210304014036, 
    -0.0026253477353556614, -0.0028205801828442493, -0.0029654716135376303, 
    -0.0030605335376075972, -0.0031070142183428498, -0.0031067406865007163, 
    -0.0030620035762687313, -0.0029755050882168833, -0.0028503245762518197, 
    -0.0026899103698074175, -0.0024980708674117854, -0.0022789736215470193, 
    -0.0020371198163291072, -0.0017773089086575438, -0.0015045662407750962, 
    -0.0012240453017988762, -0.00094089956421230202, -0.00066012726463125651, 
    -0.00038641382538971551, -0.00012397187978610395, 0.0001235848833805453, 
    0.0003533455757966928, 0.00056315142824581838, 0.00075160380161468174, 
    0.00091803357022332685, 0.001062435889645805, 0.0011853934887308991, 
    0.0012879958567620594, 0.0013717681241842022, 0.0014386128912925852, 
    0.001490769235438436, 0.0015307780518904143, 0.0015614468782727078, 
    0.0015857929544666361, 0.0016069620707859563, 0.0016281073945047934, 
    0.0016522335143987221, 0.0016820037660952064, 0.0017195407349645518, 
    0.0017662302232495624, 0.0018225573982001081, 0.0018879860630369358, 
    0.0019609154907919051, 0.0020387033671494187, 0.0021177679110561272, 
    0.0021937435681200412, 0.0022616991973727881, 0.002316394223507226, 
    0.0023525650863865238, 0.0023652324086439287, 0.0023500126679911956, 
    0.0023033991119653621, 0.0022229954873502831, 0.0021076787431034269, 
    0.0019576751095923143, 0.001774554130503449, 0.001561170618750976, 
    0.0013215509134718603, 0.0010607644700028076, 0.0007847692388499351, 
    0.0005002272440908053, 0.00021428187524534021, -6.5711466731866678e-05, 
    -0.00033248182657082706, -0.00057915097687195167, 
    -0.00079950424716046216, -0.00098820291115583989, -0.0011409202108118072, 
    -0.0012544010464021656, -0.0013264656083387507, -0.0013559747368986144, 
    -0.0013427855888896829, -0.0012876900093025476, -0.0011923509929703145, 
    -0.0010592205091061455, -0.00089143523364765016, -0.00069270770725803413, 
    -0.00046721223551917724, -0.00021948526770337664, 4.5678195203385389e-05, 
    0.00032330881203416014, 0.00060834382295687638, 0.00089571238833551447, 
    0.001180406055231986, 0.0014575265503128981, 0.0017223158786249517, 
    0.0019701651757963634, 0.0021966242405625103, 0.0023974474514403404, 
    0.0025686916676051119, 0.0027068736085746467, 0.0028091960991609597, 
    0.0028737829795584743, 0.0028998827537653499, 0.0028879936016796993, 
    0.0028398554154999175, 0.0027583244979474341, 0.002647117167919961, 
    0.0025104889388967789, 0.0023528608483692095, 0.0021784802661559436, 
    0.0019911249309087415, 0.0017938941266359277, 0.001589101920863923, 
    0.001378278449668167, 0.0011622609741666796, 0.00094137890718448312, 
    0.00071570766374506151, 0.0004853700088308468, 0.00025084069018231397, 
    1.3231842914960293e-05, -0.0002255049546828598, -0.00046246917974263546, 
    -0.00069382774877860156, -0.00091493633427815993, -0.0011205492926605416, 
    -0.0013050823440211253, -0.0014629065501833788, -0.0015886576099080601, 
    -0.0016775416520058571, -0.001725641427776838, -0.0017301995628061996, 
    -0.0016898787926904963, -0.0016049579546508724, -0.0014774429201908541, 
    -0.0013110721647326389, -0.0011111959953343338, -0.00088455909167314611, 
    -0.00063898390269098541, -0.0003830040980265972, -0.00012547405477677717, 
    0.00012482242143481339, 0.00035954673047829371, 0.00057114489323162386, 
    0.00075314214045925408, 0.00090038439947696686, 0.0010092250888995217, 
    0.0010776453682427977, 0.0011053115503794285, 0.001093548781317059, 
    0.0010452597175846703, 0.00096476112498495431, 0.00085756467920939934, 
    0.00073009952260794586, 0.00058938187707613518, 0.00044266315746633006, 
    0.00029706949491536906, 0.00015925988891516633, 3.5145854250230113e-05, 
    -7.032042589080181e-05, -0.00015325350023024959, -0.00021085436211667032, 
    -0.0002413272503546392, -0.00024374297292061606, -0.00021787075824983564, 
    -0.00016400899532444937, -8.2865157890834305e-05, 2.451653326834499e-05, 
    0.00015677744589726158, 0.00031221574236505389, 0.00048873238216529092, 
    0.0006837795586348926, 0.0008943174111875939, 0.0011168081485718631, 
    0.0013472493378132197, 0.0015812546096801901, 0.0018141644723181289, 
    0.0020411876263489673, 0.0022575462156053613, 0.0024586396434540152, 
    0.0026401916499030655, 0.0027984020548863981, 0.0029300732518055279, 
    0.0030327331462552875, 0.0031047301177056052, 0.0031453149141768928, 
    0.0031546881998521354, 0.0031340216933033625, 0.0030854374608925298, 
    0.0030119449782301621, 0.0029173219503823493, 0.0028059482599601801, 
    0.0026825833881889073, 0.002552120132766812, 0.0024193447645363066, 
    0.0022886954250294026, 0.0021640848800470475, 0.0020487590498875071, 
    0.0019452140064044393, 0.0018551524011273602, 0.0017794723609353027, 
    0.001718297494194256, 0.0016710553872313308, 0.0016365745899391865, 
    0.0016131769340831442, 0.0015987376243958126, 0.0015907213367189279, 
    0.0015862184063695421, 0.0015820306142932876, 0.0015748140966073704, 
    0.0015612892161968432, 0.0015384888911372998, 0.0015039842309666435, 
    0.0014560557958658491, 0.0013937891194158777, 0.0013170744303287298, 
    0.0012265340556428693, 0.0011233893855699343, 0.0010093153336092095, 
    0.00088628223944251427, 0.00075641265638264218, 0.00062185480830052159, 
    0.00048467102218080721, 0.00034675619891678868, 0.00020977630527825814, 
    7.5126450306279175e-05, -5.6078744757875854e-05, -0.00018300062005174465, 
    -0.00030504808302920378, -0.00042183542840763165, 
    -0.00053312881590303189, -0.00063878142979394517, 
    -0.00073867596781521181, -0.00083265474689161773, 
    -0.00092046982391705149, -0.0010017275737657675, -0.0010758417274353083, 
    -0.0011419905222938473, -0.0011990813694623943, -0.0012457428910143343, 
    -0.0012803481261265039, -0.0013010928278747193, -0.0013061159555405647, 
    -0.0012936587555844657, -0.001262223893908995, -0.0012107292454680257, 
    -0.0011386085809872823, -0.0010458732557708005, -0.00093311875877516719, 
    -0.00080149497456846719, -0.00065262628734065096, 
    -0.00048852800495432472, -0.00031148355016330981, 
    -0.00012393702881044379, 7.1620875460329443e-05, 0.00027273830182707518, 
    0.00047705334550335332, 0.00068231195904518063, 0.00088633615657911463, 
    0.0010869933299384816, 0.0012821663069492938, 0.0014697606813582733, 
    0.0016477620989872811, 0.0018143207218476571, 0.0019678684072995433, 
    0.0021072237461057727, 0.0022316781136259454, 0.0023410459685284735, 
    0.002435660238946852, 0.0025163162818730741, 0.0025841636214517286, 
    0.0026405748106703257, 0.0026869834607155412, 0.002724739261968962, 
    0.0027549978061824189, 0.0027786638304947977, 0.0027963948518310933, 
    0.0028086690613055004, 0.0028159073440749073, 0.0028186079855654455, 
    0.0028174770673509049, 0.0028135090685081666, 0.0028079899325151574, 
    0.0028024226597134858, 0.0027983806707578942, 0.0027973075971948311, 
    0.0028003046334035718, 0.0028079276271343449, 0.0028200200955565092, 
    0.0028356149087190039, 0.0028528914534816339, 0.0028692018089169552, 
    0.0028811541923357185, 0.0028847462126824828, 0.0028755391128578735, 
    0.0028488891741801844, 0.0028002192757432412, 0.0027253551698232219, 
    0.0026208773824761122, 0.0024844913853639414, 0.002315363608619858, 
    0.002114362732320533, 0.0018841935848535587, 0.0016293760420658971, 
    0.0013560772365780215, 0.0010718025180630844, 0.00078499838315607931, 
    0.00050460388193019528, 0.0002395681934184556, -1.6280321926792326e-06, 
    -0.0002114241714757451, -0.00038358088076574897, -0.00051348204958538625, 
    -0.00059833213467965808, -0.00063722086920261914, 
    -0.00063107125086090494, -0.00058245500999982937, 
    -0.00049531731828791816, -0.00037462228304230158, 
    -0.00022595773379071503, -5.5131682387158645e-05, 0.00013219800317569762, 
    0.00033083570176651298, 0.00053626908337997992, 0.00074479326751298669, 
    0.00095353214217781237, 0.0011603778248154943, 0.0013638621242373606, 
    0.0015629900226857211, 0.0017570717658188665, 0.0019455757482585501, 
    0.002128009181087998, 0.0023038528305830133, 0.0024725311301115483, 
    0.0026334062675902078, 0.0027857904577904585, 0.0029289583596915367, 
    0.0030621557713472933, 0.0031845910839549151, 0.0032954215740646597, 
    0.0033937198980521525, 0.0034784345639924299, 0.0035483566779023956, 
    0.0036020901901105988, 0.0036380424190339518, 0.0036544469793177038, 
    0.0036494114291574574, 0.0036210204943796192, 0.003567462827557581, 
    0.0034871984259682151, 0.0033791559873764219, 0.0032429240845406339, 
    0.0030789298422424175, 0.0028885807177047602, 0.0026743377905227889, 
    0.0024397373682510013, 0.0021893274400471311, 0.0019285452663109848, 
    0.0016635287049823373, 0.0014008689188486473, 0.0011473210535369114, 
    0.00090946945846889196, 0.0006933876723940384, 0.00050429200222861827, 
    0.00034624720857291262, 0.00022193337196231561, 0.00013251467400718689, 
    7.7633317548670105e-05, 5.5521804679995921e-05, 6.323245195394441e-05, 
    9.6936866538716184e-05, 0.00015228737827220279, 0.00022474466210291598, 
    0.00030986748023132321, 0.00040351696056808165, 0.00050196171911836608, 
    0.00060191991511153041, 0.0007005334874606126, 0.0007953144079201628, 
    0.00088406612272562293, 0.00096482937133093622, 0.0010358445397225312, 
    0.0010955803133076132, 0.0011428193669995427, 0.0011767974205554282, 
    0.0011973701311740882, 0.0012051645644912136, 0.0012016858845701884, 
    0.0011893412597478099, 0.0011713740099900849, 0.0011517136464524584, 
    0.001134748277314291, 0.0011250436893357816, 0.0011270355763202543, 
    0.0011447099421887682, 0.0011813002020371029, 0.0012390231747712935, 
    0.0013188698328649388, 0.0014204518172285863, 0.0015419413696187482, 
    0.0016800974767510095, 0.0018303810325699271, 0.0019871730990541473, 
    0.0021440786065828866, 0.002294292405572892, 0.0024310132885392026, 
    0.0025478595890570414, 0.0026392736768792203, 0.0027008563468884274, 
    0.0027296242979386806, 0.002724146336067892, 0.0026845641524003705, 
    0.0026124905070378434, 0.0025108142198780005, 0.0023834376539804613, 
    0.0022349728680544239, 0.0020704172958429055, 0.0018948489909893936, 
    0.0017131488580288739, 0.0015297716207063974, 0.0013485692094835737, 
    0.0011726929913670621, 0.0010045470413418132, 0.00084580879490834952, 
    0.00069747717355562685, 0.00055994046981284844, 0.00043304407985229377, 
    0.00031615452198848902, 0.00020822163512931535, 0.00010785181793801567, 
    1.3384179883775267e-05, -7.7023792257927893e-05, -0.00016530966397719824, 
    -0.00025342952351845282, -0.00034328276234014076, 
    -0.00043664936604029725, -0.00053510309485341851, 
    -0.00063989662226938103, -0.00075180480147735726, 
    -0.00087094010119177486, -0.00099656487163378351, -0.0011269537363047253, 
    -0.0012593402871349387, -0.0013899978810741147, -0.0015144422844987036, 
    -0.001627738304228434, -0.0017248602533455962, -0.0018010692021598288, 
    -0.0018523075848628965, -0.0018755608175929639, -0.0018691916360461841, 
    -0.0018332005112133367, -0.0017693644346985387, -0.001681247407647628, 
    -0.0015740528135235934, -0.0014543293958421103, -0.0013295488630987052, 
    -0.001207603166349771, -0.0010962626651459593, -0.0010026546731133287, 
    -0.0009328084240369332, -0.00089131264070918363, -0.00088110565752260383, 
    -0.00090340563878024661, -0.0009577695064120692, -0.0010422623222927591, 
    -0.001153702440142906, -0.0012879496505555418, -0.0014402076006223711, 
    -0.0016053130407136505, -0.0017779984756396022, -0.0019531157690976433, 
    -0.0021258084414744818, -0.002291655730335314, -0.0024467741097321475, 
    -0.0025878838143757149, -0.0027123599551680073, -0.0028182517386808369, 
    -0.0029042791632003955, -0.0029698169233079814, -0.0030148459903765424, 
    -0.0030399131567262518, -0.0030460795613374263, -0.0030348839621877244, 
    -0.0030083063386509919, -0.002968703856654441, -0.0029187365012057999, 
    -0.0028612286908138648, -0.0027990141458567007, -0.0027347605136559734, 
    -0.0026708088202346421, -0.0026090394054044765, -0.0025507910276947876, 
    -0.0024968216526803275, -0.0024473153880276897, -0.0024019149177662907, 
    -0.0023597586841769547, -0.0023195106043198688, -0.0022793694539194036, 
    -0.0022370745855867218, -0.0021899219962024422, -0.0021348200393146357, 
    -0.0020684196991201638, -0.001987334003300238, -0.0018884346331392327, 
    -0.0017691963738870639, -0.0016280147652346191, -0.001464461924077146, 
    -0.0012794350789524581, -0.0010751748684827709, -0.00085516108099008953, 
    -0.0006238851375168367, -0.00038652920365097411, -0.0001485802830894437, 
    8.4580894423134332e-05, 0.00030804893779576726, 0.00051768622410497357, 
    0.00071028808890972019, 0.00088362319050710732, 0.0010363296440821504, 
    0.0011677282857316131, 0.0012775761202199389, 0.0013658248930391375, 
    0.0014324093584857777, 0.0014771044255677385, 0.0014994489043753958, 
    0.0014987380742092673, 0.0014740757608299705, 0.0014244811242396973, 
    0.001349021403252007, 0.001246973852545224, 0.0011179956623736567, 
    0.00096229319932193073, 0.00078076447540872658, 0.0005751110874700889, 
    0.00034789192116838107, 0.00010251081158224601, -0.00015687156592718657, 
    -0.00042548511786978568, -0.0006981712269768989, -0.00096962736131610868, 
    -0.0012346823889467168, -0.001488565348406439, -0.0017271419429832897, 
    -0.0019471008601227616, -0.0021460806628292931, -0.002322709333453504, 
    -0.0024765760957628576, -0.0026081355981284718, -0.0027185705531090551, 
    -0.002809626214735812, -0.00288344086736016, -0.0029423717750734915, 
    -0.0029888386654907703, -0.003025195788935257, -0.0030536211794897875, 
    -0.0030760249672486988, -0.0030939872217518962, -0.0031087008023262591, 
    -0.0031209354527462251, -0.0031310013199731461, -0.0031387511366387216, 
    -0.0031435954890632134, -0.0031445570695212287, -0.0031403585741271436, 
    -0.0031295476801845613, -0.0031106373391395106, -0.0030822544312096994, 
    -0.0030432874008156866, -0.0029930097282795096, -0.0029311793868201149, 
    -0.0028580916878959504, -0.002774601741013781, -0.0026820933474952526, 
    -0.0025824081886750795, -0.0024777401006319789, -0.0023704935000506363, 
    -0.0022631190280440702, -0.0021579347443690857, -0.0020569269981303147, 
    -0.0019615557801255998, -0.0018725602365882955, -0.0017897842821340225, 
    -0.0017120517093560657, -0.0016371133529259603, -0.0015616728425177934, 
    -0.0014815210241225323, -0.0013917719159076618, -0.001287168049322131, 
    -0.0011624521846380846, -0.0010127500794529761, -0.00083396359028547204, 
    -0.00062309934742476474, -0.00037856226861657976, -0.0001003468169343952, 
    0.00020983480559484541, 0.00054852464201364721, 0.00091056522640355563, 
    0.0012892335743364498, 0.001676457046092714, 0.0020631143080249723, 
    0.0024394098933141805, 0.0027953084328253869, 0.0031210080442743574, 
    0.003407410884041711, 0.0036465606524013457, 0.003832026361890028, 
    0.0039591916777550933, 0.0040254625243238912, 0.0040303582962766347, 
    0.0039755211996674675, 0.0038646214323963604, 0.0037031876687450131, 
    0.0034983609375602771, 0.0032585999850980049, 0.0029933318186905035, 
    0.0027125361845891523, 0.0024263107356416336, 0.0021443978780806144, 
    0.0018757192054656225, 0.0016279559563033336, 0.0014071996936042806, 
    0.0012177127635541137, 0.0010618191711968057, 0.00093991413899910663, 
    0.00085059322536174442, 0.00079088257854627428, 0.00075652386708021193, 
    0.00074231917014690348, 0.00074246330148784929, 0.00075087893011915494, 
    0.00076151225878970624, 0.00076859045962458686, 0.00076683206552885172, 
    0.00075161895138687977, 0.00071912669821761659, 0.00066642145352339987, 
    0.00059152208470544311, 0.00049342284562108724, 0.00037206999246606267, 
    0.00022830451256913435, 6.3756581837368356e-05, -0.0001192955978988036, 
    -0.00031809150942344294, -0.00052956278700493466, 
    -0.00075050054929496712, -0.00097770077077196922, -0.0012080775708266679, 
    -0.0014387262970362808, -0.0016669511539561506, -0.0018902476783150708, 
    -0.0021062467052307384, -0.0023126414897684062, -0.0025070974044593972, 
    -0.0026871807277332382, -0.002850318449979954, -0.0029938349257591737, 
    -0.0031150465195673494, -0.0032114476893763066, -0.003280963868762048, 
    -0.003322223060887931, -0.0033348208684106043, -0.0033195245767488279, 
    -0.0032783738110365771, -0.0032146483793615531, -0.0031327231628860042, 
    -0.003037796237219012, -0.0029355338575240064, -0.002831672665024093, 
    -0.0027316025923239113, -0.0026399795020529233, -0.0025604144488419753, 
    -0.002495262386462898, -0.0024455385815090342, -0.0024109817358592195, 
    -0.0023902345078409002, -0.0023811237602762553, -0.0023809938722105946, 
    -0.002387052764062206, -0.0023966848605691802, -0.0024076850497773612, 
    -0.0024184169387263662, -0.0024278550063655427, -0.0024355232885742363, 
    -0.0024413554360650709, -0.0024454833977195383, -0.0024480058691176386, 
    -0.0024487550098623257, -0.0024471069157992104, -0.002441837368331604, 
    -0.0024310577484771565, -0.0024122103906284408, -0.0023821613220621611, 
    -0.002337352340064078, -0.0022740173421017082, -0.0021884336971008007, 
    -0.0020771962188889034, -0.0019374748052232845, -0.0017672790480425281, 
    -0.0015656859363199921, -0.0013330439770180807, -0.0010711335588817384, 
    -0.00078324639032369104, -0.00047416408257258376, 
    -0.00015001339208099682, 0.000182042016100298, 0.00051422679190453674, 
    0.00083868648189878189, 0.0011480593026235782, 0.0014360156780792196, 
    0.0016976953984739085, 0.001929997251786364, 0.0021316760356435175, 
    0.0023032513686803207, 0.0024467486146782409, 0.0025653190661675757, 
    0.0026627902552775976, 0.0027432335088709743, 0.0028105762919812898, 
    0.0028683337196802067, 0.0029194510056068912, 0.0029662661056782105, 
    0.0030105735420923201, 0.0030537665568925029, 0.0030969956362750816, 
    0.003141347639343618, 0.0031879706653575104, 0.0032381604497672485, 
    0.0032933707446429132, 0.0033551451865740313, 0.0034249998971035197, 
    0.0035042651154444369, 0.0035939204725568461, 0.0036944629155144962, 
    0.0038058312511894186, 0.0039273946808397716, 0.0040579693343878488, 
    0.004195879496566181, 0.0043390127139184154, 0.0044848858232700295, 
    0.0046307330246017318, 0.0047736081794072021, 0.0049105063261360741, 
    0.0050385155253581046, 0.0051549311865191514, 0.005257333428677873, 
    0.0053436119979655338, 0.0054119511605570502, 0.0054607882233021947, 
    0.0054887798778947058, 0.0054947844986639903, 0.0054778680575178172, 
    0.0054373433145849205, 0.0053727963273328778, 0.0052841309961823594, 
    0.0051715956333707597, 0.0050357988622818269, 0.0048777102598148757, 
    0.004698642200503509, 0.0045002087191097738, 0.004284271117197461, 
    0.0040528914787425182, 0.0038083189712086645, 0.003553055229374452, 
    0.0032899701909200585, 0.0030224686679091524, 0.0027546333242512351, 
    0.0024912911267603701, 0.0022379624032267849, 0.0020006644414269819, 
    0.0017855744912913954, 0.0015985928104132157, 0.0014448513717441674, 
    0.0013282310391176117, 0.0012509400441581037, 0.0012132240919786501, 
    0.0012132571817254109, 0.0012472392418371257, 0.0013097062883461767, 
    0.0013940438749220209, 0.0014931247590465602, 0.0016000314073333259, 
    0.0017087340234832717, 0.0018146668792264785, 0.0019150954758270422, 
    0.0020092461036412272, 0.002098171258225168, 0.0021843918699878694, 
    0.002271366465111641, 0.0023628775483795885, 0.0024624196611769626, 
    0.0025726596651947636, 0.0026950365418806424, 0.0028295275247472986, 
    0.0029745993409597835, 0.0031273422237938246, 0.0032837520862529705, 
    0.0034391276778844848, 0.0035885078557393547, 0.0037270906537612298, 
    0.003850589010654772, 0.0039554849157179724, 0.0040391769739853284, 
    0.0041000451042629673, 0.0041374464005756494, 0.0041516529397620143, 
    0.0041437710359944592, 0.0041155921712099069, 0.0040694208952862703, 
    0.0040078542708939999, 0.0039335332139260465, 0.0038489227754456286, 
    0.0037561035746556137, 0.0036566211996562504, 0.0035514132137048366, 
    0.0034407918779159235, 0.003324505432369197, 0.0032018766790619349, 
    0.0030719756699618054, 0.0029338347020936247, 0.0027866614826841103, 
    0.002630053178818165, 0.0024641678998433649, 0.0022898683937061948, 
    0.0021087964731343993, 0.0019233766956631866, 0.001736701756626266, 
    0.0015523120226738245, 0.0013738497431274785, 0.0012046299980634986, 
    0.0010471861467392775, 0.00090284486719614679, 0.00077140568854123376, 
    0.00065098100555648444, 0.00053804084964897503, 0.00042763702414194324, 
    0.00031380573216271241, 0.00019008224661342031, 5.0074478782253124e-05, 
    -0.00011196691062540203, -0.00030063003940937927, 
    -0.00051893599139075171, -0.00076806459137977821, -0.001047238951311095, 
    -0.0013537524203067919, -0.0016831066126615916, -0.0020292452360243093, 
    -0.0023848228905578193, -0.0027414993154630256, -0.0030902259884552697, 
    -0.0034215439804660243, -0.0037258622271009009, -0.003993735486343953, 
    -0.0042161393214619741, -0.0043847571914834458, -0.0044922577892510147, 
    -0.0045325792497968847, -0.0045012050304862683, -0.0043954152125287929, 
    -0.0042145179826302013, -0.0039600337196085827, -0.0036358175206138836, 
    -0.0032481038725637327, -0.0028054589920790663, -0.002318585195765287, 
    -0.0017999970658046632, -0.0012635416865195996, -0.00072379371293297256, 
    -0.00019535291743789831, 0.00030789809835328008, 0.00077349114076293588, 
    0.0011909720323360082, 0.0015523152330733309, 0.0018521434425977476, 
    0.0020877310451573542, 0.0022588142287755675, 0.0023672625046132403, 
    0.00241667576985299, 0.0024119437018101557, 0.0023588380464561335, 
    0.002263662498140283, 0.0021329787203990011, 0.0019734209580808439, 
    0.0017915984475931253, 0.0015940573631292312, 0.0013872759323136953, 
    0.0011776683910034004, 0.00097156092266059138, 0.0007751426017259277, 
    0.00059438016425501349, 0.00043491697808747942, 0.00030197051655959798, 
    0.00020022283072362933, 0.00013375181372794236, 0.00010598279634553798, 
    0.0001196576301367249, 0.00017681743159201789, 0.00027878251921736565, 
    0.00042607737095807591, 0.00061833969861182592, 0.00085417240543843071, 
    0.0011309936604392947, 0.001444874738112835, 0.0017904295826974774, 
    0.0021607625153152953, 0.0025475165946577502, 0.0029410344167714866, 
    0.003330635612080403, 0.0037050170108583135, 0.0040527401127149788, 
    0.0043628031117817299, 0.0046252427913048679, 0.004831728010493589, 
    0.0049760855135551306, 0.0050547299169273118, 0.0050669354331709946, 
    0.0050149281776584072, 0.0049037821470612466, 0.0047411337344756502, 
    0.0045367125996936628, 0.0043017363119994094, 0.0040481958090295483, 
    0.0037880958001854249, 0.0035326907292925268, 0.0032917993980226667, 
    0.0030732431093130255, 0.0028824538296510966, 0.0027222865596153406, 
    0.002593030143392413, 0.0024926034080009901, 0.0024169105442176167, 
    0.0023603054213539852, 0.0023161168863874352, 0.0022771838682478433, 
    0.0022363707690538333, 0.0021869898842470782, 0.0021231533689937106, 
    0.0020400093364814388, 0.0019338744862281518, 0.001802293587529234, 
    0.001644022350768735, 0.0014589677929042995, 0.0012480977199725344, 
    0.0010133329496970918, 0.00075741619152628952, 0.00048377740117665127, 
    0.00019638158900465947, -0.00010042053450429178, -0.00040204071302650936, 
    -0.00070382263883817387, -0.0010011744765045562, -0.001289744471021358, 
    -0.0015655601487449477, -0.0018252044273909165, -0.0020659712167542623, 
    -0.0022860248426221238, -0.0024845251810026903, -0.0026617165127885375, 
    -0.0028189469744723749, -0.0029586118205727754, -0.0030840080437000731, 
    -0.0031990664393172653, -0.0033079862435736987, -0.0034147565237323419, 
    -0.0035226403921584707, -0.0036336656740620604, -0.0037482219113662207, 
    -0.0038648197072846005, -0.0039800701531989861, -0.0040888887115679354, 
    -0.0041849185333455467, -0.0042611042910512551, -0.0043103663442711979, 
    -0.0043262861633334227, -0.0043037638039803748, -0.0042395281997062292, 
    -0.0041325177591693442, -0.0039840475975380912, -0.0037977854976093514, 
    -0.0035795171536443272, -0.0033367332333044185, -0.0030780748192794369, 
    -0.0028126865603863927, -0.0025495393845787568, -0.0022967696055826306, 
    -0.0020611161983495386, -0.0018474720911454113, -0.0016586221908391355, 
    -0.0014951689197062943, -0.0013556538144019637, -0.0012368523642282401, 
    -0.0011342256122605292, -0.001042456463719873, -0.00095603533382171662, 
    -0.00086983583836891391, -0.00077963396466269354, 
    -0.00068252886852053713, -0.0005772253502545232, -0.00046420519665330148, 
    -0.00034570066112384556, -0.00022553859033725348, 
    -0.00010881386238192504, -1.4428708797492329e-06, 9.0361453699249662e-05, 
    0.00016062058393499559, 0.00020408554444759612, 0.00021663248176766677, 
    0.00019554583209687208, 0.00013963784418574059, 4.9247340258296241e-05, 
    -7.3865978570694147e-05, -0.0002266985708986349, -0.00040521192327831485, 
    -0.00060457389342096824, -0.0008193936436817589, -0.0010439692092080437, 
    -0.001272491456229852, -0.0014992296822971759, -0.0017186779059728441, 
    -0.001925663848071771, -0.0021154469900256626, -0.0022838191712871692, 
    -0.0024272052659884053, -0.0025428035937844701, -0.0026287247986683361, 
    -0.0026841286572256194, -0.002709354832889279, -0.0027059913772939149, 
    -0.0026768749314551232, -0.0026259819075571391, -0.0025582129453202503, 
    -0.0024790737758473491, -0.002394264954175847, -0.0023092592801478712, 
    -0.002228883996522713, -0.0021569974438393202, -0.0020962879247283014, 
    -0.0020482101185012721, -0.0020130498980694767, -0.0019900855302081143, 
    -0.0019777921674540306, -0.001974039266832909, -0.0019762742598893619, 
    -0.0019816724860684462, -0.0019872658890047047, -0.001990095102249323, 
    -0.0019873809497849173, -0.0019767340427323046, -0.0019563824646525634, 
    -0.0019254079297378443, -0.0018839375099170103, -0.001833286608840697, 
    -0.0017759703459148055, -0.0017156277129159077, -0.001656790970754693, 
    -0.0016045312545117469, -0.0015639711392139996, -0.0015397091954773498, 
    -0.0015352403898451386, -0.0015524448940999187, -0.0015912724156998692, 
    -0.0016496423321487287, -0.001723581349682579, -0.0018075387833723249, 
    -0.0018948500677006654, -0.0019782611332820597, -0.0020504609068586511, 
    -0.0021045233023539319, -0.0021342554090934087, -0.0021343923388346714, 
    -0.0021006769321037983, -0.0020298571775437878, -0.0019196581086905005, 
    -0.0017687636688206109, -0.0015768321013429577, -0.0013445135221998806, 
    -0.001073520923651471, -0.00076668898221094004, -0.00042803615869081019, 
    -6.2791336696863291e-05, 0.00032264354669986307, 0.00072080990754679573, 
    0.0011234088678699111, 0.0015215922917927941, 0.0019063413814287037, 
    0.0022688877248180977, 0.0026011505503048728, 0.0028961412442217774, 
    0.003148296564506397, 0.0033537080983427219, 0.0035102249001520559, 
    0.0036174246081549701, 0.003676461920809363, 0.0036898328804455651, 
    0.003661101654537684, 0.0035946080871753208, 0.0034952115222427037, 
    0.0033680709322033413, 0.0032185061625707913, 0.0030518938244204494, 
    0.0028736290255162726, 0.0026891097642101972, 0.0025037148117448334, 
    0.0023227630153393355, 0.0021514026662957254, 0.0019944475377821915, 
    0.0018561492939029095, 0.0017399520909701636, 0.0016482809604291908, 
    0.0015824178738238425, 0.0015424856158192347, 0.0015275314430567338, 
    0.0015356715870064048, 0.0015642446548487, 0.0016099479766712021, 
    0.0016689698507054208, 0.0017371147004368443, 0.0018099730918395421, 
    0.0018831092095299654, 0.0019522924309274214, 0.0020137117683050243, 
    0.0020641608974472335, 0.0021011611720927899, 0.0021230194951933883, 
    0.0021288171306405299, 0.0021183455141866284, 0.0020919884760596868, 
    0.0020505729627211746, 0.0019951853234630966, 0.0019269952923350975, 
    0.0018470931614689603, 0.0017563549533357249, 0.0016553996277833543, 
    0.0015445922452830599, 0.0014241410448528247, 0.0012942073644463085, 
    0.0011550709149363118, 0.0010072758742260721, 0.0008517561214741304, 
    0.00068993590973897895, 0.00052375229256496644, 0.00035564514158533338, 
    0.00018848561682079877, 2.5469387022319001e-05, -0.00013000991859237875, 
    -0.00027446565715309268, -0.00040444421718290079, 
    -0.00051661715761177436, -0.00060786189735502494, 
    -0.00067535146845534378, -0.00071665090417495929, 
    -0.00072981648536204775, -0.00071353267656491261, 
    -0.00066725640181921741, -0.00059140369507134499, 
    -0.00048752235133824701, -0.0003584597772025632, -0.00020845398006655381, 
    -4.3121455944497621e-05, 0.00013070505050820857, 0.00030529203836446523, 
    0.0004724662933682642, 0.00062419752085617031, 0.00075321649822325488, 
    0.00085363689795923937, 0.0009214739018122165, 0.00095503220885081942, 
    0.00095509362340258689, 0.0009248837961200922, 0.00086982052779751488, 
    0.00079704621621288271, 0.00071482078973373274, 0.000631784088452201, 
    0.00055619875359210337, 0.00049521004306133873, 0.00045417820807008472, 
    0.00043615602757190872, 0.00044153196034522934, 0.00046786666666459998, 
    0.00050997467773547718, 0.00056022535207307341, 0.00060904557548764984, 
    0.00064561509030552444, 0.00065866365930531334, 0.00063732703970898429, 
    0.0005719847159442841, 0.00045502838281737189, 0.0002815228672933994, 
    4.9691697497596717e-05, -0.00023879270588176801, -0.00057872737868218654, 
    -0.00096154710394187766, -0.0013757544720509527, -0.001807567740642531, 
    -0.0022417931713953516, -0.0026628226070573606, -0.0030556411099475567, 
    -0.0034067562563533356, -0.0037049286324563001, -0.0039417175106223629, 
    -0.0041117669620531335, -0.0042128970934252295, -0.0042460065452277901, 
    -0.0042147938153815042, -0.0041253386758342819, -0.0039855800458408613, 
    -0.0038047160061323577, -0.003592595739064688, -0.0033591525665010026, 
    -0.0031139210377943861, -0.0028656773711385618, -0.0026221502857165071, 
    -0.002389850223454578, -0.0021739247674749723, -0.0019780503099142287, 
    -0.0018043798163408225, -0.0016535172257394024, -0.0015245573695925525, 
    -0.0014151577055342612, -0.0013216751914682794, -0.0012393650065239295, 
    -0.0011627112000975816, -0.0010858485825043908, -0.0010030568863686944, 
    -0.0009092214369397513, -0.0008002359207547403, -0.0006732545991345758, 
    -0.0005268609419369697, -0.00036112663956641689, -0.00017760502768881701, 
    2.0719136494911879e-05, 0.00022956238092324401, 0.00044352239496580823, 
    0.0006563305708731298, 0.00086119122926959363, 0.0010511221901147554, 
    0.0012193166390639179, 0.0013594932838514103, 0.001466213973361477, 
    0.0015351860493183715, 0.0015635126601058202, 0.0015498986551306191, 
    0.0014947813346993229, 0.0014003992056172334, 0.0012707635507121784, 
    0.0011115243476759367, 0.00092973024541267958, 0.00073348234170282048, 
    0.00053151267830349263, 0.00033271150300899445, 0.00014565204855641564, 
    -2.1861073496563408e-05, -0.00016320503935911214, 
    -0.00027327086585644838, -0.00034869319931621801, 
    -0.00038796891631723664, -0.00039139239005324714, 
    -0.00036086389020067663, -0.00029954140604706431, 
    -0.00021140681632451894, -0.00010079847228041473, 2.802028415965107e-05, 
    0.00017119904659265489, 0.00032551587769582044, 0.00048847554813579721, 
    0.00065827002908034173, 0.0008336744362909365, 0.0010138682864853459, 
    0.0011982067332497808, 0.0013860155445448654, 0.0015763804341821686, 
    0.001767980756746706, 0.0019589799513943249, 0.0021470020408719381, 
    0.0023291979486452044, 0.0025024097714916051, 0.0026633978454869756, 
    0.0028091447664761304, 0.0029371498603340727, 0.0030457259856638032, 
    0.0031342143084896286, 0.0032031041014619053, 0.0032540610350329088, 
    0.003289800270470997, 0.003313884733850411, 0.0033304398024508134, 
    0.0033437972338155506, 0.0033581210778558077, 0.0033769891247506828, 
    0.0034029727399525651, 0.0034371884951958994, 0.0034789131502157584, 
    0.0035253346726437135, 0.0035715840450376954, 0.0036111378035848262, 
    0.003636602966154606, 0.0036407436333040603, 0.0036175222705530858, 
    0.0035628977748538037, 0.0034752356181940113, 0.0033552927215526316, 
    0.0032059319360729808, 0.0030317318349677783, 0.0028385249358573528, 
    0.0026329889964504961, 0.002422301322298836, 0.0022137941987768555, 
    0.0020147039363589995, 0.0018319111148853262, 0.001671731299467243, 
    0.0015397168549705731, 0.0014404513778872841, 0.0013773763994658177, 
    0.0013526103699028913, 0.0013668079533747358, 0.0014190049335903493, 
    0.0015065524357602243, 0.0016250914858359986, 0.0017686350335374649, 
    0.0019297432886445373, 0.0020997929954581639, 0.0022693545823279349, 
    0.0024286282078465954, 0.0025679410606725167, 0.0026782359950251254, 
    0.0027515714983105304, 0.0027815311993401107, 0.0027635305678551637, 
    0.0026949543394955713, 0.0025751347169652022, 0.0024051581452435369, 
    0.0021875405343086485, 0.0019258385044716884, 0.0016242479837934888, 
    0.0012872290701060882, 0.00091923395806644019, 0.00052451218074141303, 
    0.00010698619867289833, -0.00032975003894334829, -0.00078237087626025165, 
    -0.0012477055935299192, -0.0017225698849892696, -0.0022036110875512699, 
    -0.0026871498427592888, -0.0031691189015878125, -0.0036450686533954098, 
    -0.004110259120185724, -0.0045598363376144141, -0.0049890880485250443, 
    -0.0053937136678499573, -0.0057700534285265205, -0.006115245762753266, 
    -0.0064272320975350501, -0.0067046263423373477, -0.0069464606816269907, 
    -0.0071518886753937708, -0.0073198892781724794, -0.0074490485756149097, 
    -0.0075375187201547986, -0.0075831303971431582, -0.0075836259532091983, 
    -0.0075369261207668863, -0.0074413287783939731, -0.00729567091257231, 
    -0.0070994790105419047, -0.0068531266073552193, -0.0065579593633484853, 
    -0.0062163461296703771, -0.0058315774131601113, -0.0054076220865052968, 
    -0.0049487944521043065, -0.0044593745362113196, -0.0039434035206570963, 
    -0.0034046011331787516, -0.002846530883481576, -0.0022729540395096297, 
    -0.0016882696024519452, -0.0010978818003777981, -0.00050838972510574502, 
    7.2480311179590651e-05, 0.00063624955569517594, 0.0011742880423332839, 
    0.0016784948779906431, 0.0021419607077821576, 0.0025594734944848646, 
    0.0029277875292926152, 0.0032456785041420607, 0.003513777844683826, 
    0.003734247970204589, 0.0039103586755490638, 0.0040460004081748976, 
    0.0041451825841624362, 0.0042115468055167332, 0.0042479482378856293, 
    0.0042561966945029173, 0.0042368787320742592, 0.0041893559387107997, 
    0.004111899331635996, 0.0040019746890474807, 0.0038565980830819156, 
    0.0036728516240759493, 0.0034483414188324073, 0.0031816782758786119, 
    0.0028728464413051583, 0.0025234993798633433, 0.0021370986725049237, 
    0.0017189786818050832, 0.00127626466558889, 0.00081768323544335257, 
    0.0003532538055153868, -0.00010615709274417693, -0.00054936472737981295, 
    -0.00096550182999535013, -0.0013446783415244719, -0.00167862863942683, 
    -0.001961268097957485, -0.0021890894566797179, -0.0023613459467859122, 
    -0.0024800437075670743, -0.0025496682916027317, -0.0025767455940266274, 
    -0.0025692741516463238, -0.0025361042279406333, -0.0024863023244201705, 
    -0.0024286523328362125, -0.0023711970471148695, -0.0023209730653095447, 
    -0.0022838254972879692, -0.0022643721139206951, -0.0022660205639748725, 
    -0.0022910363347925962, -0.002340657501041293, -0.0024152297572165608, 
    -0.00251433933020673, -0.0026370095364351806, -0.0027819055719524861, 
    -0.0029475594755880834, -0.0031325953648108193, -0.0033358736490275379, 
    -0.00355656038875492, -0.0037940772257122682, -0.0040478999542605427, 
    -0.0043173182051231464, -0.0046011688496182144, -0.004897574456873964, 
    -0.0052037946777653615, -0.0055161460436070689, -0.0058300897647701778, 
    -0.006140405173515817, -0.0064415279371206032, -0.0067278987565423552, 
    -0.0069943166690905638, -0.0072362433569000103, -0.0074500468792626975, 
    -0.0076331894715065424, -0.0077843595738726484, -0.0079035338995436417, 
    -0.0079919376815215624, -0.0080519273696356853, -0.0080867825797494054, 
    -0.0081003730243163902, -0.0080968169213981693, -0.0080800512653183068, 
    -0.0080534271560171126, -0.0080193183632209439, -0.0079787656127901004, 
    -0.0079312562272866108, -0.0078745843119769187, -0.0078048966526845058, 
    -0.0077168866145803016, -0.0076042412944940449, -0.00746014471324144, 
    -0.0072779606551959383, -0.0070519360653014899, -0.0067778711978287156, 
    -0.0064537056230235985, -0.0060799162560257591, -0.0056597317495533823, 
    -0.0051990911827024073, -0.0047063816066584309, -0.0041919763934621769, 
    -0.0036675601940694934, -0.0031453513365280344, -0.0026372605812407038, 
    -0.0021540726659772134, -0.0017047839820701989, -0.0012961976897569473, 
    -0.00093272080865103714, -0.00061651819795103288, 
    -0.00034784721347596984, -0.00012551301130993395, 5.2631544676971309e-05, 
    0.00018929853014218586, 0.0002874746870754636, 0.00035027397422802812, 
    0.00038092381743332364, 0.00038285432782623113, 0.00035985725360482306, 
    0.00031622674700921736, 0.00025695404262231247, 0.00018786149116376932, 
    0.00011567247803886136, 4.797920708447985e-05, -6.9338851152497393e-06, 
    -4.0408894708143534e-05, -4.3891126673253813e-05, -9.534193600990986e-06, 
    6.9174191353929418e-05, 0.00019676676987783587, 0.00037526659254753878, 
    0.00060382888257349936, 0.00087857565209676898, 0.0011927149233918377, 
    0.0015368354867141688, 0.0018994268288314727, 0.0022675273490529385, 
    0.0026274360251862298, 0.0029655088525209032, 0.0032688620282676018, 
    0.0035260961231683282, 0.0037278559822210592, 0.0038672792396744725, 
    0.0039402678937819936, 0.003945575912593596, 0.0038847293574748466, 
    0.0037617655439581088, 0.0035828907724225734, 0.0033560272909485857, 
    0.0030903356851555187, 0.0027957098784791826, 0.0024822830122726326, 
    0.0021599610204364734, 0.0018380022978519842, 0.0015247078540820882, 
    0.0012271552271844127, 0.00095113725675908026, 0.00070119946391765452, 
    0.00048079911119436694, 0.00029262333826612008, 0.00013885777450019351, 
    2.1535341259415301e-05, -5.7236394029027294e-05, -9.51292024660229e-05, 
    -8.965602943249119e-05, -3.8317185340816648e-05, 6.1028964232775302e-05, 
    0.00020973290731072136, 0.00040783205262996647, 0.00065355761445401407, 
    0.00094301175699665774, 0.0012699738234800328, 0.0016258716145148928, 
    0.0019999469679230879, 0.0023795975256275135, 0.0027507782773844242, 
    0.0030985688232405065, 0.0034077957294817657, 0.0036637655624267313, 
    0.0038530420467554429, 0.0039642693332897451, 0.0039888556903150008, 
    0.0039215372348123407, 0.0037606588395393478, 0.0035082971870847813, 
    0.0031701122153123852, 0.0027549758145455914, 0.0022743716740386642, 
    0.0017416914373824229, 0.0011712985526375606, 0.00057759583221617746, 
    -2.5896592315973258e-05, -0.0006272748728446268, -0.0012167782014274129, 
    -0.0017869832686598171, -0.0023327579791931979, -0.0028509965632410135, 
    -0.0033401750618070603, -0.0037998292482437435, -0.0042299568923906735, 
    -0.0046305532259523713, -0.005001282036501787, -0.0053415284142843376, 
    -0.0056508905265575948, -0.0059299810782457588, -0.0061810306873953114, 
    -0.0064079312601453831, -0.0066156011509064918, -0.0068090096783556715, 
    -0.0069922629065403774, -0.0071681424267640223, -0.0073379987282716566, 
    -0.0075019298540377815, -0.0076591524943432398, -0.0078083188736766109, 
    -0.0079478668864725009, -0.0080762185130928144, -0.0081919614917590009, 
    -0.0082940085015786886, -0.0083816782424931558, -0.0084548030309815735, 
    -0.0085138023683239451, -0.0085598197216000486, -0.0085948698213392984, 
    -0.0086220796338446724, -0.0086458006714753913, -0.0086715700757847829, 
    -0.0087057881417626198, -0.008755031357600038, -0.0088251578873323085, 
    -0.0089202553902827421, -0.009041724513961874, -0.0091875082616334636, 
    -0.0093518703369004745, -0.0095256013609727446, -0.009696827840283858, 
    -0.0098522057414680859, -0.009978439563205866, -0.010063828510405687, 
    -0.010099566933316649, -0.010080702479303609, -0.010006453704908, 
    -0.009880094646316704, -0.0097083775514588272, -0.0095007339159365409, 
    -0.0092682507962710513, -0.0090227406200621592, -0.0087756545762329337, 
    -0.0085371542399110406, -0.0083151633717536734, -0.008114691406429406, 
    -0.0079374869240116993, -0.0077819855976075381, -0.00764372051470554, 
    -0.0075158518916015275, -0.0073899877400807421, -0.0072570072797316131, 
    -0.0071081462476822871, -0.0069359039657088586, -0.0067350567000722446, 
    -0.0065035150686866428, -0.006242852976573475, -0.005958594305247868, 
    -0.0056600590888630578, -0.0053599115320824876, -0.0050733895082288021, 
    -0.0048174142236867869, -0.0046096316886629291, -0.0044674731639603917, 
    -0.0044073285659677747, -0.0044438586227746714, -0.0045893617800823946, 
    -0.0048531505270352935, -0.0052410888540350828, -0.0057550818481848613, 
    -0.0063927939850656462, -0.0071476209547979598, -0.0080088175143943983, 
    -0.0089619937968950132, -0.0099897436388933815, -0.011072401427138783, 
    -0.012188701609562348, -0.013316522056874596, -0.014433432759218507, 
    -0.015517437078786103, -0.016547865644892912, -0.017506266186224733, 
    -0.018377453176014608, -0.019150276288271102, -0.019818211218333666, 
    -0.020379709201794282, -0.02083809510280971, -0.021201318421605154, 
    -0.021481212511267542, -0.021692578812614379, -0.021851865920279039, 
    -0.021975542927843289, -0.022078435683907854, -0.022172128681068014, 
    -0.022263597375968922, -0.022354508773659552, -0.022441328720494536, 
    -0.022516244578106543, -0.022568933214471509, -0.022588740953870368, 
    -0.022566783583699547, -0.022497296966630092, -0.022378181284097354, 
    -0.022210756943085101, -0.021999027663466522, -0.021748866637554768, 
    -0.021467370425274617, -0.021162375240528934, -0.02084248790096048, 
    -0.020517173575890432, -0.020197198956135282, -0.019894874709617226, 
    -0.019623884645220475, -0.019398881856808159, -0.019234443836667125, 
    -0.019143550424138626, -0.019135988463222849, -0.019216423360112426, 
    -0.019382943038944028, -0.019625851332599156, -0.019927065990185944, 
    -0.02026042107322195, -0.020592337267704239, -0.020883400858204282, 
    -0.021090155649029534, -0.021167563615034583, -0.021071429131471562, 
    -0.020761387398734871, -0.020203629995558702, -0.019373836315335714, 
    -0.018259784835948707, -0.016863151381948716, -0.015200226368960823, 
    -0.013301006719115308, -0.011207138017706777, -0.0089685241096347131, 
    -0.0066397540349104264, -0.0042764253424455983, -0.0019318815776843742, 
    0.00034593119194151363, 0.0025166983002619095, 0.0045506668477820564, 
    0.0064298061159288869, 0.0081482262626489665, 0.009710342033727698, 
    0.011127271095542483, 0.01241161308417366, 0.013571809132688689, 
    0.014607505243712631, 0.015506483256396924, 0.016244458731769714, 
    0.016787342421815996, 0.017095793217048204, 0.017130812557909044, 
    0.016859777542705782, 0.016260980534396341, 0.015326392212354366, 
    0.014062085951894857, 0.012487318350881908, 0.010631915536137822, 
    0.0085334093148129592, 0.0062340390873036394, 0.0037788494882908677, 
    0.0012135927341574513, -0.0014165591035159291,
  // Fqt-Na(8, 0-1999)
    1, 0.99221783324621937, 0.96927742686805929, 0.93235650495169542, 
    0.88329282331829662, 0.82441723834983116, 0.75835397107509095, 
    0.68781375605388506, 0.61540357844435967, 0.54347133085725863, 
    0.47399633141534697, 0.40852887059871551, 0.34817535686433759, 
    0.29362089881784204, 0.24517862092718026, 0.20285470286379548, 
    0.16641919906276256, 0.13547490780175467, 0.10951897254689129, 
    0.087994383653861946, 0.070330344239891596, 0.055971958930212888, 
    0.044400478871448081, 0.035145701722665866, 0.027792234583777845, 
    0.02198113611669026, 0.017408302318662364, 0.013820702802576419, 
    0.011011336648282249, 0.0088135584137464563, 0.0070952057602476576, 
    0.0057528363596886139, 0.0047063160917559894, 0.0038938813204592109, 
    0.0032678283008879916, 0.0027908989857895815, 0.0024334214318172138, 
    0.0021711684039492714, 0.0019838657256748987, 0.0018542359049075661, 
    0.0017674140456942122, 0.0017106165981640453, 0.0016729136485195673, 
    0.0016450660258217108, 0.0016193486447245548, 0.0015893818855485138, 
    0.0015499621378757813, 0.0014969130248527651, 0.0014269545048872876, 
    0.0013375926139952278, 0.0012270355575359575, 0.0010941532952160539, 
    0.00093846400880889715, 0.00076016230460951035, 0.00056017522148660488, 
    0.00034021535544694092, 0.00010283172449516319, -0.00014858512024301443, 
    -0.00040985796191904595, -0.00067612421299820063, 
    -0.00094200926112476672, -0.0012018526617464068, -0.0014499876207561308, 
    -0.0016810624908045369, -0.0018904039138780988, -0.0020743757254786041, 
    -0.0022307025810685776, -0.0023586693570319811, -0.0024591584925110644, 
    -0.0025345066470636251, -0.002588215770174125, -0.0026245780008125499, 
    -0.0026482717936203337, -0.0026639407410604375, -0.0026757904152368175, 
    -0.0026871867221443836, -0.0027002972957139207, -0.0027157958156620895, 
    -0.0027326896997503982, -0.0027483055101367171, -0.0027584686942609938, 
    -0.0027578711174803369, -0.0027405828143137862, -0.0027006498875831054, 
    -0.002632696852062578, -0.0025324380406607293, -0.0023970322347716092, 
    -0.0022252349744645255, -0.0020173595478273506, -0.0017750626204039107, 
    -0.0015010623759548684, -0.0011988486847644021, -0.00087245189216646082, 
    -0.00052631197029708553, -0.00016522439818087971, 0.00020565000240503091, 
    0.00058075334312323625, 0.00095411201703094687, 0.0013193482101060724, 
    0.0016697523417776195, 0.0019984271000337791, 0.0022984888503448479, 
    0.0025633309948635873, 0.0027869054926267412, 0.0029640214786935863, 
    0.0030906201802465691, 0.0031640378317254413, 0.0031832342234434626, 
    0.0031489977368274915, 0.0030640874294519862, 0.0029333123901890174, 
    0.002763496165372979, 0.0025632967500939657, 0.0023428738312212902, 
    0.0021133835835567749, 0.0018863495251341285, 0.0016729557882637488, 
    0.0014833509787062359, 0.0013260486115240983, 0.0012074924703897184, 
    0.0011318207138496495, 0.0011008307141366102, 0.001114130283379414, 
    0.0011694091598220603, 0.0012627793714136881, 0.0013891179237204465, 
    0.0015423831394376045, 0.0017158778487067151, 0.001902486852624225, 
    0.0020949046045628272, 0.0022858822596140294, 0.0024684976370456281, 
    0.0026364267462115668, 0.0027841864009730973, 0.0029073105425342512, 
    0.0030024352869798352, 0.0030672771239707119, 0.0031005328274155502, 
    0.0031017089204814223, 0.0030709328421283013, 0.0030087914904804625, 
    0.0029162181509713872, 0.0027944791336783552, 0.0026452504606112363, 
    0.0024707828734168449, 0.0022740973673873624, 0.0020591889301833487, 
    0.0018311541947882348, 0.0015962068605343662, 0.0013615345240036594, 
    0.0011349644284545807, 0.00092447177196028092, 0.00073755286315970077, 
    0.00058054504419681246, 0.00045799137226812836, 0.00037214293968223892, 
    0.00032269109884774342, 0.00030678852066099663, 0.00031937762596073401, 
    0.00035377174683590476, 0.00040240088771189078, 0.00045760589285826056, 
    0.00051233743634920121, 0.00056069328487249475, 0.00059825756334698759, 
    0.00062223422401861165, 0.00063144189719639579, 0.00062619911164304141, 
    0.00060815565812885304, 0.00058008239571551482, 0.00054562984799980628, 
    0.00050905228087398365, 0.00047488762232907202, 0.00044761755722661504, 
    0.00043132307687847944, 0.00042935721677649053, 0.00044406440955092939, 
    0.00047655854335029192, 0.00052659530088816566, 0.00059254385661371091, 
    0.00067146334898198238, 0.00075929534867199319, 0.00085114670706951958, 
    0.00094165515680322308, 0.0010254044436015521, 0.0010973576459567293, 
    0.0011532748133261245, 0.0011900927249934125, 0.0012062279604626285, 
    0.0012017878717753934, 0.0011786432178793502, 0.0011403603868016267, 
    0.0010919615308981996, 0.0010395260944082688, 0.000989663028277774, 
    0.00094890503765627512, 0.00092311446128665823, 0.0009169701764816261, 
    0.00093361013540413276, 0.00097446048768390922, 0.0010392765338492331, 
    0.0011263701905683471, 0.0012329617982055337, 0.0013556030725485916, 
    0.0014905919103468303, 0.0016343126816797029, 0.0017834643952507232, 
    0.0019351583035066996, 0.0020869018513019612, 0.0022365151953392644, 
    0.0023820128021102643, 0.0025215105926058813, 0.0026531881074766902, 
    0.0027753169527034633, 0.0028863457276149538, 0.002985021295638312, 
    0.0030705259363025491, 0.0031425812666575114, 0.0032015109564340377, 
    0.0032482208042818889, 0.0032841079520722774, 0.0033108743688494095, 
    0.0033302881904558831, 0.0033439032604949334, 0.0033528021720881747, 
    0.0033573803022327086, 0.0033572422732738648, 0.0033512028630418868, 
    0.003337410254287508, 0.0033135630354386471, 0.0032771826766911706, 
    0.0032259051827363194, 0.0031577382073126391, 0.0030712720882370478, 
    0.0029658256277671677, 0.0028415216542268785, 0.0026993161075628313, 
    0.0025409845211175515, 0.0023690785559611067, 0.0021868607218254806, 
    0.0019982130979444585, 0.0018075101804153931, 0.0016194376518833555, 
    0.0014387636569879263, 0.0012700488849253168, 0.0011173228736971554, 
    0.00098376482100536638, 0.000871407708120952, 0.00078091821285881805, 
    0.00071147972777158897, 0.00066081219029517739, 0.00062531876529376817, 
    0.00060037536126570919, 0.00058070997571315177, 0.00056083384398773165, 
    0.00053545202307540949, 0.00049981435891883184, 0.00044993808864357868, 
    0.00038272335350465319, 0.00029595894155417049, 0.00018827566088775046, 
    5.9086671919866016e-05, -9.1452622002595539e-05, -0.00026242369913379715, 
    -0.00045209264885573338, -0.00065781479186394274, 
    -0.00087595356095487614, -0.0011018452113822639, -0.0013298464877199608, 
    -0.001553507713456031, -0.0017658742960593335, -0.0019598937528944732, 
    -0.0021289128500976175, -0.002267195849542685, -0.0023704151378066847, 
    -0.0024360567992535516, -0.0024636855209907598, -0.0024550484438099662, 
    -0.0024139697744913705, -0.0023460544638274042, -0.0022582042112136796, 
    -0.0021580047056390475, -0.0020530365986127035, -0.0019502137460657135, 
    -0.0018552161507815852, -0.0017721020991571959, -0.0017031128913014856, 
    -0.0016487005238066837, -0.0016077248126475589, -0.0015777810495280738, 
    -0.0015555890270294657, -0.001537382955338363, -0.0015192563101587679, 
    -0.0014974283083899207, -0.0014684301008363854, -0.0014292126879203188, 
    -0.0013772006900383913, -0.001310309680961701, -0.0012269662820831237, 
    -0.0011261262297132561, -0.001007326928633456, -0.00087076808913020523, 
    -0.00071741347173169231, -0.00054910348333973077, 
    -0.00036864768203758369, -0.00017988394151782257, 1.2340931896057412e-05, 
    0.00020226694961611357, 0.00038343179967607438, 0.00054897922004774273, 
    0.0006920609946964735, 0.00080628738411474754, 0.00088617706264583376, 
    0.0009275318602720605, 0.00092768075739909533, 0.00088555544520096258, 
    0.00080160197542431672, 0.00067755462167579821, 0.00051614999370001077, 
    0.00032084418852908848, 9.5607362497466121e-05, -0.0001551789554182383, 
    -0.0004267375096956023, -0.00071386000091220149, -0.0010108553353476127, 
    -0.0013115435039562167, -0.0016092769948037313, -0.0018970084290634425, 
    -0.0021673920400941669, -0.0024129297828633474, -0.0026261904461307739, 
    -0.0028001192007456634, -0.0029284475497563306, -0.0030061811684273828, 
    -0.0030301044549487367, -0.0029992340177033166, -0.0029151388424119547, 
    -0.002782053916824778, -0.0026067477837222529, -0.0023981385006700429, 
    -0.0021666747043332054, -0.0019235612565768989, -0.001679907216550582, 
    -0.0014459288756108861, -0.0012302773180251215, -0.0010395926895841493, 
    -0.00087829093100951004, -0.0007485966521114611, -0.00065074408550752866, 
    -0.00058332178190160285, -0.00054366389458180295, 
    -0.00052825608258123499, -0.00053309791546691707, 
    -0.00055399569459695368, -0.00058676547280990966, 
    -0.00062735438540850751, -0.00067188830554461493, 
    -0.00071668300800406017, -0.00075824795998296625, 
    -0.00079329751831252321, -0.00081880378411935246, 
    -0.00083206966263079675, -0.00083083439133512383, 
    -0.00081337600458656636, -0.00077863906435043353, 
    -0.00072634879725652548, -0.00065712753382958533, 
    -0.00057259887034751531, -0.00047543492975401212, 
    -0.00036933307161073249, -0.00025887525900660543, 
    -0.00014926531872523109, -4.5941282667732021e-05, 4.5885342870312666e-05, 
    0.00012172125227330439, 0.00017824737544692629, 0.00021366614498180634, 
    0.00022791498581230626, 0.00022269994598496444, 0.00020135271646050883, 
    0.00016853181414135202, 0.00012980424932459045, 9.1152782652864227e-05, 
    5.8466329053799473e-05, 3.7060968427137257e-05, 3.1297768793784122e-05, 
    4.4299452574509367e-05, 7.7807113048646937e-05, 0.00013214792073975646, 
    0.00020632459232827004, 0.00029817754953854233, 0.00040459947142190608, 
    0.00052174329850152457, 0.00064520691910631433, 0.00077016502151339248, 
    0.00089146622992242609, 0.0010037171400769582, 0.001101382482198376, 
    0.001178917085154096, 0.0012309414840706041, 0.0012524470873715634, 
    0.0012390143571012736, 0.0011870284697259456, 0.0010938631000934076, 
    0.00095802529562448468, 0.00077924243393598771, 0.00055850056652203704, 
    0.00029803163277992246, 1.2450584673118084e-06, -0.00032735305154932856, 
    -0.00068226146466412031, -0.0010570983538717351, -0.0014447072198040659, 
    -0.0018372902066322852, -0.0022265566327925425, -0.0026039221149554512, 
    -0.0029607435959781332, -0.0032886007094338207, -0.0035796120182287968, 
    -0.003826794009600626, -0.0040244222264230294, -0.0041683800657932833, 
    -0.0042564377157335975, -0.0042884148845334438, -0.0042662045230279335, 
    -0.0041936418273212624, -0.0040762658567682413, -0.0039209871609923912, 
    -0.0037357091740948256, -0.0035289328393434422, -0.0033093639094900484, 
    -0.0030855494838032765, -0.002865554403559263, -0.0026566512018670616, 
    -0.002465031968842952, -0.0022955194699204574, -0.0021513024959379009, 
    -0.0020337367229940418, -0.0019422643526083394, -0.0018744932997422647, 
    -0.0018264523781051246, -0.0017930107466118646, -0.0017683897022047553, 
    -0.0017467079345290784, -0.0017224982126653899, -0.0016911454920975203, 
    -0.0016492190868024142, -0.0015946974342424466, -0.001527073419425391, 
    -0.0014473385027909103, -0.0013578644739446039, -0.0012621935551612859, 
    -0.0011647523586582058, -0.0010705453371590346, -0.00098483769716007242, 
    -0.00091285023483311345, -0.00085948416718416212, 
    -0.00082908249579758851, -0.00082523870494125408, 
    -0.00085066115297216332, -0.00090706971070516219, 
    -0.00099511881890514261, -0.0011143118351837917, -0.0012629278558813084, 
    -0.0014379529427331963, -0.0016350562074458157, -0.0018486367273475746, 
    -0.0020719518987106543, -0.0022973513946106016, -0.002516592221631832, 
    -0.002721240534684631, -0.0029031264354345671, -0.0030548393995908849, 
    -0.0031702145687682909, -0.0032447661714477133, -0.0032760308367064893, 
    -0.0032637586567571069, -0.0032099214049635429, -0.0031185135419741538, 
    -0.0029951563866775352, -0.0028465304812391378, -0.002679713227815832, 
    -0.0025015010348167274, -0.0023178020802228408, -0.0021331937204396786, 
    -0.0019506829879373691, -0.0017716851839040873, -0.0015962115545889591, 
    -0.0014232256768988516, -0.0012510753096266378, -0.0010779800215135798, 
    -0.00090245216565478089, -0.00072363298638025871, -0.0005414570473382213, 
    -0.00035665152827942036, -0.00017056217043891743, 1.5139717000747002e-05, 
    0.00019876713077650744, 0.00037888779595690109, 0.00055445180148088239, 
    0.00072476728721747015, 0.00088934004652173576, 0.00104760305922616, 
    0.0011986475604569505, 0.0013410061868203657, 0.0014725756568776962, 
    0.001590677950801101, 0.0016922624104294022, 0.0017741972904285318, 
    0.0018336114855217454, 0.0018682572764999899, 0.0018768578737764765, 
    0.0018594042911597836, 0.0018173725817849139, 0.0017537940171541912, 
    0.0016731457857262241, 0.001581045744762448, 0.0014837618747900766, 
    0.0013876069024235699, 0.0012982870663017022, 0.0012203070251089537, 
    0.0011564853820983548, 0.0011076725743490753, 0.0010726860413872738, 
    0.0010484770335194467, 0.0010305144566402833, 0.0010133325351235965, 
    0.00099118050184122237, 0.00095869829622403945, 0.00091155064673457574, 
    0.00084694292119228288, 0.00076398274616639383, 0.00066383447479779621, 
    0.00054965328100749038, 0.00042628450037832767, 0.00029978335393644078, 
    0.00017678032728516747, 6.3796359366250215e-05, -3.3415927202665928e-05, 
    -0.0001104047136437512, -0.00016435423755656976, -0.0001942053327353089, 
    -0.00020057386425596156, -0.00018552603976081035, 
    -0.00015226648058284665, -0.00010479935993436891, 
    -4.7606148118719172e-05, 1.4621199889006098e-05, 7.7206616638849702e-05, 
    0.00013564296923831813, 0.00018572450432639435, 0.00022366220981518618, 
    0.00024623647836382424, 0.0002509856272564278, 0.00023645664165903885, 
    0.00020245599215619296, 0.00015027283146699558, 8.2812546711670976e-05, 
    4.5984384329219924e-06, -7.8398930196682298e-05, -0.00015908875384443202, 
    -0.00022974511128911091, -0.00028260343473843783, 
    -0.00031053438665489105, -0.00030772924280349028, 
    -0.00027033073889314854, -0.00019693615866375497, 
    -8.8905999992834215e-05, 4.9563484423023152e-05, 0.00021163516220139929, 
    0.00038828964235325717, 0.00056901443239741958, 0.00074266934217229338, 
    0.00089841418520209416, 0.0010266421739767041, 0.0011197641377259559, 
    0.0011727995331661802, 0.0011836773741002206, 0.0011532574630188802, 
    0.0010850643920016852, 0.0009848124798494081, 0.00085977140623632947, 
    0.00071806107882723704, 0.00056795829980573202, 0.00041726620723317443, 
    0.00027279389566367361, 0.00013998199299235009, 2.2701858032897417e-05, 
    -7.6779488465701065e-05, -0.00015768168393732334, 
    -0.00022045433665406479, -0.00026643807781354936, 
    -0.00029747380385416176, -0.00031551873943780345, 
    -0.00032231267954006045, -0.00031914198505123193, 
    -0.00030671739940139501, -0.00028518401372562108, 
    -0.00025423810014608858, -0.00021335095916809695, -0.0001620072934352099, 
    -9.9948696026471335e-05, -2.7375383830753939e-05, 5.4914707183706298e-05, 
    0.00014544607478716437, 0.0002420247667656652, 0.00034173974964781976, 
    0.00044098408246849683, 0.00053551307722109578, 0.00062052572473488845, 
    0.00069082136332147652, 0.00074101727964883464, 0.00076583875925078087, 
    0.000760489878214978, 0.00072108088368613048, 0.00064506332476744262, 
    0.0005316189079354809, 0.00038194492108668929, 0.00019936859967621069, 
    -1.0750760780041738e-05, -0.00024132052742664538, 
    -0.00048399475152027669, -0.00072976402710932318, 
    -0.00096958622751718839, -0.0011949841449546993, -0.001398561451489084, 
    -0.0015743827303958831, -0.0017182319785168936, -0.0018277365472871268, 
    -0.0019023669538456296, -0.0019433269870269285, -0.001953332141844745, 
    -0.0019362830476290513, -0.0018968718332968565, -0.0018401331496329279, 
    -0.0017709819367023433, -0.0016937824156127582, -0.0016119700070317215, 
    -0.0015277938863200423, -0.0014422027509968882, -0.001354924008473896, 
    -0.0012647144259861612, -0.0011697795690299552, -0.0010682512572742899, 
    -0.00095868717530377232, -0.00084046818475169455, 
    -0.00071407614111138713, -0.00058119658770452239, 
    -0.00044468075748605135, -0.00030836848076832906, 
    -0.00017680307016281112, -5.4870240257836658e-05, 5.2611053569970239e-05, 
    0.00014132111640438751, 0.00020787067750515712, 0.00025018004396308856, 
    0.00026778461163092204, 0.00026200488698041542, 0.00023598355333463697, 
    0.00019453734824576306, 0.0001438490138471043, 9.1015400662687742e-05, 
    4.346498248763685e-05, 8.3383224101426243e-06, -8.1381586063973663e-06, 
    -1.192058301586823e-06, 3.2083472354538375e-05, 9.2501056067702389e-05, 
    0.00017874420836569671, 0.00028754040517262909, 0.00041398404456193585, 
    0.0005519935215390283, 0.00069482112971042511, 0.00083556781846621912, 
    0.00096766670453884453, 0.001085289482891964, 0.0011836670156517874, 
    0.0012593109198982609, 0.0013101363655386631, 0.0013354996570432748, 
    0.0013361625231021342, 0.0013141820739488953, 0.0012727144568336042, 
    0.0012157422699396664, 0.0011477086448864727, 0.0010731159005183976, 
    0.00099612991123335559, 0.00092024294526459158, 0.00084804726591267935, 
    0.00078112432427525271, 0.00072002271895024663, 0.00066433734573373231, 
    0.0006128240600173807, 0.00056355489955391982, 0.0005140915944116468, 
    0.00046164419861197917, 0.00040322608248534903, 0.00033581489232875362, 
    0.00025653011172822469, 0.00016283143452793745, 5.2747493203671387e-05, 
    -7.4879694005597591e-05, -0.00022014852173456048, 
    -0.00038190868653105328, -0.00055764048503995902, 
    -0.00074348256238198729, -0.00093441887082770813, -0.0011246378241821407, 
    -0.0013080456961837095, -0.0014788754454232876, -0.0016322993021433072, 
    -0.0017649565855427452, -0.0018752764744767046, -0.0019635482469778638, 
    -0.0020316982252425019, -0.0020828141102814586, -0.0021205028195129165, 
    -0.0021481907555342046, -0.0021684792573528492, -0.0021826470937689633, 
    -0.0021903846806323821, -0.0021897669789967648, -0.0021774618069531878, 
    -0.0021491528065575105, -0.0021000951949025027, -0.0020257498946194873, 
    -0.0019224127985104341, -0.0017877985419436314, -0.0016214999490734652, 
    -0.0014253154794226174, -0.0012033699091110145, -0.00096205062548079725, 
    -0.00070968383097713716, -0.00045600209491084584, 
    -0.00021141168735606703, 1.3849709827176308e-05, 0.00021056687916503022, 
    0.00037131616888334042, 0.00049106762607182696, 0.00056754029952635397, 
    0.00060132537723014729, 0.00059577436565743107, 0.00055668441941487826, 
    0.00049183547003540831, 0.00041042275984556008, 0.0003224364449568608, 
    0.0002380279611167144, 0.00016691804302496749, 0.00011788081935591214, 
    9.8344890259673061e-05, 0.00011413950139856556, 0.00016938505754850937, 
    0.00026650999915145889, 0.00040634196476457964, 0.00058823433976524836, 
    0.00081018849382474421, 0.0010689420810248637, 0.0013600363226780074, 
    0.0016778428788387109, 0.002015587941299427, 0.0023653898568309884, 
    0.0027183597055474734, 0.0030647866498790411, 0.0033944342643861939, 
    0.0036969503989820471, 0.0039623579687643783, 0.0041815943328421951, 
    0.0043470247034106384, 0.0044528951975895169, 0.0044956413692416588, 
    0.0044740473810683289, 0.0043892391163529321, 0.0042445316394771277, 
    0.0040451626702271148, 0.0037979646259447331, 0.0035110081458303742, 
    0.0031932396533204976, 0.0028541358375329543, 0.0025033749009736048, 
    0.0021505079559058604, 0.0018046565102491133, 0.0014742106386224718, 
    0.0011665600761747599, 0.00088787763458682886, 0.00064298413453127391, 
    0.00043530628016658058, 0.00026694177607008903, 0.00013880393474887984, 
    5.0821022323222881e-05, 2.1232703815485103e-06, -8.8022747423578533e-06, 
    1.59550871785445e-05, 7.3708159309547236e-05, 0.00016110255512539128, 
    0.00027399506521068795, 0.00040733280054069623, 0.0005550745346454873, 
    0.00071017099795806795, 0.00086465259003121848, 0.0010098334377969668, 
    0.0011366317033390063, 0.0012359970918404016, 0.0012994299076255936, 
    0.0013195230165584874, 0.001290490423381909, 0.001208635975097068, 
    0.0010727154074078905, 0.00088416512208036981, 0.00064717156634269755, 
    0.00036856534754754994, 5.7542124256790836e-05, -0.00027480866638174024, 
    -0.00061612380428693111, -0.00095350657113490458, -0.0012743153727362362, 
    -0.0015669311285508266, -0.0018214326722124756, -0.0020300993307340552, 
    -0.0021877264591353479, -0.0022917173209113452, -0.0023419710403532927, 
    -0.0023406003363943542, -0.0022915300628963769, -0.0022000303466208834, 
    -0.0020722345136905034, -0.0019146939078181166, -0.00173400182083233, 
    -0.0015364950765511531, -0.0013280336458549868, -0.0011138683424256983, 
    -0.00089856763821875873, -0.00068600737100196155, 
    -0.00047940155410274168, -0.00028138223490210319, 
    -9.4110634794387118e-05, 8.0580715322424833e-05, 0.0002410422468971006, 
    0.00038566696406915627, 0.00051277638639869022, 0.00062057366216311722, 
    0.00070716757385120036, 0.00077068740634231184, 0.00080946476656174266, 
    0.00082228180708410138, 0.00080861391595548465, 0.00076884640151294757, 
    0.00070441330821647847, 0.00061783457259823667, 0.00051263571281990586, 
    0.00039316569860162805, 0.00026432469015128174, 0.00013123541211011733, 
    -1.1192019507048304e-06, -0.00012826787427446369, 
    -0.00024660587019515985, -0.00035370605867159207, 
    -0.00044854523319354337, -0.0005316014790095133, -0.00060478383637040155, 
    -0.00067117617073842481, -0.00073461750892567072, 
    -0.00079916435891345733, -0.00086853408064993336, 
    -0.00094560066438972856, -0.0010320238692871578, -0.0011280610655934635, 
    -0.0012325600014326881, -0.0013431288976843451, -0.0014564279671433358, 
    -0.0015685433011101645, -0.0016753868762171943, -0.0017731019047295025, 
    -0.0018584041938972888, -0.0019288386585267626, -0.0019829052092512683, 
    -0.0020200369129007197, -0.0020404591940420139, -0.002044951346532483, 
    -0.0020345841266006734, -0.0020104695564377695, -0.0019735573300068985, 
    -0.001924534348266192, -0.0018638091102705103, -0.0017915859311257581, 
    -0.0017080181218958827, -0.0016133678877523739, -0.001508158044285667, 
    -0.0013932534806742423, -0.0012698453599819313, -0.0011393594787523754, 
    -0.0010032737555375456, -0.00086289519335884372, -0.00071912794028993366, 
    -0.00057228291431214793, -0.00042195072257589423, 
    -0.00026698426403759317, -0.00010559346835678698, 6.4444034291695929e-05, 
    0.00024544873993055064, 0.000439429697641974, 0.00064760434854087355, 
    0.00086993953937762082, 0.0011047430052843329, 0.001348392693716173, 
    0.0015952654098967639, 0.0018378758698576166, 0.0020672505581552018, 
    0.0022734987853576926, 0.0024464907273511194, 0.0025766060782863188, 
    0.0026554374717419837, 0.0026764144697044648, 0.0026353114003703931, 
    0.0025306263388341602, 0.0023638154528006117, 0.0021393592698459286, 
    0.0018646413061793052, 0.0015496178115212732, 0.0012062974483020223, 
    0.00084806694797796129, 0.00048892654260558653, 0.00014270991953538201, 
    -0.0001776287914606946, -0.00046062178435040443, -0.00069675433843796781, 
    -0.0008787871097142852, -0.0010019357065605495, -0.0010639406533336816, 
    -0.0010650236724729411, -0.0010077678524402073, -0.00089692945630309555, 
    -0.00073917923884220054, -0.00054280979381844522, 
    -0.00031737991977033217, -7.333249048323566e-05, 0.0001783966938469746, 
    0.00042675858602661174, 0.00066094339485504904, 0.00087069885671535864, 
    0.0010466509317232672, 0.0011806313615517405, 0.0012660315671070529, 
    0.0012981607982053549, 0.0012745778919715394, 0.0011953193785348467, 
    0.0010629786791306012, 0.00088258771389482043, 0.00066130068442382868, 
    0.00040788701305817954, 0.00013207738121360726, -0.00015616290461521011, 
    -0.00044733934796067052, -0.00073305969208298412, -0.0010065127842511607, 
    -0.0012627595242706599, -0.0014988436358154542, -0.0017137298937065244, 
    -0.0019081064632300363, -0.0020840775248248248, -0.0022447895154668867, 
    -0.0023940003217540178, -0.0025356253113046315, -0.0026733022591741611, 
    -0.0028099840251069141, -0.0029476045199515045, -0.003086844473412701, 
    -0.0032270204941171991, -0.0033661129045366176, -0.0035009311728570018, 
    -0.0036274150137092656, -0.003741039609678665, -0.0038372749060902097, 
    -0.0039120579531386288, -0.0039622027065608374, -0.0039856975132394777, 
    -0.0039818488373911561, -0.0039512456840391959, -0.0038955594200602759, 
    -0.003817222893580231, -0.0037190645855335858, -0.0036039744912020879, 
    -0.003474654660317481, -0.0033335187207862269, -0.0031827269510623073, 
    -0.0030243336717466303, -0.002860501261425381, -0.0026937203945211008, 
    -0.002526975577075991, -0.0023638147926665189, -0.0022083125322559473, 
    -0.0020649287678496, -0.0019382873163288246, -0.001832883381448542, 
    -0.0017527420006738185, -0.0017010351436556543, -0.0016796804806475491, 
    -0.0016889544002196082, -0.0017272086778389534, -0.001790718289460667, 
    -0.0018737315624150557, -0.00196874498074796, -0.0020669819828238668, 
    -0.002159052982792673, -0.0022357134488911099, -0.0022886434591190921, 
    -0.0023111408982063085, -0.0022986872395814005, -0.0022492951798647022, 
    -0.0021636292309955055, -0.0020449014698051835, -0.001898567952620586, 
    -0.0017318838479582338, -0.001553355237902124, -0.0013721217664415457, 
    -0.0011972983619104867, -0.0010373035256562163, -0.00089923999513615396, 
    -0.00078836744866996533, -0.00070771220455470194, 
    -0.00065786566858410365, -0.00063696282376661073, -0.0006408561501811199, 
    -0.00066347662666541279, -0.00069735171792846876, 
    -0.00073426950182550201, -0.00076603264611161998, -0.0007852220381936039, 
    -0.0007859174072359145, -0.00076424583956623976, -0.00071872813074985806, 
    -0.00065032548887054733, -0.00056218442454156171, 
    -0.00045912508400204616, -0.0003469126174651735, -0.00023144995682085548, 
    -0.00011801207980824082, -1.0638991824360667e-05, 8.8205494679937583e-05, 
    0.00017766310272925994, 0.00025822008151435183, 0.00033122332559254637, 
    0.00039829760640596411, 0.00046078358610426872, 0.00051932622605947417, 
    0.00057367045442998396, 0.00062269473538531799, 0.00066463485595574909, 
    0.00069745302493742106, 0.00071923637610192635, 0.00072855552564233064, 
    0.00072474535884395786, 0.00070806109344994815, 0.00067973791804771936, 
    0.00064194932973288092, 0.00059768678196652652, 0.00055056810721412124, 
    0.00050458864326849765, 0.00046384128689419676, 0.0004322411769592935, 
    0.00041328396751155185, 0.00040985779754199373, 0.00042413827396093701, 
    0.00045752633654248971, 0.00051060064624562022, 0.00058307839272206462, 
    0.00067375777717891571, 0.00078046931818310779, 0.00090005567604077791, 
    0.0010284074754579352, 0.0011605588887794664, 0.0012908593133359515, 
    0.0014132233306120379, 0.0015214408872868566, 0.0016095557698330568, 
    0.0016722701359393336, 0.0017053623326121689, 0.0017060431522780497, 
    0.0016732099611049059, 0.0016075405982316339, 0.0015114105393793824, 
    0.0013886164552740399, 0.0012439637018984687, 0.001082778719907058, 
    0.00091044774574438757, 0.00073202891449891823, 0.00055203421015054255, 
    0.00037435624136337547, 0.0002023530431585335, 3.9023012811250306e-05, 
    -0.00011277383997431619, -0.0002501361992704345, -0.00037002829442000785, 
    -0.0004693207171949464, -0.00054494838303683539, -0.00059417513529021746, 
    -0.00061493334476158974, -0.00060619045269021858, 
    -0.00056830257779754366, -0.00050330812347858787, 
    -0.00041507268968373308, -0.00030924590004381106, 
    -0.00019297562651590091, -7.4374897125525997e-05, 3.8195796544563181e-05, 
    0.00013695060584950728, 0.00021550101886892191, 0.00026955001147469464, 
    0.0002973677167406146, 0.00029997456224407736, 0.00028102073032781492, 
    0.00024637756880134889, 0.00020349723245896017, 0.000160609038643135, 
    0.00012585997088761816, 0.00010647522444671856, 0.0001080231622907388, 
    0.00013385867182900594, 0.00018479062340950517, 0.00025903333684914259, 
    0.00035241024260729417, 0.00045884798997964396, 0.00057105341573417362, 
    0.00068134539068457635, 0.00078247507324254477, 0.00086836639169399405, 
    0.00093466944659652317, 0.00097909332995875704, 0.001001519860731253, 
    0.0010039121815106579, 0.00099008079098795586, 0.00096532957865120715, 
    0.00093600437833279851, 0.00090894456743346834, 0.00089084840205940993, 
    0.00088756993553722565, 0.0009034172406366521, 0.00094052199101940038, 
    0.00099837978016956955, 0.0010736544185600719, 0.0011602817119909796, 
    0.0012498883435799054, 0.0013324857564839961, 0.001397364873956506, 
    0.0014340824487835584, 0.0014334231535917995, 0.0013882587192084305, 
    0.0012941953165919483, 0.0011499774305427429, 0.00095762327605497998, 
    0.00072227571569183618, 0.00045180434608559615, 0.0001562072939458599, 
    -0.00015311799216763156, -0.00046414290069914733, 
    -0.00076495594196381088, -0.0010444128339252945, -0.0012926650249389681, 
    -0.001501507041227331, -0.0016645905280014163, -0.0017774632686115496, 
    -0.0018374966350205083, -0.0018437192680710503, -0.0017966144863742835, 
    -0.0016979431984050811, -0.0015506102212604854, -0.0013586007193805709, 
    -0.0011269925881656543, -0.00086199192870246291, -0.00057094180789686686, 
    -0.00026224660490341061, 5.4838076854547444e-05, 0.00037055696901374063, 
    0.00067514124969010288, 0.00095938180562051521, 0.001215216832570875, 
    0.0014362677886337939, 0.0016182549684979927, 0.001759262947020995, 
    0.001859824304449945, 0.0019228154128515126, 0.0019532004198405855, 
    0.001957617840166721, 0.0019438734417347977, 0.0019203705848123199, 
    0.0018955118081386882, 0.0018771262528530582, 0.0018719832450994859, 
    0.0018854312211629247, 0.0019211711731527878, 0.0019811982593047664, 
    0.0020658728690693233, 0.0021740975534034297, 0.0023035362118557097, 
    0.0024508437564562482, 0.0026119039409136062, 0.0027820692246794468, 
    0.0029564026844329742, 0.0031299554951258412, 0.003298037778551107, 
    0.0034564872830778327, 0.0036018928823981591, 0.0037317568289309188, 
    0.003844561826527123, 0.003939769172463377, 0.0040177067675152226, 
    0.0040794147278192128, 0.0041264447102005719, 0.0041606512148468578, 
    0.0041840135394324756, 0.0041984664066456951, 0.0042057883901233254, 
    0.0042075027669075359, 0.0042047873687665292, 0.0041983784254160392, 
    0.004188452911316109, 0.0041745015832971568, 0.0041552371674525865, 
    0.0041285835059832526, 0.0040917866901009573, 0.0040416507202590988, 
    0.0039748642434782053, 0.003888383222017898, 0.0037797674658871985, 
    0.0036474370961401257, 0.0034908354184415543, 0.0033104568520959093, 
    0.0031077933462571724, 0.0028852289441613781, 0.0026459061626392371, 
    0.0023935859727807584, 0.002132495957115212, 0.0018671421691011008, 
    0.0016020810427044073, 0.0013416240598653662, 0.001089514681307833, 
    0.00084860685715180929, 0.00062061693517907995, 0.000405992292261085, 
    0.00020394950143826966, 1.2681684556326483e-05, -0.00017024525956028225, 
    -0.00034739745436226786, -0.00052092100874526486, 
    -0.00069201421725760418, -0.00086052117549622448, -0.0010247033284716415, 
    -0.0011812149580524168, -0.0013253000374211015, -0.0014511861671254866, 
    -0.0015526523056686426, -0.0016237142440972919, -0.0016593045077991214, 
    -0.0016558700963970011, -0.0016117737901192631, -0.00152747685107938, 
    -0.0014054324859172729, -0.0012497245222326222, -0.0010655494064934511, 
    -0.00085857998072553165, -0.00063437536539122635, 
    -0.00039794241250835851, -0.00015349476571819957, 9.5536831576416737e-05, 
    0.00034630661542587216, 0.00059622514424455427, 0.00084263771695561383, 
    0.0010825681205886492, 0.0013126107983969999, 0.0015290010000147385, 
    0.0017278406408332168, 0.0019054923068456044, 0.0020590373535281422, 
    0.0021867637599134299, 0.0022885709695293988, 0.0023662202870309425, 
    0.0024233981488499083, 0.0024655783946179836, 0.0024997384956268734, 
    0.0025339887664640195, 0.0025771527557950538, 0.0026383200083734217, 
    0.0027264038449672334, 0.002849654867345802, 0.0030151520339578718, 
    0.0032282613820769591, 0.0034920900234533103, 0.0038069849262280537, 
    0.0041701724694591016, 0.0045755603985300798, 0.0050137791445107613, 
    0.0054724486286054494, 0.0059366638276440011, 0.0063896428121623513, 
    0.0068134728374393671, 0.0071899263939309123, 0.0075012676374497768, 
    0.0077310496176203882, 0.0078648584281876266, 0.0078909930875806535, 
    0.007801062276264612, 0.0075904761206679839, 0.0072587961251441759, 
    0.0068099357001899152, 0.0062521655343646242, 0.0055978957705276992, 
    0.0048632471652344383, 0.004067369185965241, 0.0032315298550529203, 
    0.002378013583980057, 0.0015289265702394207, 0.00070505667694170085, 
    -7.5127443402548267e-05, -0.00079621158202624427, -0.001446316825908294, 
    -0.0020172945141952482, -0.0025046658123839259, -0.0029073476614030458, 
    -0.0032271613354438785, -0.0034682632730739993, -0.0036364974794751309, 
    -0.0037388011844608389, -0.0037827100952159878, -0.0037759702759847828, 
    -0.0037262369580391441, -0.0036408447274721002, -0.0035266329398665852, 
    -0.0033898066450291212, -0.0032358419984397676, -0.0030694167938872126, 
    -0.0028943660410539833, -0.0027136632026325633, -0.0025294159187805644, 
    -0.0023428446381255959, -0.0021542763418344827, -0.0019631095218125161, 
    -0.0017678375337338813, -0.0015661064201818108, -0.0013549144457886213, 
    -0.0011308901278258207, -0.00089068300332504702, -0.00063144100435027258, 
    -0.00035130582324548307, -4.9854273883803658e-05, 0.00027156076932565809, 
    0.00060964835460081287, 0.00095923291524232775, 0.0013135073793903683, 
    0.0016644718455762512, 0.0020034953852584819, 0.0023219741582085327, 
    0.0026119817001294967, 0.002866869703456934, 0.003081762437619436, 
    0.0032538842869816197, 0.0033826519835505019, 0.0034695612845383654, 
    0.003517801981819738, 0.003531680339516105, 0.0035159003576033482, 
    0.0034747876292141522, 0.0034116275038538198, 0.003328200458320859, 
    0.0032246833673465649, 0.003099920366564641, 0.0029520028770140491, 
    0.0027790231171001488, 0.0025798505146922396, 0.0023547230910150839, 
    0.0021055817056864399, 0.0018360792147382003, 0.0015512603924284533, 
    0.0012569676373340893, 0.00095906391036979714, 0.00066262395605114763, 
    0.00037119328838035434, 8.6366088161619084e-05, -0.00019224358274467503, 
    -0.0004665849253649119, -0.00073932898578435587, -0.0010128090980481058, 
    -0.001287936183812087, -0.001563303913947879, -0.0018346405839530346, 
    -0.0020946655242244433, -0.0023333491966842507, -0.0025385850982871223, 
    -0.0026972087689814397, -0.002796270068273161, -0.0028244223120282223, 
    -0.0027732262173234988, -0.0026381736055837088, -0.0024192811905727075, 
    -0.0021211381389103535, -0.0017524589197057006, -0.0013252123569554182, 
    -0.00085352995819581393, -0.00035255948463495045, 0.00016254954829899324, 
    0.00067744841300619802, 0.0011791172107199896, 0.0016561775915508556, 
    0.0020990517717883552, 0.0025000695198373127, 0.0028535796786839313, 
    0.0031560556989439449, 0.0034062248779574483, 0.0036051010378349542, 
    0.0037559047116104303, 0.0038637896090137486, 0.0039353805802442455, 
    0.0039781497385724916, 0.0039996888654988422, 0.0040069747579094157, 
    0.0040057044193140736, 0.0039997727831744111, 0.0039909479714513264, 
    0.0039787604186486761, 0.003960608193663135, 0.0039320279937718359, 
    0.0038871184835624364, 0.0038190126312833373, 0.003720409896644794, 
    0.0035840934009974072, 0.0034034620185113646, 0.003173063605179713, 
    0.0028890721643698271, 0.0025497177755324555, 0.0021555615567260748, 
    0.0017096020401331622, 0.0012172153711772949, 0.00068594179015838363, 
    0.00012516881117549452, -0.00045423726381004366, -0.0010403167808188619, 
    -0.0016203833305330755, -0.0021813957662950309, -0.0027103217529066284, 
    -0.003194521418286596, -0.0036221882242098045, -0.0039828136841685733, 
    -0.0042676755842361103, -0.0044702975956422558, -0.0045868613087806046, 
    -0.0046164985778243597, -0.0045614100815873004, -0.0044268009720519978, 
    -0.0042205723966709848, -0.0039527909720272689, -0.003634979233126087, 
    -0.0032793130790565415, -0.0028978524765787819, -0.0025019332310491759, 
    -0.0021017722503747175, -0.001706332041298579, -0.0013233686242386299, 
    -0.00095958442833955944, -0.00062075306870736395, 
    -0.00031178061971758985, -3.6683523973302383e-05, 0.00020147826812898218, 
    0.00040063800612849608, 0.00055971506564739802, 0.00067857058191676388, 
    0.00075798442836032829, 0.00079970882288741608, 0.00080655239440955654, 
    0.0007825099884149892, 0.00073279760858941442, 0.00066375218356980832, 
    0.00058255163367667499, 0.00049676531237255375, 0.00041380516330352017, 
    0.00034040834558068408, 0.00028219248473868171, 0.00024336545339120164, 
    0.00022657859750490077, 0.00023292346370132815, 0.00026209311344679441, 
    0.00031264782560676318, 0.00038237787844064091, 0.0004686357126315818, 
    0.00056864733182180596, 0.00067970518356646288, 0.0007992775912970656, 
    0.00092504296819809358, 0.0010548880673459742, 0.001186900346943531, 
    0.0013193708778449001, 0.0014508160027107216, 0.0015800083965847272, 
    0.0017060113490689377, 0.0018281877991571346, 0.0019462223364337338, 
    0.0020601220744315765, 0.0021701598221378149, 0.0022767747269554785, 
    0.0023803622720353873, 0.0024810510273055018, 0.0025784346837311738, 
    0.0026714081307455183, 0.0027581362873766056, 0.0028361906634061132, 
    0.0029027757369236729, 0.0029550147211862198, 0.0029902504124988353, 
    0.0030062997903873307, 0.0030016352377312421, 0.0029755059239999792, 
    0.0029279555172621778, 0.0028597758415990133, 0.0027723454587417567, 
    0.0026674319764569167, 0.0025469593249911773, 0.0024128052873312596, 
    0.0022666689809176452, 0.002110018467015046, 0.0019441334968944486, 
    0.0017702001920688654, 0.0015894424028044701, 0.0014032449428909685, 
    0.0012132902671621077, 0.0010216634598420892, 0.0008309476452391456, 
    0.00064430331129958706, 0.00046548063222961024, 0.00029879716948757649, 
    0.00014899840216924209, 2.1025567935707912e-05, -8.0306680266715625e-05, 
    -0.00015067187970038028, -0.00018665158665053812, 
    -0.00018610937207218101, -0.0001485461255424571, -7.5393690632570164e-05, 
    2.9763882623919379e-05, 0.00016107180002784591, 0.0003103657509704867, 
    0.00046731069977962826, 0.00061973904013782959, 0.00075425354790308811, 
    0.00085708811624027586, 0.00091521972326746674, 0.00091760838795261425, 
    0.00085648847769236513, 0.0007285231516653319, 0.00053565325044670664, 
    0.00028549823550417798, -8.8328623834206012e-06, -0.00032958019817393516, 
    -0.0006557424502808886, -0.00096487647791475815, -0.0012350135074574243, 
    -0.0014464254096413251, -0.0015831272864543985, -0.0016340111375346715, 
    -0.0015935927544658279, -0.0014623830864775357, -0.0012469010760780097, 
    -0.00095931548481427876, -0.00061674415645370114, 
    -0.00024018469265022391, 0.00014693941654910251, 0.00052052026562571913, 
    0.000857716911806912, 0.0011388555775220172, 0.0013491248152339127, 
    0.0014798195230645236, 0.0015289615465172023, 0.0015013066374782568, 
    0.0014076721986203645, 0.0012637230386786835, 0.001088330008562051, 
    0.00090164115456095118, 0.00072313886149521448, 0.00056985073349122425, 
    0.00045495061974391355, 0.00038683832009844365, 0.00036884163560991503, 
    0.00039940087058283993, 0.00047274545988267095, 0.0005798869594475796, 
    0.0007097528294399048, 0.00085038568774050056, 0.0009900187369551363, 
    0.001118037451188038, 0.0012257228115180791, 0.0013068430777055779, 
    0.0013580359952310721, 0.0013789887104086547, 0.0013723583343288662, 
    0.0013434039283338911, 0.0012994249255647071, 0.001249058383438334, 
    0.0012015623084198363, 0.0011661371231741309, 0.0011513432631680425, 
    0.0011645729375475851, 0.001211636674462049, 0.0012964088936906581, 
    0.0014205588419341517, 0.0015833711418530502, 0.0017816763458080125, 
    0.0020099307819173773, 0.0022604309793076548, 0.0025237471049678159, 
    0.0027893172308288941, 0.0030462086826471076, 0.0032839675028345215, 
    0.0034934301172449174, 0.0036674305554347973, 0.003801296148566979, 
    0.0038930594842376091, 0.0039433903828383398, 0.0039552308812932689, 
    0.0039332261945337395, 0.0038830978598150476, 0.003811008674736379, 
    0.0037230365654210085, 0.0036247649070437421, 0.0035209739891307514, 
    0.0034155363260291254, 0.0033114616222474627, 0.003211153385153852, 
    0.0031167495292153688, 0.0030304550108943345, 0.0029547152765925437, 
    0.002892141807740813, 0.0028451914377956729, 0.0028156273855381472, 
    0.002803953662616532, 0.0028089136784536679, 0.0028272970546227437, 
    0.0028540827791097133, 0.0028828982002621724, 0.0029067345914217161, 
    0.0029187053371301352, 0.0029127023651174099, 0.0028839131461732169, 
    0.0028291145448587863, 0.0027467862400009984, 0.0026370933136519899, 
    0.0025017905172601287, 0.0023440745560279735, 0.002168350741307847, 
    0.0019800005702559544, 0.0017850167612385507, 0.0015896131682317117, 
    0.0013998194278082524, 0.0012211414073012906, 0.0010583574049441409, 
    0.00091552865093348439, 0.00079618468747650012, 0.00070363901554806776, 
    0.00064135024900552372, 0.00061315349506880796, 0.00062333865884708526, 
    0.00067646484268943808, 0.00077695731891853611, 0.00092856157402030845, 
    0.0011336484179758841, 0.0013925603132464192, 0.001703038257342781, 
    0.0020598898755395927, 0.0024549207704757446, 0.0028771798786319646, 
    0.0033134790751810704, 0.0037490687978125178, 0.0041684865589574887, 
    0.0045564339114854526, 0.0048986214741126802, 0.0051826016817411152, 
    0.0053984532802900395, 0.0055393702518760548, 0.0056021093386358226, 
    0.00558726864264124, 0.0054994072305360603, 0.0053469085856776505, 
    0.0051416171689922484, 0.0048981568677242378, 0.0046330506082479473, 
    0.0043636779614393975, 0.0041071884787800264, 0.0038794814168921403, 
    0.0036943767480550793, 0.0035629947034252155, 0.0034933423724739345, 
    0.0034900846909680771, 0.0035544884401713149, 0.0036844494827488069, 
    0.0038746781539058047, 0.004116981494772908, 0.0044006618966161738, 
    0.004713038722948956, 0.0050400640132682948, 0.0053670103085676499, 
    0.0056792428924785834, 0.0059630162238703197, 0.0062062499478131531, 
    0.0063991669354334021, 0.0065348070072560067, 0.0066092644740609018, 
    0.0066217376602185178, 0.0065743234440113311, 0.0064716179978871876, 
    0.0063201578437553632, 0.0061277496902154126, 0.0059027669371540291, 
    0.0056535230835232826, 0.0053877318227827991, 0.0051121294672063092, 
    0.0048323217067666535, 0.0045528076141333673, 0.0042771696765707672, 
    0.0040084081731854926, 0.0037493350069976953, 0.0035029445437770399, 
    0.0032727162480629237, 0.0030627688542560431, 0.0028778262393752596, 
    0.0027229800527706432, 0.0026032244495367961, 0.0025228325874598018, 
    0.0024845817439097116, 0.0024890707636890611, 0.0025341684702427356, 
    0.0026147245049565537, 0.0027227306775354115, 0.0028477722752541122, 
    0.0029778657482289637, 0.0031004180766685888, 0.003203306567602344, 
    0.0032757442101248816, 0.00330893351694819, 0.0032963335263407386, 
    0.0032335895416241867, 0.0031181036065146593, 0.0029484492129255523, 
    0.0027237931472239314, 0.0024434722342816999, 0.0021069158666885191, 
    0.0017139499607872115, 0.0012653999621265485, 0.00076387746361402048, 
    0.00021447234309433197, -0.00037472882395543714, -0.0009926142422010053, 
    -0.0016253888460555218, -0.002257456762126667, -0.0028725779565569958, 
    -0.0034553217268043445, -0.0039924670578877636, -0.0044742070141667069, 
    -0.0048948484239446834, -0.0052529478684003048, -0.0055507956899823498, 
    -0.0057934448348346008, -0.005987420353973095, -0.0061393752322792487, 
    -0.0062549543900281817, -0.0063379689196838875, -0.0063899686541015058, 
    -0.0064102956391425764, -0.0063964769224341151, -0.0063450026468336957, 
    -0.0062522898844090688, -0.0061156841646895508, -0.0059343738368241488, 
    -0.0057099039479175922, -0.0054463231248595839, -0.0051498381701213531, 
    -0.004828097679788073, -0.0044892806155430905, -0.004141138219904728, 
    -0.0037902154220768197, -0.0034412533074493577, -0.0030969681277430807, 
    -0.0027580866999999641, -0.0024236576876460244, -0.0020916212428145186, 
    -0.0017594364609349608, -0.0014248490751029659, -0.0010864707479622457, 
    -0.00074434654632872033, -0.00040020780951242885, 
    -5.7524019112929135e-05, 0.00027869129924521104, 0.00060227201857195013, 
    0.00090648905199180627, 0.0011847374003525978, 0.0014311969188708249, 
    0.0016414355986013509, 0.0018128527706404373, 0.0019449910974896169, 
    0.0020395966038624495, 0.0021005324961589121, 0.0021336070292022713, 
    0.0021462095703802262, 0.0021469179507953148, 0.0021450202920171167, 
    0.0021498679722827731, 0.0021701619604330888, 0.0022131427312844527, 
    0.0022838415549191887, 0.0023842656029713894, 0.0025129050689560724, 
    0.0026644174593521723, 0.0028297448898324555, 0.0029965615427949709, 
    0.0031501185667373159, 0.0032744582799631937, 0.0033537609892358776, 
    0.0033738519319039682, 0.0033236604617765276, 0.003196587575565618, 
    0.0029915272983079642, 0.0027134481806129524, 0.0023733565677268786, 
    0.0019875389436306581, 0.0015761426664195298, 0.0011612047565981317, 
    0.00076446033235804149, 0.00040507392474477787, 9.7726445059284801e-05, 
    -0.00014872201269709511, -0.00033184729145124261, 
    -0.00045548088835270983, -0.00052880734890649794, 
    -0.00056475815843129136, -0.0005780125702076087, -0.00058277102767068318, 
    -0.00059048944056002903, -0.0006080647980147365, -0.00063670904783206693, 
    -0.00067184346651225752, -0.0007039480414029783, -0.0007199992079063109, 
    -0.00070508224748538949, -0.0006439500956656706, -0.00052243523648463626, 
    -0.00032877936906114662, -5.4701096196397517e-05, 0.00030376006065169236, 
    0.00074585307356226087, 0.0012660582282107606, 0.0018544087885356683, 
    0.0024971498047561286, 0.0031776036993109301, 0.0038771539464259016, 
    0.0045762106936219097, 0.005254995932461399, 0.0058941990521416609, 
    0.0064754896879792223, 0.0069821579133742149, 0.0073997635054583828, 
    0.00771691632329674, 0.0079259344742972082, 0.0080232956655683519, 
    0.0080096465875196289, 0.00788938326689273, 0.0076698847917891898, 
    0.0073606221587497727, 0.006972090254262096, 0.0065149694344688591, 
    0.0059994423056112366, 0.0054348408899759096, 0.0048294643636971344, 
    0.0041907198191206531, 0.0035252846557403614, 0.0028393292459745539, 
    0.0021386638152999077, 0.0014289143681114446, 0.00071575501383491042, 
    5.2567994788513175e-06, -0.00069573940189455183, -0.0013794141032408664, 
    -0.0020370185246160123, -0.0026592018690101346, -0.0032365209049454767, 
    -0.0037599266214866744, -0.0042211226666063655, -0.0046126954174351559, 
    -0.0049279136962521036, -0.005160353949532669, -0.0053033409341923573, 
    -0.0053494051990022121, -0.0052901272657019209, -0.0051165070991559345, 
    -0.0048198374234388781, -0.0043930644749754048, -0.0038323302154411707, 
    -0.0031384026423036029, -0.0023177996384909538, -0.0013832861602674112, 
    -0.00035376099385831731, 0.00074643367942051281, 0.0018889004224897966, 
    0.0030430066094034964, 0.0041779456463509612, 0.005264858442005603, 
    0.0062788068797946387, 0.0072003358865214053, 0.0080163516925541699, 
    0.0087202708444738177, 0.0093112588398592093, 0.0097928936060855381, 
    0.010171300429915913, 0.01045335359837327, 0.010645208886923786, 
    0.01075135845765568, 0.010774354463594208, 0.010714788420493152, 
    0.01057137749373524, 0.010340844162040719, 0.010017552692987861, 
    0.0095933228866316167, 0.009057606061701402, 0.0083984192301509771, 
    0.007603729650498884, 0.0066635521684207969, 0.0055720213255976625, 
    0.0043296543678288321, 0.0029452365009934004, 0.0014371032316822761, 
    -0.00016644496904930398, -0.0018279998989277613, -0.0035032436878654431, 
    -0.0051442295542587996, -0.0067034799588610184, -0.0081379618013445558, 
    -0.0094123974697689732, -0.010501006823960941, -0.011387565564652216, 
    -0.012063968942186721, -0.01252808839513086, -0.012782100933891535, 
    -0.012831825566629564, -0.012687194159092606, -0.012362985631728163, 
    -0.011879332973461623, -0.011261474281429979, -0.010538735346644125, 
    -0.0097430231410246971, -0.0089073012024570922, -0.0080637882868102324, 
    -0.0072425034390615995, -0.0064698560195123721, -0.0057677111388747156, 
    -0.0051525670626363347, -0.004635036352368129, -0.004219622141978777, 
    -0.0039047048736142271, -0.0036828011196423441, -0.003541004728926829, 
    -0.0034616785835500036, -0.0034235796905820537, -0.0034032137040769456, 
    -0.0033765359893487964, -0.0033208909310479579, -0.0032170129364305234, 
    -0.0030511736975671342, -0.0028175298365939452, -0.0025199369653558764, 
    -0.002173094511958764, -0.0018021020159714196, -0.0014401766980463059, 
    -0.0011242524670064032, -0.00088905808978875919, -0.00076083266486316943, 
    -0.00075186004800772846, -0.00085778285809022449, -0.0010585100392369181, 
    -0.0013224111291887835, -0.0016129806182446796, -0.0018963896786758922, 
    -0.0021489225357505812, -0.0023624657081512727, -0.0025483555970082158, 
    -0.0027382152981976797, -0.0029827793946227239, -0.0033466913928722405, 
    -0.0039006918456644538, -0.0047102940645081942, -0.0058233455745795261, 
    -0.0072586840884125581, -0.0089984838456853358, -0.010987438655257349, 
    -0.013138771567120792, -0.015345134700747651, -0.017494080324160163, 
    -0.019484279198014598, -0.021237547747770782, -0.022707163205792493, 
    -0.023879069586414725, -0.024768902844104646, -0.02541705253004798, 
    -0.025882207696477463, -0.026236589809176387, -0.026560206619105027, 
    -0.026934367607977034, -0.027433962785997187,
  // Fqt-Na(9, 0-1999)
    0.99999999999999989, 0.99040742321880726, 0.96223180144907561, 
    0.91720972088628461, 0.85801877204030685, 0.78799231111268753, 
    0.71078729265802876, 0.6300538591733692, 0.54914906984793166, 
    0.47092419712103012, 0.39759899872660953, 0.3307210667882633, 
    0.27119672156409352, 0.21937315434044966, 0.17514962241399143, 
    0.13809776396506379, 0.10757558854115666, 0.082825325976946806, 
    0.06305047002815703, 0.047471593724292729, 0.035363052816771878, 
    0.026074170353497204, 0.019038725957462678, 0.013776229769951319, 
    0.0098878628164419946, 0.0070492257613861018, 0.0050014469889423929, 
    0.0035417195039913782, 0.0025139450689155417, 0.0017999506793509343, 
    0.0013115084058623148, 0.00098334157128917958, 0.00076720702453887614, 
    0.00062709227077973489, 0.00053554977710167269, 0.0004711162135883994, 
    0.00041672486634551333, 0.00035891657759653346, 0.00028762357894275553, 
    0.0001962423507172769, 8.1755361512740729e-05, -5.5300741578293662e-05, 
    -0.00021111812044213261, -0.00037918670862289316, 
    -0.00055111417740651906, -0.00071763949330425568, 
    -0.00086972235758753713, -0.00099962363083933329, -0.0011018259365436042, 
    -0.0011736922072224693, -0.0012157411396203285, -0.0012314778187808113, 
    -0.0012268054744970771, -0.0012090798733692346, -0.001185957203813729, 
    -0.0011642047756923229, -0.0011486577108718958, -0.0011414855172472104, 
    -0.0011418632490059694, -0.0011460966579247122, -0.0011481778053986367, 
    -0.0011407003995837473, -0.0011160128624130039, -0.0010674660331305595, 
    -0.00099060663216601463, -0.00088413592990274799, 
    -0.00075050707602060689, -0.00059601495142127116, 
    -0.00043031663667946114, -0.00026538705372258152, 
    -0.00011406169879556188, 1.1612481811191675e-05, 0.0001019123594836739, 
    0.00015061828010554188, 0.00015563904929433462, 0.00011906168146275423, 
    4.6650774226263486e-05, -5.3071740085648046e-05, -0.00016998301499564884, 
    -0.00029357625717496279, -0.00041406399019130319, 
    -0.00052324340181387715, -0.00061503891450327285, 
    -0.00068570322665170832, -0.00073368854742186221, 
    -0.00075928100546924506, -0.00076405410064574056, 
    -0.00075029249837445721, -0.00072047409614837954, 
    -0.00067690216124406352, -0.00062157787773448124, 
    -0.00055627748913380549, -0.00048280464857771024, 
    -0.00040331453150861717, -0.00032058891351199989, 
    -0.00023817540213321451, -0.00016033446951448934, 
    -9.1789486751409468e-05, -3.7314815599061313e-05, 
    -1.2314979942972502e-06, 1.3113998390595167e-05, 3.7968429811255258e-06, 
    -2.936406606124267e-05, -8.466414921970395e-05, -0.00015855318211787815, 
    -0.00024585488676858618, -0.00034012694177573959, -0.0004341187380306463, 
    -0.00052027053828733385, -0.00059119863790305701, 
    -0.00064011524908947725, -0.00066116498954178966, 
    -0.00064966251928479351, -0.00060225227543633277, 
    -0.00051702210401663527, -0.00039356947611715636, 
    -0.00023304902370823691, -3.8170866038999272e-05, 0.00018686171811771251, 
    0.00043648346165263706, 0.00070397779610391689, 0.00098174967476260958, 
    0.0012616461134868668, 0.0015353141529332766, 0.0017945668572184161, 
    0.002031760105756582, 0.0022401807892391142, 0.0024144147745701738, 
    0.0025507038560490334, 0.0026472694026658207, 0.0027045507163481254, 
    0.0027253056337609993, 0.002714501277200348, 0.0026789587229827795, 
    0.0026267412677836474, 0.0025663593114281891, 0.0025059008844195894, 
    0.002452215610814908, 0.0024102675937565134, 0.0023827753925707205, 
    0.00237015600109206, 0.0023707829210529137, 0.0023814825833364459, 
    0.0023981658025701001, 0.002416500035983231, 0.002432472992473499, 
    0.002442817061596356, 0.0024452113482699659, 0.0024382885669129331, 
    0.0024214829136794706, 0.0023947644703450825, 0.0023583635382728669, 
    0.002312495437394136, 0.002257162106485416, 0.0021920085233094835, 
    0.0021162492251574237, 0.0020286667030859377, 0.0019276987086304877, 
    0.0018116306328423756, 0.001678872645957497, 0.0015282827065725064, 
    0.0013594494604670074, 0.0011728476422009412, 0.0009698335404537368, 
    0.00075249852480815732, 0.00052347480099817318, 0.00028579090149019457, 
    4.2856390800621869e-05, -0.00020143144895917199, -0.00044252721503730162, 
    -0.00067510326946546224, -0.0008930218803319906, -0.0010894429976975753, 
    -0.0012570778077444235, -0.0013885823052040963, -0.0014770390490793893, 
    -0.0015164903643428891, -0.0015024782670711736, -0.001432517114876576, 
    -0.0013064646385635332, -0.0011267597074293661, -0.0008984654715999971, 
    -0.00062913432221061805, -0.00032846251682507868, 
    -7.7418645478537912e-06, 0.00032084449676870991, 0.00064505613811060777, 
    0.00095347223248824873, 0.0012363441140523894, 0.0014863099381625072, 
    0.0016988740115021724, 0.001872563328473626, 0.0020087221085189431, 
    0.0021109606937526697, 0.0021843538423180148, 0.0022345000773363872, 
    0.0022666152459832286, 0.0022847785970556232, 0.002291460957548945, 
    0.0022873750708088791, 0.0022716832139803014, 0.002242505548043503, 
    0.0021976450204701341, 0.0021354002460520025, 0.0020553228006014567, 
    0.0019587855061794913, 0.0018492788692296195, 0.001732372559391861, 
    0.001615362228845866, 0.0015066609153445056, 0.0014149972240747443, 
    0.0013485625806382694, 0.0013141877513528214, 0.0013166491021724118, 
    0.0013581900006584908, 0.0014382896558264374, 0.001553700160125488, 
    0.0016987182494313641, 0.0018656497016995947, 0.0020453910672778878, 
    0.0022280562990724187, 0.0024035738126697709, 0.0025622118783036009, 
    0.0026950112109656752, 0.0027941424161388069, 0.0028532132458725483, 
    0.0028675758286737579, 0.0028346537079701941, 0.0027542764236332014, 
    0.0026290031867205409, 0.0024643407676407277, 0.0022687825645747433, 
    0.002053586352793874, 0.0018322562337981642, 0.0016197031955634427, 
    0.001431173213563044, 0.0012810323401775299, 0.0011815432335377397, 
    0.0011417964150265492, 0.0011669037506783914, 0.0012575624372929786, 
    0.0014100066538467052, 0.0016163290938159972, 0.0018651061242761688, 
    0.0021422349339349214, 0.0024318646803468198, 0.0027173486408606376, 
    0.0029821300185672523, 0.003210525892718496, 0.0033884036890693154, 
    0.0035037526391564263, 0.0035471901198353109, 0.0035123998422339352, 
    0.0033965212149007101, 0.0032004305474023298, 0.0029288597024192103, 
    0.0025902590377301859, 0.0021963436468002335, 0.0017613255781308967, 
    0.0013008667257102791, 0.00083087974127620608, 0.00036630317660026214, 
    -7.9987241847648467e-05, -0.00049801731274714774, 
    -0.00088119881113351141, -0.0012263880078559122, -0.0015335267634421124, 
    -0.0018049110684182816, -0.0020442337571356401, -0.0022555473336465519, 
    -0.002442340877070744, -0.0026068770746020867, -0.0027498640432860708, 
    -0.0028704835795810061, -0.0029667194710129839, -0.0030359100296668134, 
    -0.0030753981667845996, -0.0030831724465326684, -0.0030583879229392668, 
    -0.0030017095882396193, -0.0029154267703222127, -0.0028033403276326984, 
    -0.0026704641522392646, -0.0025225883821371935, -0.0023657786329413211, 
    -0.0022058977539911643, -0.0020482057785603117, -0.0018970920598743554, 
    -0.0017559364110368624, -0.0016271129184022132, -0.0015120762209504548, 
    -0.0014114893188963927, -0.0013253770453113556, -0.0012532559413994048, 
    -0.0011942683015720833, -0.0011473219700908401, -0.0011112457575045214, 
    -0.0010849680934718743, -0.0010676887163400543, -0.0010590400587630249, 
    -0.0010591946549287439, -0.0010689093890759536, -0.0010894944236266037, 
    -0.0011226984690431475, -0.00117053483155148, -0.0012350335451959832, 
    -0.0013179370774177414, -0.0014203652420074426, -0.0015424719806729238, 
    -0.001683122585861068, -0.0018396534711708386, -0.0020077481331281532, 
    -0.0021814565543151034, -0.0023533874783045962, -0.0025150627843438327, 
    -0.0026574369258191141, -0.0027715179378463291, -0.0028490463348409501, 
    -0.0028831018161556612, -0.0028685534868591045, -0.002802276116628314, 
    -0.0026831296606749863, -0.002511754721903031, -0.0022902994938058126, 
    -0.0020221799465665819, -0.0017119341579158386, -0.0013651513165209503, 
    -0.00098843739930894918, -0.00058933967440236721, 
    -0.00017619239358397421, 0.0002421270023141045, 0.00065648093009356269, 
    0.0010577994227296136, 0.0014374048565009398, 0.0017873456020112461, 
    0.0021007368483876858, 0.0023720952609866037, 0.0025976205998869415, 
    0.0027753897553301574, 0.0029054068027596805, 0.0029894982129767145, 
    0.0030310489161571169, 0.0030346164073652756, 0.0030054662579585608, 
    0.0029490974389496786, 0.0028708271119859304, 0.0027754838462646166, 
    0.0026672617729167044, 0.002549731580226795, 0.0024260175150979868, 
    0.0022990674665787207, 0.0021719484950565044, 0.0020480730764042407, 
    0.0019313032907080844, 0.0018258888184999979, 0.0017362452794743328, 
    0.0016665703172450278, 0.0016203395517782372, 0.0015997459237999108, 
    0.0016051705724078216, 0.0016347692562413809, 0.0016842553798766878, 
    0.001746954968701108, 0.0018141288466074061, 0.001875585058758052, 
    0.0019204982394606101, 0.0019383459194396921, 0.0019198330163156083, 
    0.0018576752897511476, 0.0017471301060211482, 0.0015862380970651934, 
    0.001375749003884162, 0.0011188219342276244, 0.0008205478440176891, 
    0.00048739571518564026, 0.00012666123784858357, -0.00025403928596615658, 
    -0.00064717634631951014, -0.0010455800401398731, -0.001442559455973343, 
    -0.0018318637080668898, -0.0022075130446492946, -0.0025635390074643374, 
    -0.0028937213780291277, -0.0031913823035107656, -0.003449312766004417, 
    -0.0036598838155425016, -0.0038153831612884785, -0.0039085581624455808, 
    -0.0039333487404265679, -0.003885718442718648, -0.0037644822395103, 
    -0.003571956034970862, -0.0033142738659135487, -0.0030012662519097108, 
    -0.0026458802202181503, -0.0022632250784941146, -0.0018693849814302682, 
    -0.0014801746028269161, -0.0011100010229120778, -0.00077097237872230794, 
    -0.00047235412208418431, -0.00022039632181743098, 
    -1.8499453657457873e-05, 0.00013238862866956944, 0.00023328465734851335, 
    0.00028672442645453881, 0.0002964736270735495, 0.00026741102768063361, 
    0.00020557453486283993, 0.00011824570844357833, 1.3970324522681165e-05, 
    -9.7596246933185846e-05, -0.00020608213030259598, -0.0003010164773245889, 
    -0.00037262004967697233, -0.00041267666965445684, 
    -0.00041536004017486878, -0.00037788216101806635, 
    -0.00030084201596909281, -0.00018821404588045912, 
    -4.6936381412859222e-05, 0.00011380497231057993, 0.00028351848196604646, 
    0.00045139444274608993, 0.00060724545693324609, 0.00074224698631240849, 
    0.00084945337456866494, 0.00092404569948842928, 0.00096330846510712107, 
    0.00096641779296715072, 0.00093407664559656324, 0.0008681070593679497, 
    0.00077108596409237768, 0.00064610772647379013, 0.00049672206739522265, 
    0.0003270543864981324, 0.00014205293146883521, -5.2246650533370866e-05, 
    -0.00024857216565623235, -0.00043848050098054415, 
    -0.00061269924500965218, -0.00076172933023773977, -0.000876630922106754, 
    -0.00094988430296296907, -0.00097619329716576257, 
    -0.00095310749750657231, -0.00088137001968519599, 
    -0.00076490834176760295, -0.00061044603014222992, 
    -0.00042675272166877815, -0.00022363938528444818, -1.086729499527955e-05, 
    0.00020283271456440346, 0.00041045992623600067, 0.00060710872515896074, 
    0.00079003593845809153, 0.0009584607653470125, 0.0011131552988001734, 
    0.0012558637282364708, 0.0013886284469577543, 0.0015131335701517163, 
    0.0016301802965768479, 0.0017393912650814755, 0.0018391850251747298, 
    0.0019269986249217874, 0.001999706234391233, 0.0020541495022524895, 
    0.0020876885525583011, 0.0020987005504420442, 0.0020869752701824546, 
    0.0020539441180771369, 0.0020027277482168706, 0.0019379715501511244, 
    0.0018654835377725758, 0.0017917207243307177, 0.0017231651178710409, 
    0.0016656982687812052, 0.0016240343755009163, 0.0016013254275731316, 
    0.0015989662972964635, 0.0016166557735761713, 0.0016526686802832316, 
    0.0017042859951885176, 0.0017683104814106537, 0.0018415285963315042, 
    0.0019210648581214184, 0.0020045460699526741, 0.0020900446406307213, 
    0.0021758507017237728, 0.0022601130844065479, 0.0023404791736601127, 
    0.0024138344219704106, 0.0024762351477221394, 0.0025230510470821087, 
    0.0025492976846015983, 0.0025500498933329376, 0.0025208526796533428, 
    0.0024580405229012491, 0.0023589226440251863, 0.0022218438663152555, 
    0.0020461587704287366, 0.001832159458812078, 0.0015810147976883118, 
    0.0012947507611311309, 0.00097630197866031897, 0.00062960417826712868, 
    0.00025967675320601115, -0.00012735098258609287, -0.00052430302197524503, 
    -0.00092314698269467402, -0.0013153071655969423, -0.0016920466484617366, 
    -0.0020449001949995951, -0.0023660770440697169, -0.0026488132057553501, 
    -0.0028876535416846004, -0.0030786647244271759, -0.0032196000239074138, 
    -0.0033100002899363857, -0.0033512270983823019, -0.0033463809272745977, 
    -0.0033001183375122008, -0.0032183382081071715, -0.00310780587218926, 
    -0.0029757478814200133, -0.0028294836107071535, -0.0026761135317479199, 
    -0.0025222648684962864, -0.0023738830662715081, -0.0022360556506701209, 
    -0.0021128669030504722, -0.0020072954504378403, -0.0019211607503523351, 
    -0.0018551387744293484, -0.0018088255317460029, -0.0017808882135976526, 
    -0.0017692794264155493, -0.0017714993097236779, -0.0017848247171578895, 
    -0.0018064854306462125, -0.0018337418331480593, -0.0018638692089680759, 
    -0.0018940933679818302, -0.0019215065753060553, -0.0019430265228774835, 
    -0.0019554270671128006, -0.0019554896912017936, -0.0019402467403112334, 
    -0.0019072774090079661, -0.0018549868305565019, -0.0017828165046100512, 
    -0.0016913361964006281, -0.001582252709441644, -0.0014583480255445282, 
    -0.0013233844279505653, -0.0011819491913075109, -0.0010391896860610947, 
    -0.00090040264849832125, -0.00077046360266758433, 
    -0.00065315525557884551, -0.00055050466825364117, -0.0004622421802786919, 
    -0.00038550218952128432, -0.00031484920067281384, 
    -0.00024266289042896834, -0.00015985384792861491, 
    -5.6865242986928557e-05, 7.5142741161783578e-05, 0.00024305732069344996, 
    0.00045066160732585138, 0.00069772915742710262, 0.00097949360128512727, 
    0.0012866074077823903, 0.0016056545000073693, 0.0019201772689010608, 
    0.0022121528178168075, 0.002463730856142939, 0.0026590281665754265, 
    0.0027857450794696501, 0.0028363636238947594, 0.0028087800289037842, 
    0.0027062743434340237, 0.002536866580048478, 0.0023121565361893105, 
    0.0020458726801231915, 0.0017523535402491814, 0.0014451821775059903, 
    0.001136171994253615, 0.00083480657175329163, 0.00054815533714327807, 
    0.00028121411160347446, 3.7527391325019706e-05, -0.00018005778750916868, 
    -0.00036872256503422463, -0.00052522770872625918, 
    -0.00064580166598476809, -0.00072639966159804325, 
    -0.00076328971121956404, -0.00075384926875865824, 
    -0.00069741171920000705, -0.0005959627653384608, -0.00045455170960274704, 
    -0.00028126794912600877, -8.6799440124278934e-05, 0.00011639895790564842, 
    0.000315206721060334, 0.00049702150844739914, 0.00065087808860914381, 
    0.00076834235734719815, 0.00084412178145529433, 0.00087632780698458624, 
    0.00086643978468250603, 0.00081899686427378362, 0.00074108842106951117, 
    0.00064169349071467065, 0.00053091109836923833, 0.00041912228856398235, 
    0.00031613503408958087, 0.00023036272079075427, 0.0001681064567304244, 
    0.00013301769969398288, 0.00012583035216218191, 0.00014442724620460185, 
    0.00018424748452543368, 0.00023898567279171713, 0.00030145463166812454, 
    0.00036440958598890931, 0.00042119427336885149, 0.00046612058220068831, 
    0.00049457910130655059, 0.00050298966303747921, 0.00048868771413636649, 
    0.00044988377545987707, 0.00038574633825015593, 0.00029662400507564097, 
    0.00018433591233523266, 5.2419407636429387e-05, -9.3815557457136057e-05, 
    -0.00024750398400937891, -0.0004007549809637967, -0.00054540452512474825, 
    -0.00067388196923082741, -0.00077998341598046366, 
    -0.00085941860253207244, -0.00091002899829588509, 
    -0.00093165835960001787, -0.00092573364084397986, 
    -0.00089469818643840712, -0.00084140990052925186, 
    -0.00076861261700739082, -0.00067859538508755184, 
    -0.00057306895297711447, -0.00045327742017739221, 
    -0.00032030068348227591, -0.00017548733001733193, 
    -2.0905288371930817e-05, 0.00014028789292581728, 0.00030364845636424555, 
    0.00046345069122746401, 0.00061294964220104777, 0.00074483436291420562, 
    0.00085186298510123919, 0.0009275768365490523, 0.00096699757589586988, 
    0.00096719984388164986, 0.00092764296845685964, 0.0008502077754963277, 
    0.00073891498500137237, 0.00059940187099658709, 0.00043825163623234888, 
    0.00026228743883632187, 7.7962194461420365e-05, -0.00010908279516594589, 
    -0.00029423681057431456, -0.00047392968669098532, -0.0006454981912945041, 
    -0.00080697841109444134, -0.0009569143112950272, -0.0010942208926803425, 
    -0.0012181303193366212, -0.001328228897521261, -0.0014245539529478455, 
    -0.0015077121730033829, -0.0015789359489493189, -0.0016400042621278553, 
    -0.0016930133562332698, -0.0017399965730861369, -0.0017824978341798216, 
    -0.0018211987357206968, -0.0018556659426500371, -0.0018843248010693156, 
    -0.0019046383455858051, -0.0019134902271945281, -0.0019076884693245474, 
    -0.0018845114230696849, -0.0018421979108462802, -0.0017803042922226466, 
    -0.0016998635202126432, -0.0016033403746435794, -0.0014943811960969372, 
    -0.0013774426489294167, -0.0012573713496964159, -0.0011390229384803194, 
    -0.0010269669814151694, -0.00092527619630694341, -0.00083739167623555545, 
    -0.00076601302918344089, -0.00071298905786627734, 
    -0.00067920637387973892, -0.00066448928259089631, 
    -0.00066755902124558837, -0.00068606726591612728, 
    -0.00071677705765685784, -0.00075585000835338197, 
    -0.00079924678040388169, -0.00084318643535924681, 
    -0.00088457148569469259, -0.00092133560938093895, 
    -0.00095260091850077723, -0.00097862388188501149, -0.0010004971441562765, 
    -0.0010196756482702745, -0.0010374255086098979, -0.0010543192028873321, 
    -0.0010699283878113886, -0.0010827945613219665, -0.001090691089763879, 
    -0.0010910932618410961, -0.001081733893916271, -0.0010610877478113214, 
    -0.0010286910873066012, -0.00098527988536864074, -0.00093275249826353743, 
    -0.00087404486299593419, -0.00081292708658541653, 
    -0.00075378365119279863, -0.00070136084770413068, 
    -0.00066051300148052441, -0.00063596495704739938, 
    -0.00063209846104606709, -0.00065273922384268815, 
    -0.00070091102953359879, -0.00077853772039161999, 
    -0.00088612372439901142, -0.0010224638777762108, -0.0011844603861110058, 
    -0.0013671282445580748, -0.0015638260345989022, -0.0017667175263424764, 
    -0.0019673852086658258, -0.0021575174956697373, -0.0023295433614250491, 
    -0.0024771450455601256, -0.0025955904418654228, -0.0026818699570346043, 
    -0.0027346857423656418, -0.0027543064512783083, -0.0027423554795660264, 
    -0.0027015396257670616, -0.0026353661806387992, -0.0025478679243655842, 
    -0.0024433757961665847, -0.0023263492200351803, -0.0022013031731909953, 
    -0.0020727771640627907, -0.0019453637675222414, -0.0018236939165360126, 
    -0.001712364114842549, -0.0016157634967241892, -0.0015377982581905748, 
    -0.001481561123554918, -0.0014490010712957433, -0.0014406388044648237, 
    -0.0014554138757472046, -0.0014906538327679394, -0.0015421948382844087, 
    -0.0016046263645573011, -0.0016716643112573649, -0.001736602359303454, 
    -0.0017928494376780726, -0.0018345031212096915, -0.0018569268331757841, 
    -0.0018572672009707551, -0.0018348455578740379, -0.0017913538114126622, 
    -0.0017307817584971009, -0.0016590731911256642, -0.001583510023669168, 
    -0.0015119127852477429, -0.0014517398689712459, -0.0014092271896213443, 
    -0.0013886638740904947, -0.0013919101696386188, -0.0014182124801547539, 
    -0.0014643324097690612, -0.0015249948229812873, -0.0015935628493984558, 
    -0.0016628460574022326, -0.001725912331317354, -0.001776772797159702, 
    -0.0018108481171708725, -0.0018251472758829843, -0.0018181781238110943, 
    -0.0017896295632855237, -0.0017399214115014882, -0.0016697454868743111, 
    -0.0015797064467993032, -0.0014701474309424178, -0.0013411970299318184, 
    -0.0011930134733477862, -0.0010261945203314574, -0.00084222842486065077, 
    -0.00064390254330146698, -0.00043554543671898093, 
    -0.00022302247946845251, -1.3444556644196871e-05, 0.0001853786602099892, 
    0.00036564974104632403, 0.00052033561360358127, 0.00064382310570485803, 
    0.00073236772059108858, 0.0007842706775049058, 0.00079978890802002967, 
    0.0007808303025750549, 0.00073051651759925671, 0.00065272072427698493, 
    0.00055164778984670535, 0.00043152018169235291, 0.00029639302063639357, 
    0.00015007303582356641, -3.8942127990561001e-06, -0.00016219816719035209, 
    -0.00032174731842775454, -0.00047969682270508705, 
    -0.00063352859854884066, -0.00078118698631991475, 
    -0.00092125242605957066, -0.0010530995508142987, -0.0011769953809915466, 
    -0.0012940931826149185, -0.0014062855353277853, -0.0015159336381128576, 
    -0.0016254832212657265, -0.0017370231136903031, -0.0018518631180816998, 
    -0.0019701909747242632, -0.002090880303888939, -0.0022114873666839244, 
    -0.0023284438460603359, -0.0024374381995350899, -0.0025339511409016263, 
    -0.0026138348144590954, -0.0026738849598622527, -0.0027122867733838721, 
    -0.0027288609563297125, -0.0027250960282763407, -0.0027039393499504764, 
    -0.002669421485240419, -0.0026261729269236598, -0.0025789091955532154, 
    -0.0025319676599086789, -0.0024889539890951781, -0.0024525482958330548, 
    -0.0024244808216150522, -0.0024056658252364846, -0.0023964277613096512, 
    -0.0023967618885945446, -0.0024065317406038633, -0.0024255833179149177, 
    -0.0024536710385207176, -0.0024902559882511361, -0.0025341219315467259, 
    -0.0025829448418897179, -0.0026329042792941669, -0.0026784674808253126, 
    -0.0027124596888770365, -0.0027264523807141146, -0.0027114465811933896, 
    -0.0026587316353606713, -0.002560815441085656, -0.0024122287674860519, 
    -0.002210087410874504, -0.0019543302841681228, -0.0016476479897366133, 
    -0.0012951849748657868, -0.00090410164397854013, -0.00048311401952846325, 
    -4.2047605799789645e-05, 0.00040857489931881422, 0.00085793774637410675, 
    0.0012953345128916571, 0.001710558156205869, 0.0020942685752287555, 
    0.0024383011004492426, 0.0027359037315349169, 0.0029818798636837636, 
    0.0031726436672162872, 0.0033062050091387241, 0.0033820760157820462, 
    0.0034011357949660348, 0.0033654414734380902, 0.003278039722775075, 
    0.0031427497185000011, 0.0029639921520239515, 0.0027466505637233959, 
    0.0024959950085808348, 0.0022176668636487364, 0.0019176583703385403, 
    0.0016022711924358949, 0.0012780081914641598, 0.00095138820919295642, 
    0.00062873874868886155, 0.00031599379364554244, 1.8521739085201102e-05, 
    -0.0002589987774643322, -0.00051266639393798418, -0.00073942683674585658, 
    -0.00093715339953487809, -0.0011047327581066991, -0.0012421930858623844, 
    -0.0013508456997995315, -0.001433406371147268, -0.0014940155896012652, 
    -0.0015381176257039972, -0.001572155551892847, -0.0016030767835056949, 
    -0.0016377232188658965, -0.0016821691891791071, -0.0017410848485352385, 
    -0.0018172209923015808, -0.0019110390596137113, -0.0020205396330191298, 
    -0.002141284847864377, -0.002266635707456101, -0.0023881871673110252, 
    -0.0024964331268667412, -0.0025816056565286325, -0.00263465969904277, 
    -0.0026482922520976652, -0.0026178579162120016, -0.0025420735220876055, 
    -0.0024233694180646618, -0.0022678198708368032, -0.0020846064017387114, 
    -0.0018850893677232294, -0.0016816343052208544, -0.0014863889824055956, 
    -0.0013102090747802706, -0.0011618735820643628, -0.0010476153922048307, 
    -0.0009709817669156009, -0.00093294951869797018, -0.00093230415821050937, 
    -0.00096614375524273427, -0.0010304891867532915, -0.0011208772888758954, 
    -0.0012328386374199764, -0.0013621585202539688, -0.0015049347337757583, 
    -0.0016574340265280761, -0.0018158553013521545, -0.0019760635317215337, 
    -0.0021333742741985857, -0.0022824293554227549, -0.0024172054411144175, 
    -0.0025311604030913161, -0.0026175217670292034, -0.0026697018259269644, 
    -0.0026817891337037429, -0.0026490771561312868, -0.0025685448745167631, 
    -0.0024392564014015898, -0.002262599242204543, -0.0020423440170479128, 
    -0.0017845088719388711, -0.0014970409667195948, -0.0011893662293444248, 
    -0.00087187098788296744, -0.00055537001215354262, 
    -0.00025061115216619336, 3.2139857520223488e-05, 0.00028341227645829921, 
    0.00049473059277373166, 0.00065873032499378899, 0.00076918175241323054, 
    0.00082100646859768756, 0.00081030451709785322, 0.00073449007613493459, 
    0.00059254433084361734, 0.00038537611352615255, 0.00011624627820046765, 
    -0.0002088460034369394, -0.00058090980921967424, -0.00098793192936452007, 
    -0.0014151342666522419, -0.0018455387293890202, -0.0022608617756068572, 
    -0.0026426667790043789, -0.0029736859646338769, -0.0032391944217885008, 
    -0.0034282297181682073, -0.003534561674729726, -0.0035572312405457119, 
    -0.0035005877461521998, -0.0033738188373524203, -0.0031900047563704205, 
    -0.002964823040074482, -0.0027150794928729335, -0.002457238413004938, 
    -0.0022061018562461758, -0.0019737633787513613, -0.001768876836693528, 
    -0.0015962509269858501, -0.0014567737429805546, -0.0013476717764734224, 
    -0.0012631138933090645, -0.0011951622007938848, -0.0011349878082310551, 
    -0.0010741926924821715, -0.0010060438287552145, -0.00092642713808965783, 
    -0.00083441015290582152, -0.00073240611044433652, -0.0006259361771763514, 
    -0.00052307278365925941, -0.00043366106528103091, 
    -0.00036830884238404969, -0.00033728319840095096, 
    -0.00034933549581571578, -0.00041058490358096518, 
    -0.00052357992605322709, -0.00068667985321192628, 
    -0.00089388194521168476, -0.0011351484213418062, -0.001397234236866053, 
    -0.0016649323741540661, -0.0019225689881436528, -0.0021555542028040813, 
    -0.0023517554972702537, -0.0025025204614815433, -0.0026032079080502389, 
    -0.0026532085229256184, -0.0026554686125539084, -0.0026156873404244957, 
    -0.0025413419947570241, -0.002440754714125728, -0.0023223727051689372, 
    -0.0021943610552246228, -0.0020644844623913224, -0.0019402041811155987, 
    -0.0018288182009402539, -0.0017375226415832414, -0.0016733009386281075, 
    -0.001642649659824878, -0.0016511408344850706, -0.0017029373726714331, 
    -0.0018003202324476445, -0.0019432919864092154, -0.0021293350851801012, 
    -0.0023533499830883315, -0.0026077869227546522, -0.0028830175134550487, 
    -0.0031678988126767286, -0.0034505402226560995, -0.0037191399434554212, 
    -0.0039627825360529674, -0.0041720917684649663, -0.0043396076988272518, 
    -0.0044599029633945464, -0.0045294483567594832, -0.0045463532915026002, 
    -0.0045100368974018961, -0.0044209323111167043, -0.004280270259644431, 
    -0.0040899383048954661, -0.003852452099806307, -0.0035709835827521844, 
    -0.0032494791341936119, -0.0028928329320779354, -0.0025070747298544306, 
    -0.0020995318470996781, -0.0016789238536144703, -0.0012553095398960916, 
    -0.00083988538550314369, -0.00044456342708194753, 
    -8.1390452505882325e-05, 0.000238227877499896, 0.00050437289467351138, 
    0.00070950894647107206, 0.00084926204949485856, 0.00092304270661088688, 
    0.00093434416339252698, 0.0008907050956560085, 0.00080325310040559885, 
    0.00068585520125892692, 0.0005539778811495743, 0.00042334004290688233, 
    0.00030852812371951827, 0.00022172055225768285, 0.00017164887314037147, 
    0.00016291251101023226, 0.00019571901381867961, 0.00026605346617516524, 
    0.00036625279050352382, 0.00048590646036104321, 0.00061299638515406076, 
    0.00073515715715696925, 0.00084098720688276338, 0.00092125674561332528, 
    0.00096995208046218504, 0.0009850359214334547, 0.0009688357134379369, 
    0.00092798079573102308, 0.00087283397596599232, 0.00081644581088494096, 
    0.00077308164201799487, 0.00075650940290641899, 0.00077826642901830038, 
    0.00084613246430382627, 0.00096305690153584696, 0.0011266895961189955, 
    0.0013295372557944993, 0.0015597041524696657, 0.0018021128083591735, 
    0.0020400134075497151, 0.00225660206169028, 0.0024365646752163741, 
    0.0025673928367584489, 0.0026403146394424733, 0.0026507828144466121, 
    0.0025984906625107188, 0.00248696969840791, 0.0023228499018275771, 
    0.0021149271659604775, 0.0018732032889984596, 0.0016080607154757721, 
    0.0013296740808335821, 0.0010477056845391206, 0.00077123201944790266, 
    0.0005088178894440598, 0.0002686785188338363, 5.8791830740165284e-05, 
    -0.00011307019182000966, -0.00023943551812517322, 
    -0.00031334444833185473, -0.00032869761638635832, -0.0002806835992626194, 
    -0.00016627616865871298, 1.5300274799248426e-05, 0.000262179576598629, 
    0.00056964938676566581, 0.00093018836877934363, 0.001333746628214245, 
    0.0017682730404393759, 0.002220357079543172, 0.0026759076150842317, 
    0.0031207384966049205, 0.0035409831987887525, 0.0039233163328599076, 
    0.0042550395772215964, 0.004524116443778657, 0.0047192806743795914, 
    0.0048302890964620308, 0.004848360240811843, 0.00476676749346384, 
    0.0045815011550854262, 0.0042918992578726348, 0.0039011141904201655, 
    0.0034163464469845837, 0.0028487468555924364, 0.002212996852855247, 
    0.0015265206981813417, 0.0008084181229919236, 7.8203236601265432e-05, 
    -0.0006454906543838547, -0.0013460806455909977, -0.0020099216494625254, 
    -0.0026268346038670681, -0.0031902288029900744, -0.0036968819092121044, 
    -0.0041464217281914351, -0.0045406646405445642, -0.0048828682182164547, 
    -0.0051770123130864421, -0.0054272012871988268, -0.0056372127500792634, 
    -0.0058102199752145854, -0.0059487052744034126, -0.0060545282303919069, 
    -0.0061290893557510153, -0.0061735566618916961, -0.0061890712963741032, 
    -0.0061769069637718629, -0.0061385566232822252, -0.0060757466195631854, 
    -0.005990409131702944, -0.00588462685356926, -0.0057605679677158305, 
    -0.0056204965496032978, -0.0054668153073021992, -0.0053021927052949039, 
    -0.005129694613783385, -0.0049528720196172328, -0.0047757686999607887, 
    -0.0046027935379007942, -0.0044384760537781306, -0.0042871180753070205, 
    -0.0041523907952492377, -0.0040369359355602171, -0.0039420221486310709, 
    -0.0038673385809402882, -0.003810928397519296, -0.0037693177044529798, 
    -0.003737792732656166, -0.0037108103669585674, -0.003682510219884996, 
    -0.0036472778423618539, -0.003600267548364483, -0.0035378812918823153, 
    -0.0034581033359251672, -0.0033606539867734593, -0.0032469492925421002, 
    -0.0031198409252852608, -0.0029832004584744885, -0.0028413722398037324, 
    -0.0026986065289262904, -0.0025585415373066997, -0.0024238051120834981, 
    -0.0022957980701008617, -0.0021746934132662443, -0.0020596063118035186, 
    -0.0019489287478980698, -0.0018407408014448187, -0.0017332596240013025, 
    -0.0016252292475162832, -0.00151622736215618, -0.0014067863791452867, 
    -0.001298310180289197, -0.0011927069587598794, -0.0010917978723589232, 
    -0.00099656881582127206, -0.00090639830995384112, 
    -0.00081846536233659269, -0.00072747921476468743, 
    -0.00062586319428005184, -0.00050441995906553173, 
    -0.00035341409870780135, -0.00016390257025760194, 7.0856917482539053e-05, 
    0.00035415623385053573, 0.00068491326569807042, 0.0010572419989436522, 
    0.0014605893255516767, 0.0018804388265402947, 0.002299508611674877, 
    0.0026992793729595003, 0.0030617055871323424, 0.0033708944570418251, 
    0.0036145498148863926, 0.0037850408296028655, 0.0038799485431731161, 
    0.003902034374576274, 0.0038586425555334198, 0.0037606621857236566, 
    0.0036212029330724032, 0.0034542008739631568, 0.003273123367165268, 
    0.0030898922316000936, 0.0029141116690483285, 0.0027526250791700306, 
    0.0026094465654934638, 0.0024860082681207088, 0.0023816727630588917, 
    0.0022943999467478567, 0.0022214236606909956, 0.0021598780424426488, 
    0.0021073219080546667, 0.0020621395136813008, 0.002023832406812474, 
    0.0019931944466883298, 0.0019723315777738729, 0.0019645024837214595, 
    0.0019737363996947576, 0.0020042592265494498, 0.0020597712647721423, 
    0.0021426603659492473, 0.0022532649041249464, 0.0023893355361396321, 
    0.0025457333984655042, 0.0027144784695487438, 0.00288516426948508, 
    0.0030457392068114508, 0.0031835674969179083, 0.0032866798189528346, 
    0.0033450521507309679, 0.003351724404870532, 0.0033036217526220277, 
    0.0032019504766698827, 0.0030521254257855407, 0.0028632701224714937, 
    0.0026473597887756513, 0.0024181004673235699, 0.0021897175128801445, 
    0.0019757788925613474, 0.0017882156833226, 0.0016365659717734247, 
    0.0015275352821282752, 0.0014648016536471433, 0.0014490880954482514, 
    0.0014784205569827093, 0.0015485757994337505, 0.001653635619466888, 
    0.0017865469134502271, 0.0019396471595902608, 0.002105054336203731, 
    0.0022749074865543329, 0.0024414394846962589, 0.0025969144893120311, 
    0.0027334838368471624, 0.0028430583323175774, 0.0029173005773350303, 
    0.002947831012033989, 0.0029267018140771445, 0.0028470385286349081, 
    0.002703819794066377, 0.0024945947504336641, 0.0022200396080236016, 
    0.0018842623505193842, 0.0014947665447382805, 0.0010621019429783479, 
    0.00059922346319410836, 0.00012060853337986952, -0.00035874369768996252, 
    -0.00082433184740832307, -0.0012630851817435318, -0.0016641030617757812, 
    -0.002019064807416713, -0.002322294568506994, -0.0025704438039260303, 
    -0.0027618795801169667, -0.0028958777163156043, -0.0029718324929129099, 
    -0.0029886417285973719, -0.002944418136878547, -0.0028365466113649705, 
    -0.002662100076559358, -0.0024184953479224102, -0.0021042710107964718, 
    -0.0017198449944954867, -0.0012681386705919809, -0.00075497491413197438, 
    -0.00018923135364503827, 0.00041724572372721814, 0.0010499620648348482, 
    0.001692247952141101, 0.002325896058307349, 0.0029319458354804592, 
    0.0034916121387151521, 0.0039873214834957836, 0.0044038140517885654, 
    0.0047292477312150492, 0.0049561477192043525, 0.0050820972076323972, 
    0.005110060602458685, 0.0050482760646416375, 0.0049096892290444545, 
    0.0047109752566441825, 0.0044712082226162509, 0.0042102902715765176, 
    0.0039473077510928118, 0.0036989558518346647, 0.0034782701030965655, 
    0.0032937379945452523, 0.0031489303865542802, 0.0030425574003936874, 
    0.0029690520941709465, 0.002919477057577731, 0.0028827654077371368, 
    0.0028470978769636816, 0.0028012560579106769, 0.0027357953791229128, 
    0.002643892147628577, 0.0025218166851060648, 0.0023690046025762346, 
    0.002187790246512653, 0.0019829129971739314, 0.0017608964728106856, 
    0.0015293926525645483, 0.0012965836387313712, 0.0010706696362680112, 
    0.00085947924517954476, 0.0006701902312763791, 0.0005091748760758457, 
    0.00038192818411028639, 0.00029305012199541377, 0.00024619743436761759, 
    0.00024394397390611568, 0.00028752853602102016, 0.00037648045989546069, 
    0.00050821934068371027, 0.00067766731703332783, 0.00087708054865184523, 
    0.001096161563368774, 0.0013225867951899347, 0.0015428769276298584, 
    0.00174357711711383, 0.0019125800916128081, 0.002040366303959003, 
    0.0021209747069961893, 0.0021525564101769531, 0.0021373212990926597, 
    0.0020809359306883228, 0.0019914033091558794, 0.0018776055642931507, 
    0.0017477521557177334, 0.0016080054454370924, 0.0014615107260831154, 
    0.0013080566023935087, 0.001144418138338847, 0.00096537735324799727, 
    0.00076519024259796094, 0.0005392458959248399, 0.00028557462750241719, 
    5.9273596221756522e-06, -0.00029374406777118208, -0.00060346250315652873, 
    -0.0009100017430963849, -0.0011981195075229537, -0.0014520681095130093, 
    -0.0016571780085343909, -0.0018013145207899592, -0.0018760403227413825, 
    -0.0018773627060076057, -0.0018060023395712931, -0.0016671679110765445, 
    -0.0014699118904502009, -0.0012261406085673722, -0.00094940312742221929, 
    -0.00065362425972011889, -0.00035191635182559402, 
    -5.5586962493713358e-05, 0.00022650163084838345, 0.00048820276181629887, 
    0.00072596020842287845, 0.00093837679339967006, 0.0011256198548512866, 
    0.0012887979614281681, 0.0014294793327941601, 0.0015494012135396334, 
    0.001650357256283967, 0.001734085802445783, 0.0018020995582458553, 
    0.0018553389049813644, 0.0018938125969042267, 0.0019163514440536631, 
    0.0019207213440349579, 0.0019042166647987805, 0.0018646272902184155, 
    0.0018012490582312829, 0.0017155235275213346, 0.0016109324549325836, 
    0.0014921578025364325, 0.0013637818514203165, 0.0012290305652110612, 
    0.0010889620751868456, 0.0009423194510170224, 0.00078605628242302034, 
    0.0006163452239641566, 0.00042993806507962869, 0.00022558380251322396, 
    5.2755761580831634e-06, -0.00022491965569548626, -0.00045465990541546466, 
    -0.00066979962970028085, -0.00085354941763933208, 
    -0.00098811515624611795, -0.0010565319408767111, -0.0010445050155193912, 
    -0.00094205423380340589, -0.00074482780944576312, 
    -0.00045496981782525549, -8.141526843639035e-05, 0.00036046416950040894, 
    0.00084993686638962197, 0.0013626094407905793, 0.0018725490294255903, 
    0.0023545193641276657, 0.0027860216342566763, 0.0031488347533585891, 
    0.003429966616411042, 0.0036219642194565017, 0.0037226738519205694, 
    0.003734604006367691, 0.0036640678185178317, 0.0035202132226997912, 
    0.0033140575080513788, 0.0030575687301868746, 0.0027627712011114559, 
    0.0024409430952701057, 0.0021019189607002905, 0.0017536075675956512, 
    0.001401801599871964, 0.0010502673332483171, 0.00070111792855402167, 
    0.00035541467097277156, 1.3891113677144649e-05, -0.00032231060105553246, 
    -0.00065099116861713985, -0.00096847620995168951, -0.0012694617763867873, 
    -0.0015472440146380758, -0.0017943323503246747, -0.0020034646713931038, 
    -0.0021688996308641961, -0.0022877562980154606, -0.0023611401061612593, 
    -0.0023947684069264437, -0.0023989395124386836, -0.0023877832890517301, 
    -0.0023778624520449268, -0.0023863244195299121, -0.0024288031679338276, 
    -0.0025173877267368142, -0.0026588928966957562, -0.00285364502716005, 
    -0.0030950110161942742, -0.0033696989151220528, -0.0036588638406944854, 
    -0.0039398885018497214, -0.0041886720902329488, -0.0043820968946034671, 
    -0.0045003569163031762, -0.0045288886586664122, -0.0044595830443638282, 
    -0.0042912038115336471, -0.0040290493866291617, -0.0036839514117876044, 
    -0.0032708180976240703, -0.0028069235430945609, -0.0023101097727195275, 
    -0.001797182979451093, -0.001282698578210851, -0.00077841311557239642, 
    -0.00029346956597433319, 0.00016479907251797579, 0.00058972960206696106, 
    0.00097442263107893278, 0.0013113256983798408, 0.0015925384789958561, 
    0.0018106615073415987, 0.001959905667799005, 0.0020372251081585565, 
    0.0020432665609239967, 0.0019830885330516254, 0.001866506392009452, 
    0.0017079262872915604, 0.0015255234549856457, 0.0013397898352167004, 
    0.0011715619563384917, 0.0010397557665861904, 0.00095923879709569073, 
    0.00093907110966853606, 0.00098144478522763849, 0.0010814316475505361, 
    0.0012275775553681318, 0.0014032518165695042, 0.0015886050982681576, 
    0.001762871850457582, 0.001906739840100644, 0.0020045137523140777, 
    0.0020458098812288, 0.0020265445366717916, 0.0019491673975955341, 
    0.0018220507767293549, 0.0016581506710954695, 0.0014730692151175982, 
    0.0012828146535578597, 0.0011016085132615691, 0.00093998329027916781, 
    0.0008034640630980893, 0.00069198365031127767, 0.00060005793808882025, 
    0.00051764651277047774, 0.00043154362650775762, 0.00032710567573035942, 
    0.00019011581282843274, 8.5259422804545679e-06, -0.00022605660056915135, 
    -0.00051741154919782888, -0.00086432385593102805, -0.0012608633953656747, 
    -0.0016972487927891515, -0.002161084487796758, -0.0026387773882667188, 
    -0.0031168683978010782, -0.0035830637232838369, -0.0040268159259754695, 
    -0.0044394294052933049, -0.0048136761936647928, -0.0051431260359772303, 
    -0.0054214346755987863, -0.0056418096155166249, -0.0057968146294921684, 
    -0.005878653039511272, -0.0058799383314612225, -0.005794756276395056, 
    -0.0056199524780244986, -0.005356369828396549, -0.0050097694234902358, 
    -0.0045913214047527649, -0.0041175225223245484, -0.0036094694087516728, 
    -0.0030915901620416531, -0.002589922464951717, -0.0021300823398255416, 
    -0.0017351468285417785, -0.0014236870301409619, -0.0012081132916437532, 
    -0.0010935777986243117, -0.0010775608113055047, -0.0011502800536903072, 
    -0.0012958832455469797, -0.0014943714788904603, -0.0017238303924598099, 
    -0.0019626980795926221, -0.0021917779177650478, -0.0023957618103546065, 
    -0.002564285299237635, -0.0026925439896240549, -0.0027814161511214262, 
    -0.0028371398136989401, -0.0028704551169119116, -0.0028952148055171089, 
    -0.0029265974041036338, -0.0029791356459266437, -0.0030648335436489855, 
    -0.0031915900653779446, -0.0033621174673948264, -0.003573422568686614, 
    -0.0038169282845191368, -0.0040792188060093278, -0.0043433885698244273, 
    -0.0045909329411253251, -0.0048039452228210485, -0.0049674378847608096, 
    -0.0050713690766234307, -0.0051120854323720606, -0.0050928703891859163, 
    -0.0050234941642526452, -0.0049187615258497741, -0.0047965108801514347, 
    -0.004675264904285009, -0.0045721026706259842, -0.0045009789896069199, 
    -0.0044716183404343666, -0.0044890311477416289, -0.0045535883873396056, 
    -0.0046616131742246479, -0.0048062956589976389, -0.0049788171097432717, 
    -0.0051695400516438093, -0.0053690046098562498, -0.0055686292821195702, 
    -0.0057610494346046629, -0.0059401146970719564, -0.0061006894632949383, 
    -0.0062383637811638274, -0.0063492488940119531, -0.0064298355726747332, 
    -0.0064769217943722313, -0.0064876583686063393, -0.0064596544499140873, 
    -0.006391184580745831, -0.0062814560589701564, -0.006130917170097879, 
    -0.00594147520328477, -0.0057166431499188191, -0.0054616135617002832, 
    -0.0051832614222870679, -0.0048902077337163686, -0.004592867341495519, 
    -0.0043034171939729882, -0.0040355449857779144, -0.0038038742482880785, 
    -0.0036230409413100825, -0.0035064410781615379, -0.0034648567818646452, 
    -0.0035050766608837693, -0.0036287825655997078, -0.0038318873169415186, 
    -0.0041044686723843366, -0.0044314405736399221, -0.0047938724985055609, 
    -0.0051708139884582682, -0.0055414616007292061, -0.0058873044764230368, 
    -0.006193982828077634, -0.0064524970371700801, -0.0066596174158854594, 
    -0.0068175350740404409, -0.0069328499960161858, -0.0070152772455940029, 
    -0.007076219044048768, -0.0071274551004635069, -0.0071800241036461421, 
    -0.0072432441882583718, -0.0073239803114950319, -0.0074260150551317839, 
    -0.0075496851101485565, -0.0076917318396123348, -0.0078454743888643451, 
    -0.0080013175540960668, -0.0081475017556894673, -0.0082711199769531663, 
    -0.0083592382942304037, -0.0084000362929542386, -0.0083839033102018467, 
    -0.00830431551142247, -0.0081584347222474832, -0.0079472696065953814, 
    -0.007675429960718929, -0.007350432965809308, -0.0069817354031802299, 
    -0.0065795704160825485, -0.0061538658994329904, -0.0057133867531656592, 
    -0.0052651603985535058, -0.0048143118324390976, -0.0043642161477739942, 
    -0.0039169146786317069, -0.0034736398525486607, -0.0030352633124551111, 
    -0.002602465647757925, -0.0021757268061038289, -0.0017550453617029122, 
    -0.0013396465131159383, -0.00092784659086928771, -0.0005171113425569882, 
    -0.00010437212372386761, 0.00031354009730465192, 0.00073962022352968616, 
    0.0011765168058451509, 0.0016266608603850599, 0.0020924529338488141, 
    0.0025764203132525336, 0.0030812821222386774, 0.0036097507388502823, 
    0.0041642607761972353, 0.0047464563491132041, 0.0053566205974407309, 
    0.0059930731399928444, 0.0066517149359437552, 0.0073257341307047816, 
    0.0080057181580207373, 0.0086800400289531107, 0.0093355481283225808, 
    0.0099582601818367211, 0.010534120518728306, 0.011049562765603337, 
    0.01149192167435672, 0.011849744708049864, 0.012112978876878882, 
    0.012273138663730384, 0.012323504662711949, 0.012259326908096151, 
    0.012078094202699268, 0.011779751726690293, 0.011366909504691639, 
    0.010844946154968841, 0.010221909282713057, 0.0095083176323480009, 
    0.0087166587165712281, 0.0078608121533246186, 0.0069554244484763134, 
    0.0060153929834617917, 0.0050555350135326332, 0.0040905725676796305, 
    0.0031352270738365501, 0.0022044444528272642, 0.0013135323251960362, 
    0.00047807089512114933, -0.0002865179706965678, -0.00096566947776918007, 
    -0.0015466399070709715, -0.0020195329994534168, -0.0023782588251844675, 
    -0.0026211496310813241, -0.002751146683424978, -0.002775451890244811, 
    -0.0027047449423249778, -0.0025521052730894996, -0.002331957692555934, 
    -0.002059231791385353, -0.001748846398698667, -0.0014155335089563411, 
    -0.0010737894236996415, -0.00073789835655749638, -0.00042172419225817851, 
    -0.00013828197643652427, 0.00010099951535579802, 0.00028717879823669259, 
    0.00041475362516421935, 0.00048245997688846224, 0.00049368629760923339, 
    0.00045632681860347142, 0.00038208549894454985, 0.00028510871820207253, 
    0.0001802554437846291, 8.1260998493898774e-05, -7.3446044398335283e-07, 
    -5.8146125801267646e-05, -8.714987227715883e-05, -8.7304456672939986e-05, 
    -6.0902649904792791e-05, -1.2041050490687981e-05, 5.4229479543125734e-05, 
    0.00013281886876022721, 0.00021950576169134416, 0.00031175784688493172, 
    0.00040943143457738669, 0.00051511299121031768, 0.00063388426399649104, 
    0.00077248853281552238, 0.00093770874728588312, 0.0011345416487885424, 
    0.0013642688772665108, 0.0016231995387992306, 0.0019023055504041129, 
    0.0021878563550757789, 0.0024627591035495189, 0.0027081864852665431, 
    0.0029049579677001363, 0.0030344849827007659, 0.0030797135189793278, 
    0.0030261385753733681, 0.0028633140803626615, 0.0025861743535881667, 
    0.002195524333430269, 0.0016974654990012453, 0.0011020760286971421, 
    0.00042189060836173888, -0.00032935038307849748, -0.001137416539757016, 
    -0.0019877499357714569, -0.0028652502093296645, -0.0037540062454592101, 
    -0.0046370995484537134, -0.0054968856681673929, -0.0063155696075437584, 
    -0.007076045706531052, -0.0077629899423176689, -0.0083640180361694207, 
    -0.0088708600359153449, -0.0092802561095208357, -0.0095943229921964766, 
    -0.009820360596783026, -0.009969878502089892, -0.010057160022020046, 
    -0.010097326993592351, -0.010104425108275724, -0.010089505733331467, 
    -0.010059207662175867, -0.010014879008428627, -0.0099522728490322176, 
    -0.009861810149925182, -0.0097291677106717059, -0.0095360773566018457, 
    -0.0092614596634470834, -0.0088829359812869716, -0.0083789771442097909, 
    -0.0077314158743932368, -0.0069281876510568288, -0.0059656480108906743, 
    -0.0048501432722360639, -0.003598280452257567, -0.0022361904182518553, 
    -0.00079784787643493165, 0.00067684266085289203, 0.0021440921453772374, 
    0.0035580953736812182, 0.0048729555801277948, 0.0060447856859054848, 
    0.0070344518550942061, 0.0078101052521164817, 0.0083497244383635844, 
    0.0086429240295183042, 0.0086918664918662052, 0.0085109511088369647, 
    0.0081255378958326324, 0.0075697903264383207, 0.0068838735170938005, 
    0.0061111707897776512, 0.0052956933785971699, 0.0044798145790487728, 
    0.0037026481812431344, 0.0029988845900606209, 0.0023981134186671577, 
    0.0019244662111709463, 0.0015964724499030367, 0.0014267567383784694, 
    0.0014214686868704051, 0.001579657691215926, 0.0018926042783865798, 
    0.0023437973780291634, 0.0029098295008522105, 0.0035620578396203598, 
    0.0042686355265964294, 0.0049965600996826481, 0.0057133554726796817, 
    0.0063884526314001433, 0.0069944240924632237, 0.0075079598854598086, 
    0.0079106665752491367, 0.0081893338606399725, 0.0083359408671133048, 
    0.0083474478844320511, 0.0082258089901898063, 0.0079783909954106724, 
    0.0076183926747135306, 0.0071653096632519923, 0.0066443119343398407, 
    0.0060844665387223438, 0.0055153902428211705, 0.0049627119823551389, 
    0.0044434552915951948, 0.0039622035828985628, 0.0035094231420222922, 
    0.0030627780479657962, 0.002591326858046231, 0.002061653257588573, 
    0.0014444145412322747, 0.00071974658324736301, -0.00011949533074557101, 
    -0.001066215167275884, -0.0020985871536576199, -0.0031799533356076182, 
    -0.0042587460720684908, -0.0052699960951141916, -0.0061391618719429733, 
    -0.0067884280796707917, -0.0071448215803812326, -0.0071481709395002863, 
    -0.0067577213887641029, -0.0059562035545057592, -0.0047507488533307784, 
    -0.0031713355525408381, -0.0012675976537772052, 0.00089551815596785461, 
    0.0032420888023646519, 0.0056894583011454667, 0.0081520246447719606, 
    0.010544193152544734, 0.01278319925455388, 0.01479090395060584, 
    0.016496161071710473, 0.017836939192568471, 0.018763092644475628, 
    0.019239481271210796, 0.019248766110930619, 0.018793215726600983, 
    0.017894682710159822, 0.016591813871196719, 0.014935621983405561, 
    0.012983437314925165, 0.010793486740372352, 0.0084208130237411263, 
    0.005915456835429646, 0.0033235295892588348, 0.00068941417188216102, 
    -0.0019412597617533851, -0.0045190436315584587, -0.0069896477138472572, 
    -0.0092955247982606654, -0.011379074102195784, -0.013187329476841134, 
    -0.014677308434810927, -0.01581960773994566, -0.016600352246677788, 
    -0.017021704282829318, -0.01710230348418057, -0.016878901874609775, 
    -0.016407103866846882, -0.01576098660618537, -0.01502779550323205, 
    -0.014298315189975597, -0.013653565898587457, -0.013152370203458351, 
    -0.012821139395336356, -0.01264856756684229, -0.012587598381242435, 
    -0.012563559752672319, -0.012487170935006436, -0.012267809739140174, 
    -0.011829349794891933, -0.011120845185093847, -0.010126861074637396, 
    -0.0088723122611105917, -0.0074233425587179377, -0.0058815783446477653 ;

 Fqt-total =
  // Fqt-total(0, 0-1999)
    0.99999999999999956, 0.99985957605264542, 0.99943928103314139, 
    0.99874200616144604, 0.99777248846531141, 0.99653721116083827, 
    0.99504427182074517, 0.9933032260871314, 0.99132491292540292, 
    0.98912126874241957, 0.98670513705745955, 0.98409007845849261, 
    0.98129018591304418, 0.97831990917261313, 0.9751938902938021, 
    0.9719268120585286, 0.96853325993705597, 0.9650275994503974, 
    0.9614238656145867, 0.9577356671668652, 0.95397610340565575, 
    0.95015769418833718, 0.94629232390837914, 0.94239119774248103, 
    0.93846481362941137, 0.93452294478916897, 0.93057463268945084, 
    0.92662818935669178, 0.92269120336955712, 0.91877055290170828, 
    0.91487242551694181, 0.9110023404440597, 0.9071651783805178, 
    0.90336521067906905, 0.89960613107349552, 0.89589108800816131, 
    0.89222271745505188, 0.88860317586249704, 0.88503417314521404, 
    0.88151700680001865, 0.87805259404763658, 0.87464150719041889, 
    0.87128400623750224, 0.86798007345880102, 0.86472944633976867, 
    0.86153164984730624, 0.85838602572013478, 0.85529176077959013, 
    0.8522479120938008, 0.84925342946623894, 0.84630717383391518, 
    0.84340793567943761, 0.84055444970617099, 0.8377454085846594, 
    0.83497947288168184, 0.83225528257739267, 0.82957146296850237, 
    0.82692663214536954, 0.82431940704155471, 0.82174840934194637, 
    0.81921226873871844, 0.81670962734222496, 0.81423914341598125, 
    0.81179949198198542, 0.80938937034052072, 0.80700750168999069, 
    0.80465264119261992, 0.80232358288091665, 0.80001916601166689, 
    0.79773828060179153, 0.79547987005411847, 0.79324293231358967, 
    0.791026518346859, 0.78882972744237867, 0.78665170254580796, 
    0.78449162440529718, 0.78234870743418061, 0.78022219450596952, 
    0.77811135278204435, 0.77601547235225921, 0.77393386210947523, 
    0.77186584959999294, 0.76981077870706105, 0.76776800941192125, 
    0.76573691718802683, 0.76371689381351071, 0.76170734667570028, 
    0.75970770140717958, 0.7577174041210365, 0.75573592261306144, 
    0.75376275118038716, 0.75179741392142219, 0.74983946754992425, 
    0.7478885058457212, 0.74594416434882171, 0.74400612435198377, 
    0.74207411704240456, 0.74014792577243094, 0.73822738684275513, 
    0.73631238827765622, 0.73440286607801919, 0.73249880164248593, 
    0.73060021571608491, 0.72870716437885985, 0.72681973433615776, 
    0.72493803890534902, 0.72306221160871031, 0.7211924025893951, 
    0.71932877469513423, 0.71747149749697325, 0.71562074591616343, 
    0.7137766954463215, 0.71193952158403861, 0.71010939655294947, 
    0.70828648869109578, 0.70647095888333855, 0.70466295829043779, 
    0.70286262502739427, 0.70107008326826548, 0.69928544160674078, 
    0.6975087948054276, 0.69574022741127728, 0.69397981687614041, 
    0.69222763674104282, 0.69048375767776982, 0.68874824730544315, 
    0.68702116943208558, 0.68530258246242914, 0.68359253620379667, 
    0.68189106955310974, 0.68019820904611483, 0.67851397044848094, 
    0.67683835743013931, 0.67517136506026898, 0.67351297912622687, 
    0.67186317918933047, 0.67022193973779709, 0.66858922923297037, 
    0.66696501271322217, 0.66534925161766578, 0.66374190552436918, 
    0.66214293192856888, 0.66055228606436522, 0.65896991992782605, 
    0.65739578378464902, 0.65582982288176139, 0.65427197699296147, 
    0.65272217892510265, 0.65118035095632698, 0.64964640160641896, 
    0.64812022305449224, 0.64660168882476676, 0.64509065229045015, 
    0.64358694922221715, 0.64209039669905565, 0.64060080057187951, 
    0.63911795706980612, 0.63764165844452758, 0.63617169631548198, 
    0.63470786683978098, 0.63324997337107669, 0.63179782908409088, 
    0.63035125898996303, 0.6289101008736343, 0.6274742052304132, 
    0.62604343386063621, 0.62461766096706417, 0.62319677054433797, 
    0.62178065794338699, 0.62036923023606738, 0.61896240719032181, 
    0.61756012362539126, 0.61616232916095737, 0.61476898648620226, 
    0.6133800690921738, 0.61199555782044235, 0.61061543823581443, 
    0.60923969558197988, 0.60786831385334117, 0.60650127408568166, 
    0.60513855314751042, 0.60378012612607668, 0.60242596609980104, 
    0.60107604416581273, 0.59973033019036648, 0.59838879180259708, 
    0.5970513904950262, 0.59571808119745728, 0.59438880991353693, 
    0.59306351085775, 0.59174210525088733, 0.59042450149358039, 
    0.58911059521982911, 0.5878002689023234, 0.58649339516070809, 
    0.58518984182378031, 0.58388947420477, 0.58259216280891046, 
    0.58129778507251917, 0.58000623005835439, 0.57871739815126344, 
    0.5774312034115765, 0.57614757508969938, 0.57486646071814163, 
    0.57358782335524194, 0.57231164685064406, 0.57103793298214856, 
    0.56976670152594233, 0.56849799037976079, 0.56723185187095693, 
    0.56596835160726255, 0.56470756559261504, 0.56344957747757451, 
    0.56219447509968656, 0.56094234714387892, 0.55969328285194697, 
    0.55844736715113841, 0.5572046798341711, 0.55596529306170783, 
    0.55472926952115253, 0.55349665937706183, 0.5522674979398644, 
    0.55104180464746921, 0.54981958056178981, 0.54860080620857454, 
    0.54738544176678483, 0.54617342656439738, 0.54496467867644738, 
    0.54375909583956994, 0.54255655601956887, 0.54135691840399691, 
    0.54016002464783652, 0.53896569805731165, 0.53777374590399785, 
    0.53658395981717999, 0.53539611767222406, 0.53420998530439001, 
    0.5330253207363973, 0.53184187723633725, 0.53065940592028638, 
    0.52947766178396471, 0.52829640501226149, 0.52711540446990668, 
    0.52593443957278363, 0.52475330388438146, 0.52357180688028626, 
    0.52238977930706143, 0.52120707305514213, 0.52002356634266766, 
    0.51883916514396256, 0.5176538053494828, 0.51646745279422412, 
    0.51528010128223234, 0.51409177292307584, 0.51290251600537162, 
    0.51171240419958175, 0.51052153705086689, 0.50933003983149039, 
    0.50813806258060268, 0.50694577939992957, 0.50575338675512449, 
    0.50456110167729362, 0.50336915622631573, 0.50217779401587304, 
    0.50098726276308481, 0.49979780986627476, 0.49860967237031939, 
    0.49742307407088354, 0.49623821886006203, 0.49505528678879768, 
    0.49387443221624089, 0.49269578160324518, 0.49151943527252295, 
    0.49034546940247276, 0.4891739365000442, 0.4880048715717859, 
    0.48683829667869216, 0.48567422342158584, 0.48451265762556034, 
    0.48335360299948821, 0.48219706343620905, 0.48104304546377341, 
    0.47989156104284442, 0.47874262819702273, 0.47759627295000767, 
    0.47645253052899095, 0.47531144520256724, 0.47417307159701072, 
    0.47303747291290393, 0.47190472340190748, 0.47077490791678162, 
    0.46964812293470587, 0.46852447511683692, 0.46740408250893606, 
    0.46628707361744826, 0.4651735867071744, 0.4640637686627771, 
    0.46295777412692146, 0.46185576137965467, 0.46075789171856979, 
    0.45966432470118473, 0.45857521418776293, 0.45749070438807438, 
    0.45641092645648518, 0.45533599268342423, 0.45426599530429818, 
    0.45320100153638432, 0.45214105339749716, 0.4510861688270541, 
    0.45003634605359022, 0.4489915670698516, 0.44795180350071928, 
    0.44691702075069278, 0.4458871833925061, 0.44486225831584936, 
    0.44384222082986335, 0.44282705805650352, 0.44181676969509504, 
    0.44081137283131894, 0.43981090105611004, 0.43881540753844334, 
    0.43782496009018984, 0.43683964387950081, 0.43585955798972381, 
    0.43488481311996985, 0.43391553041080361, 0.4329518395930787, 
    0.43199387700375103, 0.43104178411412203, 0.43009570572451511, 
    0.42915578592296205, 0.42822216494999099, 0.42729497459011911, 
    0.42637433311870948, 0.42546034033998481, 0.42455307450095164, 
    0.42365258973766901, 0.42275891457767772, 0.42187205255802795, 
    0.42099198418656231, 0.4201186697737897, 0.41925205160658047, 
    0.41839205634033033, 0.41753859789788139, 0.41669157589926797, 
    0.41585087715888508, 0.41501637382133977, 0.41418792507321234, 
    0.41336537589308281, 0.41254855740500773, 0.4117372861739112, 
    0.41093136694828059, 0.41013058717853229, 0.40933471692215595, 
    0.40854350690905145, 0.40775668465198261, 0.40697395434679429, 
    0.40619499958868738, 0.40541948442085429, 0.40464705859723887, 
    0.40387736085786652, 0.4031100239231552, 0.40234467807338348, 
    0.40158095651541104, 0.40081850192929647, 0.40005697269741536, 
    0.39929605003953272, 0.39853544342078195, 0.39777489483820472, 
    0.39701418028607782, 0.39625310907900785, 0.39549152155119682, 
    0.39472928559688392, 0.39396629354615958, 0.39320245922870423, 
    0.39243771745547246, 0.39167202175100896, 0.39090534389613313, 
    0.39013767526022092, 0.38936902237031218, 0.38859940677070937, 
    0.38782886182592319, 0.38705743029166628, 0.38628515961471671, 
    0.38551210090262994, 0.3847383072734471, 0.38396383007475743, 
    0.38318871546960465, 0.38241300605500539, 0.38163673766052147, 
    0.38085994277762547, 0.38008265305866806, 0.37930490421286944, 
    0.37852673612941168, 0.3777481944263692, 0.37696932519028625, 
    0.37619017697849921, 0.37541079664209254, 0.37463123040679575, 
    0.37385152595541227, 0.37307173246471781, 0.37229190405108936, 
    0.37151210129212886, 0.37073239124277502, 0.36995284545219431, 
    0.36917353961213856, 0.36839454689495554, 0.36761593630592265, 
    0.3668377669355633, 0.36606008585957311, 0.36528292348357677, 
    0.36450629436926318, 0.3637301959027141, 0.36295461104835636, 
    0.36217951175926005, 0.36140486610788652, 0.36063064481531526, 
    0.35985682814858577, 0.35908341218018919, 0.35831041304677891, 
    0.35753786802538762, 0.35676583578123416, 0.35599439173017972, 
    0.35522362358229881, 0.35445362787321777, 0.35368450320211031, 
    0.35291634610808581, 0.35214924797627689, 0.35138329314245881, 
    0.35061856126515067, 0.34985512848470185, 0.34909307346393809, 
    0.34833247652159288, 0.34757342291868942, 0.34681599998051427, 
    0.34606029659828619, 0.34530639913853145, 0.34455439093974333, 
    0.34380434952064776, 0.34305634579667077, 0.34231044211218487, 
    0.34156669075513529, 0.34082513170374956, 0.34008579195169769, 
    0.33934868021743531, 0.3386137865765097, 0.33788107878069712, 
    0.33715050032274319, 0.33642197032380183, 0.33569538580101793, 
    0.3349706272693917, 0.3342475675853504, 0.33352608127616756, 
    0.33280605642929723, 0.33208739822440059, 0.33137003380389723, 
    0.33065391120195847, 0.3299389959459294, 0.32922526782393419, 
    0.32851271601712512, 0.32780133503003317, 0.32709112043503213, 
    0.32638206621431626, 0.32567416364614366, 0.32496740310114419, 
    0.32426177603764006, 0.32355728035820497, 0.32285392457597317, 
    0.32215173312474193, 0.32145074968352211, 0.32075104020096096, 
    0.32005269387740476, 0.3193558232073555, 0.31866056154415379, 
    0.31796706349741743, 0.31727550069871724, 0.31658605926057004, 
    0.31589893712587896, 0.31521434216215349, 0.31453248478424084, 
    0.31385357774996991, 0.31317782977953823, 0.3125054429937888, 
    0.31183661049182859, 0.31117151469404752, 0.31051032645337967, 
    0.30985320337006422, 0.30920029110981628, 0.30855172115713891, 
    0.30790761209042911, 0.30726806580741961, 0.30663316905922722, 
    0.3060029901738614, 0.30537757631647761, 0.30475695457805413, 
    0.30414113104717, 0.30353009069742348, 0.30292380009661762, 
    0.30232220541384913, 0.30172523482009, 0.30113279520407388, 
    0.30054477506767119, 0.29996104154214742, 0.29938143971425163, 
    0.2988057931757816, 0.29823390159266272, 0.29766554438751197, 
    0.29710048504409886, 0.2965384745281735, 0.29597925949526344, 
    0.29542258754189815, 0.29486821310175831, 0.29431590115712702, 
    0.29376543031729863, 0.29321659571082187, 0.29266921211288355, 
    0.2921231127300144, 0.29157815174407298, 0.29103420448731787, 
    0.29049116607005543, 0.28994895205542043, 0.2894074948026969, 
    0.2888667438124724, 0.28832666489133546, 0.28778723942376194, 
    0.2872484655611825, 0.28671035718917404, 0.28617294342819566, 
    0.28563626432329425, 0.28510037048082726, 0.28456531755073111, 
    0.28403116551216273, 0.28349797701216489, 0.28296581706305668, 
    0.28243475264783391, 0.28190485282023603, 0.28137618671642084, 
    0.28084882450919718, 0.28032283517052181, 0.2797982839721157, 
    0.27927523168317891, 0.27875373415063759, 0.27823384034220344, 
    0.27771559714729865, 0.27719904982445304, 0.27668424465391334, 
    0.27617123268060573, 0.27566007079355637, 0.27515082268455809, 
    0.27464355807915963, 0.2741383520822509, 0.27363528147902799, 
    0.27313442006921013, 0.27263583751367743, 0.27213959279337796, 
    0.27164573100191874, 0.27115428061548785, 0.27066525170237887, 
    0.27017863584840723, 0.26969440666334482, 0.26921252294487935, 
    0.26873292964191797, 0.26825556192860367, 0.26778034448996546, 
    0.26730719659692403, 0.26683603059593963, 0.26636675613360666, 
    0.26589928095678983, 0.26543351316804525, 0.26496936223540335, 
    0.2645067426749364, 0.2640455725577161, 0.26358577694097257, 
    0.26312728744212988, 0.26267004277105466, 0.26221398890727438, 
    0.26175907553905614, 0.2613052570501051, 0.26085248696773272, 
    0.26040071814598392, 0.25994989849341604, 0.25949997054661389, 
    0.25905087348597922, 0.25860254376694503, 0.25815491917917632, 
    0.25770794219337462, 0.25726156514092313, 0.2568157510432707, 
    0.2563704756067316, 0.25592572584983597, 0.2554814985000663, 
    0.25503779772843438, 0.25459463301450358, 0.25415201655826475, 
    0.25370996221535302, 0.25326848251774003, 0.25282758744557315, 
    0.25238728146294442, 0.25194756073200814, 0.25150841102805849, 
    0.25106980357441483, 0.25063169623390757, 0.25019403173412003, 
    0.24975673850612387, 0.24931973294131546, 0.24888292393192285, 
    0.24844621827134172, 0.24800952816064839, 0.24757277646077278, 
    0.24713590618470355, 0.2466988833295273, 0.24626170020858262, 
    0.24582437829921108, 0.24538696330046986, 0.24494952410019175, 
    0.24451215052722211, 0.24407494769807331, 0.24363803252011063, 
    0.24320152985057564, 0.24276556852903555, 0.24233027704098822, 
    0.24189578183625662, 0.24146220300560634, 0.24102965267791132, 
    0.24059823487059442, 0.24016804227950822, 0.2397391579004135, 
    0.23931165446421068, 0.23888559099240683, 0.23846101401284314, 
    0.23803795540863926, 0.23761643059145193, 0.23719643929844941, 
    0.23677796688592931, 0.23636098424496274, 0.23594545231717309, 
    0.23553132303507704, 0.23511854482771466, 0.23470706250005682, 
    0.2342968207315245, 0.23388776721365442, 0.23347984991657461, 
    0.23307302204102337, 0.23266723828899982, 0.23226245810416532, 
    0.23185864269313622, 0.23145575599641849, 0.23105376486323403, 
    0.23065263744780856, 0.2302523432581656, 0.22985285262988839, 
    0.22945413573664039, 0.22905616231172291, 0.22865890068254696, 
    0.22826231574727032, 0.22786636994108356, 0.22747102085903387, 
    0.22707621971376113, 0.22668191060419579, 0.22628802843353826, 
    0.22589449820467775, 0.22550123426059016, 0.2251081415011317, 
    0.22471511784100157, 0.22432205887619483, 0.22392886047734745, 
    0.22353542386607383, 0.22314165704964817, 0.22274747834495459, 
    0.22235281789721484, 0.22195761806148187, 0.2215618358642, 
    0.22116544333928342, 0.22076842462444016, 0.22037077665413679, 
    0.21997250576762342, 0.21957362447879353, 0.21917414742922192, 
    0.21877408978596888, 0.21837346363688245, 0.21797227391176602, 
    0.21757051905254404, 0.2171681899479829, 0.21676527170725948, 
    0.21636174468836705, 0.21595759107091553, 0.21555279944462269, 
    0.21514737114497212, 0.21474132480043878, 0.21433470130281559, 
    0.21392756717630432, 0.21352001936757711, 0.21311218666408444, 
    0.21270422757883783, 0.21229632634375206, 0.2118886838427782, 
    0.21148150852352213, 0.21107500901527679, 0.21066938852742773, 
    0.21026484524076086, 0.20986157436497521, 0.2094597686247317, 
    0.20905961957544111, 0.20866131797396362, 0.20826505127559491, 
    0.20787100189195254, 0.20747934620497002, 0.20709024870720869, 
    0.20670386215023584, 0.20632032517207347, 0.20593975978508378, 
    0.20556227043818956, 0.20518794271775412, 0.2048168430544598, 
    0.20444901622270911, 0.20408448627149992, 0.20372325587498658, 
    0.20336530647930121, 0.20301059831894616, 0.20265907248583098, 
    0.20231065156883404, 0.20196524036826641, 0.20162272708661994, 
    0.20128298392157201, 0.20094586555987609, 0.20061120917568748, 
    0.2002788323249636, 0.19994853050055514, 0.19962007938430251, 
    0.19929323345897154, 0.19896773155398798, 0.19864329857762877, 
    0.19831964942939939, 0.19799649444403358, 0.19767354062624493, 
    0.19735049503365482, 0.1970270700717944, 0.19670298768026512, 
    0.1963779847747521, 0.19605181727154034, 0.19572426772565593, 
    0.19539514755871845, 0.19506430016051013, 0.19473160201067433, 
    0.19439696089395067, 0.19406031558783657, 0.19372163130738365, 
    0.19338089757128424, 0.19303812424629035, 0.19269333825794938, 
    0.19234657582461465, 0.19199787747810843, 0.19164728341871778, 
    0.19129482526463032, 0.19094052578600115, 0.19058439522991691, 
    0.19022643361333885, 0.18986663145697943, 0.18950497311345435, 
    0.1891414399080982, 0.18877601280586795, 0.18840867593309682, 
    0.18803941964503137, 0.18766824331296758, 0.18729515760823412, 
    0.18692018784314532, 0.18654337540497987, 0.18616477755132435, 
    0.18578446793278924, 0.1854025331329297, 0.18501907073375048, 
    0.18463418491328654, 0.18424798220771466, 0.18386056875003001, 
    0.18347204684079099, 0.18308251344738674, 0.18269205990844545, 
    0.18230077545656864, 0.18190874728521739, 0.18151606444101945, 
    0.18112282095511817, 0.18072911858117902, 0.18033506808600774, 
    0.17994079223843687, 0.17954642492560172, 0.17915211272678983, 
    0.17875801419283324, 0.17836429921069186, 0.17797114886256829, 
    0.17757875325109845, 0.17718731091795512, 0.17679702460436569, 
    0.1764081009485903, 0.17602074598663606, 0.17563516580671862, 
    0.17525156200004369, 0.17487013204052754, 0.17449106610166867, 
    0.17411454744939284, 0.1737407482428685, 0.17336983107444906, 
    0.17300194335070584, 0.17263721814697877, 0.17227576981643847, 
    0.17191769317304972, 0.17156305882997622, 0.1712119103636521, 
    0.1708642629972259, 0.17052010102846679, 0.17017937398213356, 
    0.16984199496390703, 0.16950784004963415, 0.16917674845003225, 
    0.16884852568871106, 0.16852294464627335, 0.16819975101376608, 
    0.16787866739539076, 0.16755939692861224, 0.16724162659334274, 
    0.1669250355222221, 0.16660929716885897, 0.16629408417385588, 
    0.16597907610903448, 0.16566396445918538, 0.16534845595657435, 
    0.16503227711716406, 0.16471517531125299, 0.16439691813638413, 
    0.16407729734901433, 0.16375612742780993, 0.16343324927982958, 
    0.16310852950296448, 0.16278186208204154, 0.1624531655443644, 
    0.16212238247344682, 0.16178947587134199, 0.16145442829041898, 
    0.16111723974421185, 0.16077792425826357, 0.16043650768548204, 
    0.16009302928863078, 0.15974753496905539, 0.15940007911101051, 
    0.15905071985368038, 0.15869951962255807, 0.15834653877723132, 
    0.1579918373096271, 0.15763547144471607, 0.1572774931416028, 
    0.15691794907531734, 0.15655688362686093, 0.15619433987321973, 
    0.15583036418501153, 0.15546500813618203, 0.1550983316934087, 
    0.15473040527393128, 0.1543613125468071, 0.15399114747788553, 
    0.15362001680728038, 0.15324804075587387, 0.15287535303386049, 
    0.15250210627303964, 0.15212847114673103, 0.1517546400599617, 
    0.15138082399035482, 0.15100725060477002, 0.15063416164671764, 
    0.15026180647744558, 0.14989043646381486, 0.1495203010731527, 
    0.1491516442919763, 0.1487847000275723, 0.14841968883118739, 
    0.1480568127171222, 0.14769625479680148, 0.14733817734687199, 
    0.14698271884712963, 0.14662999638732221, 0.14628010570531588, 
    0.14593312083208299, 0.14558909590703806, 0.14524806477297664, 
    0.14491004159503565, 0.14457502297750718, 0.14424298357256499, 
    0.14391388261186511, 0.14358766504408929, 0.14326426316483609, 
    0.14294360056696856, 0.14262559533100844, 0.14231016239014807, 
    0.14199721473389909, 0.14168666457033521, 0.14137842533126946, 
    0.14107240958434195, 0.14076852976401011, 0.14046669951904814, 
    0.1401668327649111, 0.13986884844741437, 0.13957267025438125, 
    0.13927823100836315, 0.13898547623568197, 0.13869436762895587, 
    0.13840488701509382, 0.13811704230777988, 0.13783087215469123, 
    0.13754644948839992, 0.13726388713396484, 0.13698333570228172, 
    0.13670498356987029, 0.13642905228819394, 0.13615579023776736, 
    0.13588546832617809, 0.13561837092237738, 0.13535479378625018, 
    0.13509503765905728, 0.13483940340177539, 0.13458818955211044, 
    0.13434168743089717, 0.13410017841717517, 0.13386392935990582, 
    0.13363318925724957, 0.13340818467890644, 0.13318911546769527, 
    0.1329761511492297, 0.132769426355584, 0.13256903873685527, 
    0.13237504639937439, 0.13218746595876593, 0.13200627393340081, 
    0.13183140551054873, 0.13166275778000783, 0.13150018996310964, 
    0.13134352698374735, 0.13119256293771403, 0.1310470640208119, 
    0.1309067710047811, 0.13077140327888997, 0.13064066193444171, 
    0.13051423349661193, 0.13039179610720397, 0.13027302139123051, 
    0.13015757998709435, 0.1300451460771119, 0.12993540062024639, 
    0.12982803098549497, 0.12972273547929472, 0.12961922221033165, 
    0.12951721089197971, 0.1294164321538718, 0.12931662886419096, 
    0.1292175558781927, 0.12911897937282776, 0.12902067796857694, 
    0.12892244022076454, 0.12882406491577503, 0.12872535847441743, 
    0.12862613429698877, 0.12852621238952974, 0.12842541922603123, 
    0.12832359022399945, 0.12822057022039851, 0.12811621717371885, 
    0.12801040677945996, 0.1279030311411152, 0.12779400259406071, 
    0.12768325485575732, 0.1275707433044698, 0.12745644547013024, 
    0.12734035850553863, 0.12722250100693344, 0.12710290713922848, 
    0.12698162619360659, 0.1268587185885984, 0.12673425200062824, 
    0.12660829882112939, 0.1264809306598523, 0.12635221723252082, 
    0.12622222406354247, 0.12609101337087789, 0.12595864602280768, 
    0.12582518178156721, 0.12569068660636293, 0.12555523249218442, 
    0.12541889976836795, 0.12528177906149252, 0.12514396627533045, 
    0.12500556114724798, 0.12486666147792794, 0.12472735842472214, 
    0.12458772955674723, 0.12444783526774887, 0.12430771730967428, 
    0.12416739480708196, 0.12402686403444987, 0.12388609848123461, 
    0.12374504718463289, 0.1236036354823622, 0.12346176560428865, 
    0.12331931816540213, 0.12317615300907944, 0.12303211428639696, 
    0.1228870311891396, 0.12274072795443412, 0.12259302623956461, 
    0.12244375479819222, 0.12229275691826737, 0.12213989704770127, 
    0.12198506856766066, 0.12182819883417338, 0.12166925575460025, 
    0.12150824982020761, 0.12134523220989314, 0.12118029442695495, 
    0.12101355945507014, 0.12084517519896296, 0.12067530267978378, 
    0.12050410965600065, 0.12033175986759928, 0.12015840602512205, 
    0.11998418454137999, 0.11980921304195596, 0.11963358662144721, 
    0.119457379350155, 0.11928064525126511, 0.11910341839870563, 
    0.11892571733123902, 0.11874754927889852, 0.11856891023180335, 
    0.11838979156803479, 0.11821018223192087, 0.11803007335643641, 
    0.11784946048979582, 0.11766834779341001, 0.11748675195688632, 
    0.11730470435548232, 0.11712225223902821, 0.11693946284189349, 
    0.11675642049288147, 0.11657322658721006, 0.11638999678050069, 
    0.11620685693651167, 0.11602393873158789, 0.1158413739455313, 
    0.11565929283741826, 0.1154778194673324, 0.11529706680555894, 
    0.11511713930560398, 0.1149381285981553, 0.11476011476788704, 
    0.11458316543647673, 0.1144073391002989, 0.11423268223284949, 
    0.11405923284911394, 0.11388702274009917, 0.11371607860650862, 
    0.11354642457816864, 0.11337808147442106, 0.11321106656616342, 
    0.1130453941424505, 0.11288107113330506, 0.11271809812381357, 
    0.11255646497458831, 0.11239614670323411, 0.11223709927508173, 
    0.11207925463159438, 0.11192251506797984, 0.11176675443378054, 
    0.11161181975615003, 0.11145753247959912, 0.11130369489630559, 
    0.1111500970802814, 0.11099652038342284, 0.1108427442710916, 
    0.11068855169068256, 0.11053373232866832, 0.11037808571261819, 
    0.11022142364973833, 0.11006356982994168, 0.10990435788486358, 
    0.10974362993719795, 0.10958123434486448, 0.10941702169346001, 
    0.10925084291876655, 0.10908255059946133, 0.10891200025947194, 
    0.10873905282395835, 0.1085635801903566, 0.10838546776106812, 
    0.10820461755231148, 0.10802094675110936, 0.1078343900274891, 
    0.10764489459159449, 0.10745241930677946, 0.10725693230106294, 
    0.10705840677251452, 0.10685681954801025, 0.10665214887693471, 
    0.10644437224317928, 0.10623346567098317, 0.10601940368469284, 
    0.1058021596635301, 0.10558170717957231, 0.10535802129662308, 
    0.10513107951885363, 0.10490086574741034, 0.10466736981031245, 
    0.10443058851928511, 0.10419052835900326, 0.10394720743887072, 
    0.10370065555624304, 0.1034509195851218, 0.10319806312872025, 
    0.10294217242765336, 0.10268335882449353, 0.10242176217948745, 
    0.10215755301656201, 0.10189093222307154, 0.10162213195280642, 
    0.10135141159316112, 0.10107905517934813, 0.10080536554300321, 
    0.10053065921345855, 0.10025525936369531, 0.099979490537901533, 
    0.099703673212572716, 0.099428118062468984, 0.099153122937793617, 
    0.098878969812096235, 0.098605921604163052, 0.098334221002900929, 
    0.098064090228060258, 0.097795729976029269, 0.097529322991743064, 
    0.09726503102864735, 0.097003000310355122, 0.096743359109594487, 
    0.096486218620771197, 0.096231673951494845, 0.095979804103045491, 
    0.095730670966442666, 0.095484324517305097, 0.095240800946891302, 
    0.095000129112835494, 0.094762331073212941, 0.094527424566214754, 
    0.094295423623669716, 0.094066339848883893, 0.093840181702047359, 
    0.093616954705019947, 0.093396661900424116, 0.093179304444284475, 
    0.092964880088170082, 0.092753383027644937, 0.092544802752014918, 
    0.092339122212065611, 0.092136316057104914, 0.09193635067777868, 
    0.09173918322694137, 0.091544760995391439, 0.091353021267418108, 
    0.091163893710815722, 0.090977300486605364, 0.090793159933773293, 
    0.090611389368382977, 0.090431905314969432, 0.090254625443642642, 
    0.090079468916731326, 0.089906354321680898, 0.08973519591426804, 
    0.089565902036266229, 0.08939837503668778, 0.089232509630699397, 
    0.089068195486977336, 0.088905317565003306, 0.088743761359485085, 
    0.088583411719049779, 0.088424155779885993, 0.08826588366517267, 
    0.088108490222902208, 0.087951875402034571, 0.087795946395272342, 
    0.087640620392077664, 0.087485828728712481, 0.087331517893530108, 
    0.087177655905409046, 0.087024231351072831, 0.086871258429345288, 
    0.086718775387602462, 0.086566844289013206, 0.08641555160667673, 
    0.086265005571177888, 0.086115332985424078, 0.085966678577425265, 
    0.08581920001787309, 0.085673065053591763, 0.085528448077898722, 
    0.085385527544288575, 0.085244480421902996, 0.085105483285960487, 
    0.084968709176766258, 0.084834328436686021, 0.084702510320035701, 
    0.084573423120922558, 0.084447232676993306, 0.084324098565207617, 
    0.084204170756093655, 0.084087583973588564, 0.083974452857506349, 
    0.083864872329969711, 0.083758912046706976, 0.083656617601426814, 
    0.083558008573446571, 0.083463077734400676, 0.083371787537185563, 
    0.083284070152041978, 0.083199824347640408, 0.083118913573975842, 
    0.083041170915389706, 0.082966397175527548, 0.082894365795197392, 
    0.082824825381085904, 0.08275750694292755, 0.082692121303805433, 
    0.082628366344569146, 0.082565926996115022, 0.082504475352717446, 
    0.082443673542572773, 0.082383170359685023, 0.082322606367566331, 
    0.08226161504057318, 0.082199824069957086, 0.08213686227815889, 
    0.082072363625814507, 0.082005971890703508, 0.081937345268988632, 
    0.081866159152256326, 0.081792108744021375, 0.0817149107574726, 
    0.081634305501944102, 0.081550060322147566, 0.081461969558069877, 
    0.081369860046731607, 0.081273589190227022, 0.081173050714751685, 
    0.081068170588526986, 0.080958908685828265, 0.080845255110124345, 
    0.080727227322997808, 0.080604865910020335, 0.080478229835703866, 
    0.080347395009836522, 0.080212445788531914, 0.080073472712575755, 
    0.079930565888971017, 0.079783811266168528, 0.079633284251899264, 
    0.079479052341548159, 0.079321171432476134, 0.079159692112271057, 
    0.078994663143234584, 0.078826134113105489, 0.07865416044961393, 
    0.078478806089279568, 0.07830014461386535, 0.078118265216745128, 
    0.077933271597634107, 0.077745288430897327, 0.077554459214427135, 
    0.077360945959423499, 0.077164924564731119, 0.076966580550968, 
    0.076766106675750206, 0.076563694380417033, 0.076359529471575455, 
    0.076153784428561258, 0.075946617021066615, 0.075738161259800152, 
    0.075528523430515915, 0.075317776933881711, 0.075105959733826513, 
    0.074893073842033864, 0.074679088425265522, 0.074463945923289407, 
    0.074247568986446993, 0.074029873602274435, 0.07381077644925349, 
    0.073590209111795035, 0.07336812027306075, 0.073144484889045389, 
    0.072919299516749858, 0.072692585624058795, 0.072464383574861721, 
    0.07223474902660304, 0.072003747646513669, 0.071771447395627269, 
    0.071537916119463751, 0.071303213227389847, 0.071067389414263341, 
    0.070830480304410207, 0.070592510526302041, 0.070353493525310645, 
    0.070113436506490046, 0.069872345657628732, 0.069630231190349154, 
    0.069387113029395556, 0.069143027691487266, 0.068898034222046281, 
    0.068652224800998293, 0.068405728736277954, 0.068158718542343524, 
    0.067911409713483098, 0.067664057956679985, 0.06741695221454154, 
    0.067170411932323579, 0.066924779893044281, 0.066680416559170272, 
    0.066437697738308543, 0.066197007798156224, 0.065958730279748426, 
    0.065723245471307049, 0.065490919948403739, 0.065262095459592287, 
    0.06503708449235325, 0.064816160331306438, 0.064599549977425466, 
    0.064387428333768634, 0.064179918473538086, 0.063977089841853629, 
    0.063778963966118291, 0.063585519307485655, 0.063396704422894648, 
    0.063212446855745424, 0.063032666241690169, 0.062857281669532528, 
    0.062686220360665637, 0.062519418178537414, 0.062356818833868961, 
    0.062198373097719861, 0.062044034315717117, 0.061893756218079833, 
    0.061747497877876451, 0.061605220197955231, 0.061466890749502991, 
    0.061332481827336201, 0.061201966912634506, 0.061075311663040886, 
    0.060952465097087204, 0.060833350648691789, 0.060717860342323814, 
    0.060605849976995203, 0.060497142736737619, 0.060391530210846811, 
    0.060288774888914369, 0.060188622512907408, 0.060090808601989593, 
    0.059995069248066246, 0.059901149952257239, 0.059808817532942496, 
    0.059717860472288622, 0.05962809019984721, 0.059539340644647061, 
    0.059451462248150032, 0.059364318363748385, 0.059277781912407894, 
    0.05919173151036921, 0.059106052777539324, 0.059020643073244568, 
    0.058935409979159657, 0.058850278672871792, 0.058765194621510003, 
    0.058680125082618162, 0.058595060059543652, 0.058510010299258682, 
    0.058425002635217688, 0.058340074106046531, 0.058255270885610937, 
    0.058170643348931815, 0.058086243077490898, 0.058002126181927481, 
    0.057918355290892565, 0.057835001469514896, 0.057752146934776961, 
    0.05766988362597858, 0.057588310204896589, 0.057507537144981517, 
    0.057427680073283242, 0.057348862256005564, 0.057271215349224053, 
    0.057194877921346372, 0.057119996753895945, 0.057046723496659221, 
    0.056975216847618991, 0.056905632892740365, 0.056838127390158324, 
    0.056772847207002042, 0.05670992787921534, 0.056649487997843417, 
    0.056591623266081643, 0.056536406585845897, 0.056483883481158258, 
    0.056434072215771666, 0.056386960806617745, 0.05634250948304334, 
    0.056300651981911372, 0.056261294869594788, 0.056224322534959993, 
    0.056189600006822743, 0.056156985167397561, 0.056126332010354524, 
    0.056097502887704737, 0.056070375693402667, 0.056044845650993561, 
    0.056020831017983545, 0.055998271048883295, 0.055977124280816845, 
    0.055957368430931805, 0.055938995502869841, 0.055922012528332614, 
    0.055906440730495305, 0.055892310819372522, 0.055879667341087742, 
    0.055868564838764408, 0.055859072261820499, 0.055851270055248259, 
    0.055845250382027874, 0.055841119551830971, 0.055838995237524482, 
    0.055839009244761019, 0.055841304438001733, 0.055846031223060422, 
    0.055853348250786153, 0.055863412720028496, 0.055876383490445589, 
    0.055892411136055663, 0.055911638959136103, 0.055934196990512858, 
    0.055960201961050948, 0.055989757450764212, 0.05602295237487518, 
    0.056059860129138384, 0.05610053643308343, 0.056145021304686828, 
    0.05619333310595552, 0.056245467671326134, 0.056301395074395556, 
    0.056361058917008086, 0.05642437757281666, 0.056491242457162583, 
    0.05656152559938827, 0.056635077030284614, 0.056711729602275787, 
    0.056791302761532859, 0.056873604498755885, 0.05695843128035586, 
    0.057045571317392747, 0.057134802065085671, 0.057225888941455146, 
    0.057318588352295079, 0.057412641725383358, 0.057507782346609776, 
    0.057603739370998365, 0.057700241681791338, 0.057797026363116143, 
    0.057893845206282248, 0.057990468685042922, 0.058086692459033577, 
    0.0581823367313433, 0.058277252729760712, 0.058371322135816507, 
    0.058464455783542431, 0.058556592474412361, 0.05864769247044941, 
    0.058737729251474698, 0.05882668389626923, 0.058914534734470003, 
    0.059001251252465484, 0.059086791508413734, 0.059171104063826065, 
    0.059254134699090737, 0.059335830691801698, 0.059416148796444065, 
    0.059495058951414263, 0.059572547768492398, 0.059648622919445164, 
    0.059723317777861502, 0.059796696874219832, 0.059868856243486625, 
    0.059939928199981042, 0.06001007584718971, 0.060079488041012354, 
    0.060148371643745674, 0.06021693777462335, 0.06028539287955835, 
    0.060353931763786554, 0.060422736728161654, 0.060491978113613495, 
    0.060561817596294344, 0.06063241534497435, 0.06070392770278691, 
    0.060776503244517603, 0.060850277463442182, 0.060925364569052155, 
    0.06100185382253407, 0.061079805635329242, 0.061159253183892585, 
    0.061240204096384074, 0.061322640628595104, 0.061406524366041736, 
    0.061491798525278266, 0.061578388771157198, 0.061666211659224132, 
    0.061755163712287113, 0.061845128747929669, 0.061935972252419362, 
    0.062027538753186715, 0.062119651951045803, 0.062212110926505734, 
    0.062304693102256128, 0.062397157579536532, 0.062489247741227341, 
    0.062580699896557429, 0.062671247026483565, 0.06276062777612168, 
    0.062848586904896198, 0.062934881322094821, 0.063019281156798251, 
    0.063101571609114449, 0.063181553952923963, 0.063259037875011456, 
    0.063333840972002439, 0.063405779410966145, 0.063474661861524603, 
    0.063540283091373231, 0.063602417503619821, 0.063660812978106357, 
    0.063715192349820676, 0.06376525609894905, 0.063810684622848113, 
    0.063851143787352044, 0.063886301342041305, 0.063915827351183674, 
    0.063939408333136938, 0.063956749328922272, 0.063967577209526769, 
    0.063971644721728602, 0.063968729530042651, 0.063958636887081269, 
    0.063941196865357514, 0.063916270303963366, 0.063883753779752792, 
    0.063843582593968357, 0.063795744075577782, 0.063740280255398366, 
    0.063677297949156594, 0.063606965489793832, 0.063529509440888199, 
    0.063445216154959461, 0.063354422389474793, 0.06325751008398664, 
    0.063154907250242628, 0.063047076443205827, 0.062934512982873461, 
    0.062817738306443688, 0.06269730030277014, 0.062573764969824433, 
    0.062447711803485476, 0.062319728875077071, 0.062190401375879792, 
    0.062060299199400926, 0.061929965263731131, 0.061799899514609541, 
    0.061670551679829926, 0.061542308526585508, 0.061415492929052504, 
    0.061290360409199149, 0.061167101670297312, 0.061045841974521731, 
    0.060926647650065197, 0.060809531891061287, 0.060694457049236185, 
    0.060581339753848149, 0.060470058397401577, 0.060360461739308514, 
    0.060252375727543869, 0.060145615643589799, 0.060039996268038222, 
    0.059935337733896775, 0.059831473059995102, 0.059728253683020816, 
    0.059625551488957804, 0.059523258387166246, 0.059421287589445176, 
    0.059319575855306367, 0.059218083153067057, 0.059116790511370684, 
    0.05901570404333837, 0.058914848234940795, 0.058814268401627262, 
    0.058714028413966141, 0.058614204397158462, 0.058514882530765082, 
    0.05841615724154537, 0.058318125052904568, 0.058220881753228551, 
    0.058124518206812012, 0.058029118007406393, 0.05793475263678622, 
    0.057841477773198723, 0.057749331115117999, 0.057658323718167238, 
    0.057568440870495972, 0.057479642938410347, 0.057391875273631994, 
    0.057305075419182526, 0.057219178678203288, 0.057134122341990404, 
    0.057049844208801853, 0.056966277802195008, 0.056883353251706764, 
    0.056800989956285144, 0.056719100497303859, 0.056637585951410926, 
    0.05655633467718222, 0.056475228895514651, 0.056394146192179584, 
    0.056312964870788532, 0.056231573143079271, 0.056149879665383103, 
    0.056067824097321646, 0.055985387405521503, 0.055902604491245039, 
    0.055819568320945215, 0.055736435891929045, 0.055653425985465618, 
    0.055570810169321493, 0.055488901661184468, 0.055408040780398064, 
    0.055328572055444857, 0.055250831631125132, 0.055175129054462077, 
    0.05510174035356713, 0.055030891646924728, 0.054962758289033325, 
    0.05489746093523281, 0.05483506339027943, 0.054775576431680052, 
    0.054718967894631973, 0.05466517328246568, 0.054614112840114526, 
    0.054565706696885506, 0.054519884981077515, 0.054476588606378287, 
    0.05443577000144692, 0.054397384696621205, 0.054361384654733912, 
    0.054327712220901644, 0.054296289994287074, 0.054267023059567383, 
    0.054239794910717266, 0.054214474037300571, 0.054190913608310992, 
    0.054168959384599764, 0.0541484525751256, 0.054129236685729762, 
    0.05411116069870648, 0.05409408714905499, 0.05407789033912426, 
    0.054062461516902971, 0.05404770836604731, 0.054033558812446002, 
    0.054019954885277936, 0.05400685313015121, 0.053994216737113368, 
    0.053982017427301049, 0.053970235634989157, 0.053958857547896838, 
    0.053947889066687404, 0.053937357313358053, 0.053927308778984058, 
    0.053917817669055595, 0.05390897801691235, 0.05390090386892054, 
    0.053893717240641764, 0.053887551722460049, 0.053882542693964398, 
    0.053878822638800387, 0.0538765250504466, 0.053875769396765652, 
    0.053876671271345683, 0.053879334344033927, 0.053883846463394357, 
    0.053890284127435656, 0.053898709220605884, 0.053909177481872919, 
    0.05392173710081264, 0.053936445001569418, 0.053953363343404941, 
    0.053972565774765287, 0.053994138779161455, 0.054018177780425676, 
    0.054044796098833274, 0.054074118256158897, 0.054106281409624299, 
    0.054141438547003429, 0.054179745210760633, 0.054221355554549204, 
    0.054266418487185636, 0.05431507461783662, 0.054367444791845188, 
    0.054423626592443444, 0.05448369795261844, 0.05454771609413802, 
    0.054615713671657302, 0.054687710032231829, 0.054763703587870645, 
    0.054843679460823469, 0.054927601233782104, 0.055015416414478158, 
    0.055107047564308155, 0.055202394431073859, 0.055301327173773118, 
    0.055403689435646858, 0.05550928889043133, 0.055617907142930072, 
    0.055729292730665195, 0.055843175142103955, 0.05595927203665349, 
    0.056077301720588342, 0.056196994617504735, 0.056318104176982409, 
    0.05644041110375269, 0.056563723068823867, 0.056687871688634983, 
    0.056812701055184621, 0.056938051299469286, 0.057063756574255865, 
    0.057189632500518728, 0.05731546450390336, 0.057441015021973303, 
    0.057566017642719236, 0.057690193125115682, 0.057813248156647234, 
    0.057934882718635457, 0.058054799242456746, 0.058172705261138123, 
    0.058288322611869836, 0.058401397099767133, 0.058511704400872853, 
    0.058619070031428487, 0.058723374117638137, 0.058824554222463542, 
    0.058922603610376517, 0.059017561563666464, 0.059109498150540639, 
    0.059198494833273892, 0.05928462078464531, 0.059367922295530576, 
    0.059448413668959268, 0.059526077804048991, 0.059600874129094886, 
    0.05967274603498695, 0.059741628637616367, 0.059807453252905027, 
    0.059870154436180628, 0.059929657332988252, 0.059985878843386478, 
    0.0600387328811103, 0.060088120462877211, 0.060133937916612583, 
    0.060176082921126701, 0.060214460140930251, 0.06024898880609781, 
    0.060279612929996153, 0.060306294251246596, 0.060329020304865866, 
    0.06034780102727743, 0.060362669286068801, 0.060373673442856324, 
    0.060380881085646577, 0.060384380344181275, 0.06038427462148991, 
    0.06038068766513504, 0.060373761586417503, 0.060363646235558809, 
    0.060350496948930972, 0.060334460492093879, 0.060315665562081448, 
    0.060294209625794605, 0.060270154715086913, 0.060243531930943887, 
    0.060214341665659143, 0.060182562800084258, 0.060148159665078867, 
    0.060111103234631855, 0.06007136609960443, 0.060028935483917502, 
    0.059983816156120424, 0.059936025390755543, 0.05988559646322679, 
    0.059832578247278369, 0.059777033597019441, 0.059719041637952962, 
    0.059658704726075311, 0.059596146254796152, 0.059531522945375837, 
    0.059465015114943717, 0.059396838737814456, 0.059327238171427377, 
    0.059256475399310185, 0.059184824359697394, 0.059112552826645265, 
    0.059039916396330883, 0.058967150333182325, 0.058894447135532074, 
    0.058821955236653962, 0.058749771220933888, 0.058677931269343245, 
    0.058606408336859248, 0.058535115837951818, 0.058463901928036681, 
    0.058392562172522401, 0.058320849081052381, 0.058248487278810428, 
    0.058175187847413712, 0.058100664440117029, 0.058024657209006875, 
    0.057946946358348871, 0.057867369053289167, 0.057785821919540785, 
    0.05770227798280881, 0.057616787220747812, 0.057529475908686546, 
    0.057440538836925355, 0.057350211333263908, 0.057258762997185006, 
    0.057166455535676917, 0.05707351090594915, 0.056980118598766269, 
    0.056886417090980627, 0.0567925007292489, 0.056698428792842558, 
    0.056604244723409365, 0.056509983517343994, 0.056415695955350793, 
    0.056321445861064974, 0.056227320813187723, 0.05613342469495837, 
    0.056039866956500081, 0.055946755295323551, 0.055854168025721698, 
    0.055762129896248659, 0.055670596139466004, 0.055579425879075453, 
    0.055488370599260164, 0.055397069352491252, 0.055305063586003622, 
    0.055211807662467721, 0.055116710157221416, 0.055019170384776696, 
    0.054918628181847076, 0.054814595278372139, 0.054706666532191091, 
    0.054594539856491611, 0.05447799885477253, 0.054356902265730804, 
    0.05423117874543823, 0.05410079300899618, 0.0539657294009359, 
    0.05382598229675991, 0.053681532997875585, 0.05353232272528647, 
    0.053378252833101242, 0.053219174604534229, 0.053054899599372062, 
    0.052885201564778279, 0.052709853997506606, 0.052528653672431105, 
    0.052341451036932739, 0.052148176494289461, 0.051948849521712206, 
    0.05174359337339976, 0.051532601200108503, 0.051316146672773302, 
    0.051094525953162807, 0.050868079531380068, 0.050637148086262962, 
    0.050402103217515828, 0.05016332069640568, 0.04992119195717562, 
    0.049676115189346635, 0.049428516983490586, 0.049178809998681801, 
    0.048927421300386582, 0.048674765482179055, 0.048421233463290282, 
    0.04816719373242527, 0.047912972445006786, 0.047658840249985693, 
    0.047405014498398408, 0.047151642111636756, 0.046898774674587147, 
    0.046646400092751221, 0.046394391023977903, 0.046142522097695024, 
    0.045890446233603645, 0.04563770140736273, 0.045383726778723286, 
    0.045127875902556527, 0.044869464321815183, 0.044607822810198434, 
    0.044342349820917615, 0.044072580210268206, 0.04379822157004884, 
    0.043519219527132051, 0.043235781837831715, 0.042948422356891384, 
    0.042657949099458026, 0.042365469689748948, 0.042072349273875265, 
    0.041780157139230514, 0.041490598747526454, 0.041205456071318904, 
    0.040926537629314877, 0.04065560781943027, 0.040394358014661652, 
    0.040144384410701298, 0.039907146171380484, 0.039683977592739401, 
    0.039476062519950776, 0.039284448385097662, 0.039110052947695227, 
    0.038953645775668455, 0.038815859920672942, 0.038697175499821337, 
    0.038597914720312557, 0.038518190562577902, 0.038457899901368733, 
    0.038416694959630363, 0.038393961173350054, 0.038388825073036197, 
    0.038400143162084281, 0.038426517316710006, 0.038466339325072658, 
    0.03851783037203383, 0.038579109480584323, 0.03864823135851931, 
    0.038723262879960828, 0.0388023042960777, 0.038883579107167408, 
    0.038965449335966809, 0.03904641597491422, 0.039125226824585926, 
    0.039200780674352592, 0.039272226132420436, 0.039338874474055402, 
    0.039400206061491624, 0.039455827915702651, 0.039505434323618235, 
    0.039548790399330319, 0.039585667341489869, 0.039615902301079739, 
    0.039639390017175764, 0.039656161727732987, 0.039666381216839471, 
    0.039670399149400327, 0.039668709409566315, 0.03966198416197448, 
    0.039650995650231932, 0.039636584737679698, 0.039619625082935428, 
    0.039600965170790939, 0.039581418018302165, 0.039561699668672075, 
    0.039542481631678825, 0.039524404064815812, 0.039508091199917716, 
    0.039494184684316286, 0.039483313865547792, 0.03947608076892855, 
    0.039473018599609846, 0.039474527740769615, 0.039480923653701934, 
    0.039492459399181064, 0.039509366380459869, 0.039531910618627514, 
    0.039560403790019218, 0.039595242838002573, 0.039636910862529469, 
    0.039685904544034277, 0.039742818095635242, 0.039808080576058807, 
    0.039882159719303728, 0.039965164917903973, 0.040056815748194731, 
    0.040156755333129762, 0.040264002359202793, 0.040377427903482109, 
    0.040495539845685713, 0.04061642156790389,
  // Fqt-total(1, 0-1999)
    0.99999999999999956, 0.99955255870496751, 0.99821416445889921, 
    0.99599647490078835, 0.9929185774998438, 0.98900653212994838, 
    0.98429276641126995, 0.97881535848777246, 0.97261723754647611, 
    0.96574533668919105, 0.95824973051199269, 0.95018278252767951, 
    0.94159832654224052, 0.93255090009012565, 0.92309504150021904, 
    0.91328465835919459, 0.90317247079376173, 0.89280953543905184, 
    0.88224483851799496, 0.87152496647426136, 0.86069384240921187, 
    0.84979252868998256, 0.8388590938713183, 0.82792853318184956, 
    0.81703274816995508, 0.80620056628057335, 0.79545779980833586, 
    0.78482733702564922, 0.77432925120709239, 0.7639809304849583, 
    0.75379722696094886, 0.74379061076068353, 0.73397134098036476, 
    0.72434763231321464, 0.71492582451333264, 0.70571054729447058, 
    0.69670488139922648, 0.68791051300721506, 0.67932788262575639, 
    0.67095632840172292, 0.6627942193828531, 0.65483908819251235, 
    0.64708775020692633, 0.63953642074412298, 0.63218081842481222, 
    0.62501626179308123, 0.61803775089817392, 0.61124004362361761, 
    0.60461772026063554, 0.59816524180353325, 0.5918769952808266, 
    0.58574734101977854, 0.57977064640961595, 0.57394131975111096, 
    0.56825383207507096, 0.5627027417010797, 0.55728270600028695, 
    0.5519884932871808, 0.54681499153620061, 0.54175721584146608, 
    0.5368103080189458, 0.53196953940142633, 0.52723031324004499, 
    0.52258815889752908, 0.51803873893967123, 0.51357785045859727, 
    0.50920143312120558, 0.50490557971072547, 0.5006865463021607, 
    0.49654076026637467, 0.49246482341058317, 0.48845551141555094, 
    0.48450976858202566, 0.48062469598655311, 0.476797540571961, 
    0.47302568335369349, 0.46930662883110019, 0.46563799516948284, 
    0.46201750552702053, 0.45844298750400331, 0.45491236591883405, 
    0.45142366581859672, 0.44797501144604257, 0.44456463088861031, 
    0.44119085932905566, 0.43785214740271372, 0.43454706470453081, 
    0.43127431033043484, 0.42803271793905856, 0.42482125247543301, 
    0.42163901147149102, 0.41848521749743178, 0.41535920976675067, 
    0.41226043762484499, 0.40918845700137069, 0.40614292991449513, 
    0.40312362061348783, 0.40013039311575155, 0.39716320291125695, 
    0.39422208736600794, 0.39130715060437338, 0.38841855098335099, 
    0.38555648404680126, 0.38272116944286072, 0.3799128392713399, 
    0.37713172731932199, 0.3743780572240869, 0.37165203615060999, 
    0.36895385083966292, 0.36628366053056477, 0.36364159880033398, 
    0.36102777111269696, 0.35844226045369498, 0.35588512553675095, 
    0.35335640668716717, 0.35085612333863697, 0.34838427220906493, 
    0.34594082299830975, 0.34352571867696502, 0.3411388730725094, 
    0.3387801739150107, 0.33644948882655712, 0.33414667026813555, 
    0.33187156239257753, 0.32962400186706831, 0.32740381871135665, 
    0.32521083499539244, 0.32304486144025901, 0.32090569206674141, 
    0.31879309969550668, 0.31670683378185704, 0.31464662403673627, 
    0.31261218090380988, 0.31060319973454797, 0.30861936014609703, 
    0.30666032702308577, 0.30472574914066408, 0.30281525335986714, 
    0.3009284451801531, 0.29906490697425486, 0.29722419874233452, 
    0.29540585771135741, 0.29360939851831136, 0.2918343114202771, 
    0.29008006466781272, 0.28834609918415044, 0.28663183017463495, 
    0.28493664368762639, 0.28325989523238643, 0.2816009068805419, 
    0.27995896807010689, 0.2783333382584694, 0.27672325121803637, 
    0.27512792394819996, 0.27354656515332426, 0.27197839337709423, 
    0.27042264618388862, 0.26887859709388168, 0.26734556379818469, 
    0.26582292052175488, 0.26431010082853718, 0.26280660113626503, 
    0.26131197860740607, 0.25982584825835225, 0.25834787616279881, 
    0.25687777136058604, 0.25541527766500227, 0.25396016510685449, 
    0.25251222335068041, 0.25107125590729468, 0.24963707831327481, 
    0.24820951928094506, 0.24678842189853503, 0.24537364213408203, 
    0.24396504835076474, 0.24256251843848062, 0.24116593926580779, 
    0.2397752008919444, 0.23839019752070997, 0.23701082666193671, 
    0.23563698693446031, 0.23426858151823421, 0.23290551802350987, 
    0.23154770990703602, 0.23019507537144096, 0.22884753724750173, 
    0.2275050169605978, 0.22616743466741121, 0.22483470627726757, 
    0.22350674149192826, 0.2221834438048601, 0.22086471506083899, 
    0.21955045881504301, 0.21824058094197554, 0.21693499620508727, 
    0.21563363301957675, 0.21433643166246155, 0.21304335108392811, 
    0.21175436242201745, 0.21046945002262343, 0.20918860454922192, 
    0.2079118254165869, 0.20663911608046964, 0.20537049104957561, 
    0.20410596993382865, 0.20284558475763872, 0.20158937651955247, 
    0.20033739921734778, 0.19908971803862635, 0.19784640754688743, 
    0.19660755446138684, 0.19537325406036568, 0.19414361161967519, 
    0.19291874211658555, 0.19169877128279789, 0.19048383952993728, 
    0.18927410134525158, 0.18806972840841574, 0.18687090851062951, 
    0.18567784445165095, 0.18449074910261321, 0.18330984014315499, 
    0.1821353355411707, 0.18096744454411987, 0.17980636313710047, 
    0.17865227008860723, 0.17750532182003392, 0.17636565255062045, 
    0.17523337284139218, 0.17410856940603842, 0.1729913079864859, 
    0.17188163199115566, 0.17077956303299552, 0.16968510369432946, 
    0.16859823656609946, 0.16751892420856329, 0.16644710740746488, 
    0.16538270509823597, 0.16432561195239478, 0.16327569459979921, 
    0.16223279744567182, 0.16119674029577291, 0.16016732804078013, 
    0.15914435363079968, 0.15812761281979193, 0.15711690908205744, 
    0.15611206728272747, 0.15511293678775831, 0.15411940227247337, 
    0.15313138738238852, 0.1521488575587355, 0.15117182139115176, 
    0.15020032710543754, 0.14923446261094767, 0.14827435268540629, 
    0.14732016000551365, 0.14637208333205268, 0.14543036130313269, 
    0.14449526753506764, 0.143567109417299, 0.14264622099327304, 
    0.14173295694107385, 0.14082768002646903, 0.13993074821844317, 
    0.13904250199213536, 0.13816325371951046, 0.13729326966223482, 
    0.13643276643466348, 0.13558190210043419, 0.13474077385415736, 
    0.13390941934319875, 0.13308781939877351, 0.1322759062921946, 
    0.13147357340338897, 0.1306806828448539, 0.1298970797020339, 
    0.12912260249625507, 0.12835709027930714, 0.12760038965560533, 
    0.12685236033944999, 0.12611287475134408, 0.12538181771776322, 
    0.12465908618332801, 0.1239445853713645, 0.12323822792948334, 
    0.12253993248364721, 0.12184962259984558, 0.12116722766252983, 
    0.1204926829457488, 0.11982593082327402, 0.11916692237895572, 
    0.11851561768058959, 0.11787198662509607, 0.11723600624801729, 
    0.11660766379209458, 0.11598695610872878, 0.11537389212540634, 
    0.11476849287540876, 0.11417079170050191, 0.11358083387961564, 
    0.11299867171648301, 0.11242436158561686, 0.11185795794624857, 
    0.11129951091368302, 0.11074905676379812, 0.11020661786484441, 
    0.10967219651591745, 0.10914577164101898, 0.10862729594625038, 
    0.10811669603619302, 0.10761387450012369, 0.10711871376292907, 
    0.10663108458954737, 0.10615085670154874, 0.10567790682093989, 
    0.10521212916632425, 0.10475344257466961, 0.10430179478846144, 
    0.10385716516102016, 0.10341956372269677, 0.10298902963052424, 
    0.10256562443909394, 0.10214942785389504, 0.10174053050559501, 
    0.10133902616473107, 0.10094500605871039, 0.10055855278746653, 
    0.10017973718091333, 0.099808612374886377, 0.099445214249597028, 
    0.099089557472922848, 0.098741636272780486, 0.09840142456662368, 
    0.098068876226533111, 0.097743926182606175, 0.097426491482279776, 
    0.097116470332530042, 0.096813744468155008, 0.096518177905020333, 
    0.09622961828595028, 0.095947897549574293, 0.095672832502539384, 
    0.095404225736406639, 0.095141868288045647, 0.094885535588841455, 
    0.09463499140994952, 0.094389980661981218, 0.094150227422443458, 
    0.093915427274998478, 0.093685240448330473, 0.093459289188508779, 
    0.093237156608628843, 0.093018382686062745, 0.092802467049803716, 
    0.092588870575009238, 0.092377016547860499, 0.092166291742285786, 
    0.091956054117051392, 0.091745640139279605, 0.091534376095523354, 
    0.091321592383695277, 0.091106632442024882, 0.090888866140798094, 
    0.090667702236610234, 0.090442601361339331, 0.090213088181220938, 
    0.089978760495659046, 0.089739297537526796, 0.089494462938064401, 
    0.089244103037828842, 0.088988144910816941, 0.088726585988655321, 
    0.088459490861725582, 0.088186979168930715, 0.087909220904580726, 
    0.087626428630587547, 0.087338851246877139, 0.087046767567294014, 
    0.086750482094028233, 0.086450316603635044, 0.086146604171939908, 
    0.085839685612906433, 0.085529900806964737, 0.085217586853400099, 
    0.084903074850651503, 0.08458668886213315, 0.084268748873334465, 
    0.083949567315206988, 0.083629455296458377, 0.083308720632749883, 
    0.082987665897299986, 0.082666585603595508, 0.082345764105105829, 
    0.08202547372197172, 0.081705977972384936, 0.081387531976069585, 
    0.081070387690126561, 0.080754793221006413, 0.080440995388679062, 
    0.080129241796240203, 0.079819780284817093, 0.079512859940890843, 
    0.079208727806311066, 0.078907625962266234, 0.078609782830480035, 
    0.07831540511371346, 0.078024664982121031, 0.077737693802465355, 
    0.077454570391336672, 0.077175315957272464, 0.076899889225332752, 
    0.076628183865594099, 0.076360028876124753, 0.076095195384473485, 
    0.075833398626560036, 0.07557430896190552, 0.075317559253140723, 
    0.075062752521001475, 0.074809474303587087, 0.074557300358434497, 
    0.07430581031920229, 0.074054596289835392, 0.073803271042567065, 
    0.073551477869105958, 0.073298897430073548, 0.073045253597509685, 
    0.07279032016924207, 0.072533925519470036, 0.072275957468880436, 
    0.072016370283850842, 0.071755186520693598, 0.071492501184457227, 
    0.07122847723549397, 0.070963342334864732, 0.070697381588864516, 
    0.070430926236209446, 0.070164338737054785, 0.069898003461185423, 
    0.069632310714236367, 0.069367642311590705, 0.069104357069442499, 
    0.068842776135331657, 0.068583168487025142, 0.06832574047779176, 
    0.068070622008352483, 0.067817857557278538, 0.067567401497482596, 
    0.067319109951993431, 0.067072743559981648, 0.066827967649354891, 
    0.066584363781794442, 0.066341444131426203, 0.066098669391127435, 
    0.065855470700363405, 0.065611267992099181, 0.065365485641974266, 
    0.06511756656325221, 0.064866978816641094, 0.064613225688046561, 
    0.064355850102744958, 0.064094440770042949, 0.063828636304502848, 
    0.063558130932756154, 0.063282677383301247, 0.06300209659625719, 
    0.062716280902798266, 0.062425201168631247, 0.062128908070026558, 
    0.061827530041574826, 0.061521273342246802, 0.061210413913277244, 
    0.06089529258280315, 0.060576304379777922, 0.060253893137051054, 
    0.059928544343365996, 0.059600777504831684, 0.05927114341102642, 
    0.058940218571688699, 0.058608605039356651, 0.058276921610795118, 
    0.0579458054902907, 0.057615902290526919, 0.057287864331937388, 
    0.056962343920342405, 0.056639988329434302, 0.056321430405677081, 
    0.056007281347647653, 0.055698120263603212, 0.055394484171642111, 
    0.055096856725636169, 0.054805655703753044, 0.054521227883618781, 
    0.054243839392319332, 0.053973671076954916, 0.053710822082145671, 
    0.053455312628985105, 0.053207088785199613, 0.052966030241171948, 
    0.052731953217346056, 0.052504612558714435, 0.052283702471451726, 
    0.052068858630232827, 0.051859659838953895, 0.051655629561922434, 
    0.051456241957338313, 0.051260928850912144, 0.051069090858869355, 
    0.05088011252461902, 0.050693375890284269, 0.050508278311666203, 
    0.050324244562335099, 0.050140740346534665, 0.049957279651184135, 
    0.049773431583398184, 0.049588825713670126, 0.049403151755212621, 
    0.049216156582838851, 0.04902764221244249, 0.04883746151515983, 
    0.048645512351319864, 0.048451734756215933, 0.048256105942462685, 
    0.048058639148369622, 0.04785938018102668, 0.047658408309551099, 
    0.047455832905570289, 0.047251792030923834, 0.047046448816580336, 
    0.046839984292165376, 0.046632595452959551, 0.046424488511660054, 
    0.046215878807028439, 0.046006988646318893, 0.045798049255432564, 
    0.045589298273203058, 0.045380981657750064, 0.045173347453795996, 
    0.044966650412305749, 0.044761145748221993, 0.044557092943556358, 
    0.044354757333962679, 0.044154413983709478, 0.043956348635386978, 
    0.043760864554113203, 0.043568280036844625, 0.043378928571740638, 
    0.043193156041987167, 0.043011313758587667, 0.042833752928112118, 
    0.042660814498568102, 0.04249282074646283, 0.042330062029083355, 
    0.042172784327615793, 0.042021181370071568, 0.041875381106359369, 
    0.041735441024813552, 0.041601344046303744, 0.041472996757567701, 
    0.04135023559719031, 0.041232831030681052, 0.041120498997496646, 
    0.04101290547701477, 0.04090967712949832, 0.040810404529001462, 
    0.040714653642089288, 0.04062196976440164, 0.040531890911583601, 
    0.040443955027487433, 0.040357714115241743, 0.040272741099584342, 
    0.040188638643723587, 0.040105042428671842, 0.040021625329071185, 
    0.039938099439581487, 0.039854215515004954, 0.039769761445435502, 
    0.039684560051141828, 0.03959846880759281, 0.039511372212508208, 
    0.039423181324030179, 0.03933382844465156, 0.039243264498138475, 
    0.039151459477640455, 0.039058399372489415, 0.038964085863903354, 
    0.038868535129747153, 0.038771777428963553, 0.038673852168826253, 
    0.038574805863832495, 0.038474686967756612, 0.038373543181300415, 
    0.038271420111998813, 0.038168355600458344, 0.038064379109910625, 
    0.037959509917347874, 0.037853753584029898, 0.037747106363084725, 
    0.037639552408890838, 0.037531068090041121, 0.037421623960825441, 
    0.037311186123163982, 0.037199721693637472, 0.037087198819967665, 
    0.03697358852234827, 0.036858867657428421, 0.036743020128530521, 
    0.03662603952049643, 0.036507931411809275, 0.036388713956042588, 
    0.036268424173261669, 0.036147111136268908, 0.036024843645253012, 
    0.035901704143534843, 0.035777785002547573, 0.03565318574553418, 
    0.035528008918608495, 0.035402354334684756, 0.035276317414182974, 
    0.035149983761107569, 0.035023428440766058, 0.034896709946726306, 
    0.034769869588606041, 0.034642924230293484, 0.034515861999243343, 
    0.034388635084357515, 0.034261151881277804, 0.034133274190534399, 
    0.034004815359582281, 0.033875539165005866, 0.033745164671886173, 
    0.033613372939223146, 0.033479811334952009, 0.033344102603055543, 
    0.033205857048353757, 0.03306468063901305, 0.032920188761900754, 
    0.032772016265694544, 0.032619831486418907, 0.032463343577396435, 
    0.032302313980924535, 0.032136563209077026, 0.031965976552611033, 
    0.031790510250193506, 0.031610193682030593, 0.031425130412989305, 
    0.03123549763329447, 0.031041542741216139, 0.030843577257047405, 
    0.030641968537196758, 0.030437130186527425, 0.030229512311253176, 
    0.03001958667793396, 0.029807838502413034, 0.029594753611211638, 
    0.029380809285342462, 0.029166467876763458, 0.028952169275008134, 
    0.028738322927515769, 0.028525302038023378, 0.028313435575050908, 
    0.028102997545688266, 0.027894199453975539, 0.027687185837409405, 
    0.02748203932123713, 0.027278787822630785, 0.027077416194646129, 
    0.026877880645210458, 0.026680121364721213, 0.026484075038589308, 
    0.026289683257075799, 0.026096898708780108, 0.025905691750113705, 
    0.025716044332046523, 0.025527946968014227, 0.025341389783666589, 
    0.02515635388020512, 0.024972796860929642, 0.024790647261028486, 
    0.024609797073620605, 0.024430091534556723, 0.024251324784783035, 
    0.024073233219462059, 0.02389549463759464, 0.023717725393984444, 
    0.023539484866804437, 0.023360290021963069, 0.023179632074960592, 
    0.022997003805817873, 0.022811925879294124, 0.022623975625379655, 
    0.02243280992790532, 0.022238186637151575, 0.022039978864985783, 
    0.021838176837379517, 0.021632880943850106, 0.021424282615772634, 
    0.021212638918591473, 0.020998251318260948, 0.020781443063663849, 
    0.020562551151560811, 0.020341916277104632, 0.020119875916542025, 
    0.01989675884831078, 0.019672878866477218, 0.019448527853265545, 
    0.019223970235564186, 0.018999441468391779, 0.018775143161179456, 
    0.018551245657270999, 0.018327887464799526, 0.018105180278553991, 
    0.017883212421781158, 0.017662050203260993, 0.017441747732944823, 
    0.017222342298850012, 0.017003862730693646, 0.016786328081644084, 
    0.016569748438311858, 0.016354121545723327, 0.01613943511861924, 
    0.015925662800047074, 0.015712764846001717, 0.015500688576278942, 
    0.015289375080925127, 0.015078763356497575, 0.014868802497376515, 
    0.014659462901989589, 0.014450740731601684, 0.014242663365914031, 
    0.014035290548570892, 0.013828705099902361, 0.013623007116153441, 
    0.01341830293447138, 0.013214699157533221, 0.013012293321840843, 
    0.012811170648262649, 0.012611400757875557, 0.012413037489785467, 
    0.012216118910758111, 0.012020669914239206, 0.011826704488016832, 
    0.011634228208871052, 0.01144323730401671, 0.011253719431161957, 
    0.01106564989396162, 0.010878989279482932, 0.010693680543618495, 
    0.010509648094188388, 0.0103267960885167, 0.010145010463776085, 
    0.0099641577244867462, 0.0097840850918992656, 0.0096046216604747294, 
    0.009425573484132227, 0.0092467317954346585, 0.009067869008123881, 
    0.0088887472732076846, 0.0087091197613117718, 0.0085287352265776672, 
    0.008347344388602301, 0.0081647018112726549, 0.0079805705451907009, 
    0.0077947249957530124, 0.0076069545318142914, 0.0074170652285325519, 
    0.007224884538830161, 0.0070302627508688305, 0.0068330729730169387, 
    0.006633216096924883, 0.0064306190456920407, 0.0062252351516073837, 
    0.0060170484100639087, 0.0058060729392913546, 0.0055923554198782427, 
    0.0053759801846260278, 0.0051570657555731775, 0.0049357740711323001, 
    0.0047123065862248129, 0.0044869054169732253, 0.0042598497943839141, 
    0.0040314511820611623, 0.0038020503361352186, 0.0035720056811673851, 
    0.0033416902923434021, 0.0031114799299036379, 0.0028817482235118015, 
    0.0026528579179305235, 0.0024251496495560749, 0.0021989388991064127, 
    0.0019745101877909088, 0.0017521153323696085, 0.0015319707062147439, 
    0.0013142632845810484, 0.0010991533833365462, 0.00088678027043771204, 
    0.00067726557928896134, 0.00047071924928736509, 0.00026723564870560014, 
    6.6893211202166987e-05, -0.00013024785764536567, -0.00032414854775402369, 
    -0.00051479581090463507, -0.00070220104019135107, 
    -0.00088640218390759456, -0.0010674613821383451, -0.0012454677685204971, 
    -0.0014205363579688072, -0.0015928086416738796, -0.0017624541230059773, 
    -0.0019296720478005867, -0.002094694241177432, -0.0022577838953615429, 
    -0.0024192372569321026, -0.0025793801289722843, -0.0027385682819643575, 
    -0.0028971789031032916, -0.0030556089026325568, -0.0032142684981833185, 
    -0.0033735755051117382, -0.0035339442990804412, -0.0036957792214759922, 
    -0.0038594586908814806, -0.0040253255173870791, -0.0041936712945536431, 
    -0.0043647256444963771, -0.0045386504582529963, -0.0047155381457859059, 
    -0.0048954150640504205, -0.0050782452669625297, -0.0052639447319409198, 
    -0.0054523855274445513, -0.0056434105247475793, -0.0058368383659321912, 
    -0.0060324716140335195, -0.0062301025201893087, -0.0064295149346060738, 
    -0.0066304870574265167, -0.006832791990879261, -0.0070362041387855663, 
    -0.0072405003928231078, -0.0074454632294966242, -0.0076508880335868727, 
    -0.0078565837289904759, -0.0080623808163587298, -0.0082681306551693305, 
    -0.0084737124776627822, -0.0086790341000864447, -0.0088840351564344611, 
    -0.0090886884753738576, -0.0092930010923363681, -0.0094970128500623825, 
    -0.0097007981831248435, -0.0099044595922465391, -0.01010812378410181, 
    -0.010311931348939259, -0.010516028939206017, -0.010720555701133828, 
    -0.010925636265616904, -0.011131369299158811, -0.011337819915812708, 
    -0.011545014557477539, -0.011752934541004248, -0.011961519007335077, 
    -0.012170659135514912, -0.012380207339221651, -0.012589978481476739, 
    -0.012799756751012676, -0.013009306738299135, -0.013218378150448075, 
    -0.013426719182378007, -0.013634082187945793, -0.013840231319310498, 
    -0.014044949052784672, -0.014248041402691838, -0.014449337869145042, 
    -0.014648692562119802, -0.01484598541060045, -0.015041119337031785, 
    -0.015234017093040878, -0.015424618659603101, -0.015612876079603809, 
    -0.015798747441043731, -0.015982187614792382, -0.016163140643036766, 
    -0.01634153094202756, -0.016517252009171039, -0.016690159755700488, 
    -0.016860066729247804, -0.01702673675554953, -0.017189886333856676, 
    -0.017349184828670042, -0.017504262499756573, -0.01765471729037894, 
    -0.017800124160913807, -0.017940047019246525, -0.018074047238805374, 
    -0.018201694529772931, -0.018322576259891799, -0.018436302582212096, 
    -0.018542514226808651, -0.018640888351080569, -0.018731140419945624, 
    -0.018813030590534685, -0.018886362551971007, -0.01895098614696129, 
    -0.019006795038085497, -0.019053725709449385, -0.019091756197386574, 
    -0.019120905013157732, -0.019141227862040644, -0.019152821884038825, 
    -0.019155827288474661, -0.01915042933848107, -0.019136855157971359, 
    -0.019115372716997162, -0.019086284641730962, -0.019049924842160122, 
    -0.019006651737761875, -0.018956847441922057, -0.018900913245186272, 
    -0.018839266827430902, -0.018772338405505594, -0.018700566588612706, 
    -0.018624394513298309, -0.018544264458592582, -0.018460616856185674, 
    -0.01837388482238584, -0.018284493950283739, -0.018192861826043606, 
    -0.018099397446478125, -0.01800449741653647, -0.017908548985542762, 
    -0.017811928732577694, -0.017714997343870137, -0.017618098320552271, 
    -0.017521553730989615, -0.01742565914143827, -0.017330677318323363, 
    -0.017236836573634031, -0.017144328290250262, -0.01705330431562594, 
    -0.016963883811851876, -0.016876152182562873, -0.016790164176380143, 
    -0.016705950262747331, -0.016623511955123956, -0.016542829096085034, 
    -0.016463860921899293, -0.016386550904160021, -0.016310830255188584, 
    -0.01623662136707503, -0.016163840232853041, -0.01609240018656408, 
    -0.016022209129360823, -0.015953171219478587, -0.015885187626046765, 
    -0.015818155559794597, -0.015751968917402277, -0.01568651925827836, 
    -0.015621700515774398, -0.015557410816351954, -0.015493555791624099, 
    -0.015430053756468446, -0.01536683937504002, -0.015303868080479359, 
    -0.015241117939165709, -0.015178590399631705, -0.015116313004381522, 
    -0.015054336567174014, -0.014992734704597012, -0.01493160265255093, 
    -0.01487105046907157, -0.014811202314777852, -0.014752190411433283, 
    -0.014694151360773153, -0.014637222491853393, -0.014581537943767764, 
    -0.014527225834239196, -0.014474404220655252, -0.014423174608688569, 
    -0.014373621407457945, -0.014325803483378868, -0.014279753352689131, 
    -0.014235471815968846, -0.014192928938409604, -0.014152064238864562, 
    -0.014112788312346355, -0.014074990855317125, -0.014038546082537786, 
    -0.014003320492744043, -0.013969184178797179, -0.013936014026667351, 
    -0.013903705760614067, -0.013872177978265291, -0.013841375440732112, 
    -0.013811271219271337, -0.013781865797410611, -0.013753184185284194, 
    -0.013725271426822517, -0.013698191040188962, -0.013672017360256266, 
    -0.013646836916825502, -0.013622742690094263, -0.013599831895692567, 
    -0.013578203843171922, -0.013557952892146114, -0.013539165869456684, 
    -0.013521916724933832, -0.013506261810101202, -0.013492238600456808, 
    -0.01347986542539808, -0.013469146858790148, -0.013460086662775348, 
    -0.013452695601728338, -0.01344700946916504, -0.013443100744738059, 
    -0.013441090534792028, -0.013441157213896878, -0.013443535726844195, 
    -0.013448517970571896, -0.013456441587568282, -0.013467678398772867, 
    -0.013482621078226616, -0.013501667966759359, -0.013525209796813603, 
    -0.013553620103070419, -0.013587248127016106, -0.013626417013355705, 
    -0.013671419854962499, -0.013722519536038799, -0.013779950266242248, 
    -0.013843912201137398, -0.013914568891995044, -0.013992040446191836, 
    -0.014076397795415177, -0.014167651836439031, -0.014265745110431265, 
    -0.014370545897231444, -0.014481842392117243, -0.0145993406126298, 
    -0.014722667335353819, -0.014851374889503553, -0.014984944027691554, 
    -0.015122794987687897, -0.015264290478901266, -0.015408747857715933, 
    -0.015555447886951356, -0.015703649298819046, -0.015852602962421476, 
    -0.016001566346571454, -0.016149822735108257, -0.016296697339525996, 
    -0.016441571230075169, -0.016583893128654426, -0.016723192831244925, 
    -0.016859086582312575, -0.016991283430329712, -0.017119584960416604, 
    -0.017243877751250653, -0.017364129345010186, -0.017480373646645338, 
    -0.017592700608002394, -0.017701245926827439, -0.017806183266818019, 
    -0.017907721026556765, -0.01800609618452477, -0.018101572263260524, 
    -0.018194432196653607, -0.018284969298066455, -0.018373477847295767, 
    -0.01846024074407256, -0.018545516515681947, -0.018629529377533767, 
    -0.018712458228814254, -0.018794429615385001, -0.018875512197964142, 
    -0.018955712427208244, -0.019034975702217481, -0.019113188387596652, 
    -0.019190185076618078, -0.01926575295002118, -0.01933964452580015, 
    -0.019411583166173578, -0.01948127089368543, -0.019548397243445197, 
    -0.019612642571072883, -0.019673681849587888, -0.019731190305536085, 
    -0.019784846964249019, -0.019834340581471759, -0.01987937646624191, 
    -0.019919686053853608, -0.019955029804697193, -0.019985211305270267, 
    -0.020010076958369406, -0.020029524168978987, -0.0200435013427883, 
    -0.020052005864912043, -0.020055084381564371, -0.020052826020150627, 
    -0.020045362493899776, -0.020032862470737194, -0.020015527233522779, 
    -0.019993583231266619, -0.019967278657773167, -0.019936872471962727, 
    -0.019902628292400752, -0.019864805038736669, -0.019823651709057071, 
    -0.019779399624809419, -0.019732257873216433, -0.019682409324359464, 
    -0.019630006377995456, -0.019575169017732541, -0.019517982525934705, 
    -0.019458497266088223, -0.01939672806526881, -0.019332652877625443, 
    -0.01926621569645777, -0.019197328807117723, -0.019125879293525799, 
    -0.019051733295862371, -0.018974743021385312, -0.018894754686592775, 
    -0.018811616019878269, -0.018725183166575721, -0.018635328507737026, 
    -0.018541944740266991, -0.018444950704635497, -0.018344295381852126, 
    -0.018239961377519157, -0.018131965033638349, -0.018020359822729735, 
    -0.017905233622429857, -0.017786708548850162, -0.017664935363302596, 
    -0.01754009217615473, -0.01741237485743069, -0.017281993512880432, 
    -0.017149164835630767, -0.017014107189602196, -0.016877035571918254, 
    -0.01673815914426378, -0.016597678854206623, -0.016455788103283603, 
    -0.016312674566513849, -0.016168520841043237, -0.016023510200714894, 
    -0.015877828361414884, -0.015731666410332659, -0.015585223320292177, 
    -0.015438706756623065, -0.015292333437283215, -0.015146328438972156, 
    -0.01500092297940196, -0.014856353988186171, -0.014712862507034918, 
    -0.014570692937154186, -0.014430090832343591, -0.014291302574316338, 
    -0.014154574367679378, -0.014020153894319173, -0.013888288082383748, 
    -0.013759226773828771, -0.013633219088775425, -0.01351051515898479, 
    -0.013391365583631321, -0.013276013853713757, -0.013164691596432514, 
    -0.013057616152520254, -0.012954977693148904, -0.012856936574460453, 
    -0.012763617483035661, -0.012675106137082236, -0.012591450145393795, 
    -0.01251265489316231, -0.012438688605607149, -0.01236947369605006, 
    -0.012304890004342968, -0.012244772215095082, -0.012188902368256153, 
    -0.012137013888721982, -0.012088788606858769, -0.01204386110760017, 
    -0.0120018254604604, -0.011962242445048055, -0.011924654245673029, 
    -0.011888593396130709, -0.011853598414989333, -0.011819221536793538, 
    -0.011785040775618727, -0.011750663176017095, -0.011715731337032449, 
    -0.011679921546562696, -0.011642943112163443, -0.011604533271638368, 
    -0.011564454043720647, -0.011522486137830898, -0.01147842640537206, 
    -0.011432084385671039, -0.01138328371034013, -0.011331863735409209, 
    -0.011277687695747166, -0.011220649610585307, -0.011160685003192032, 
    -0.011097778197965496, -0.011031968954245372, -0.010963355230255486, 
    -0.010892091645579846, -0.010818384836385704, -0.010742484494018835, 
    -0.010664671093175789, -0.01058524370516916, -0.010504510672286756, 
    -0.010422773345388409, -0.010340317119234169, -0.010257405171967816, 
    -0.010174266941446743, -0.010091098748965964, -0.010008057686116324, 
    -0.0099252626823071507, -0.0098427938445912067, -0.0097606936023919965, 
    -0.0096789652913252741, -0.009597576792351601, -0.0095164580726390512, 
    -0.0094355056591600046, -0.0093545824659455601, -0.0092735247818776529, 
    -0.0091921455528751507, -0.0091102407817890939, -0.0090275910701365907, 
    -0.0089439731489205573, -0.0088591606814961629, -0.0087729300222835309, 
    -0.008685069494532292, -0.0085953803616094643, -0.0085036849428195595, 
    -0.0084098258191300027, -0.0083136681309420452, -0.0082150970285639474, 
    -0.0081140160873800372, -0.0080103460046190705, -0.0079040226257544709, 
    -0.0077949954373708729, -0.0076832257240087099, -0.007568682599379763, 
    -0.0074513363805598556, -0.0073311582786460688, -0.0072081115637807076, 
    -0.0070821551097655375, -0.0069532432903464305, -0.0068213386520629511, 
    -0.0066864232435980926, -0.0065485086944187679, -0.0064076525987795127, 
    -0.0062639606661196064, -0.0061175979721644182, -0.005968791553877366, 
    -0.0058178349224789674, -0.0056650822671921557, -0.0055109467781642102, 
    -0.005355889114505478, -0.0052004072142634401, -0.0050450191231808973, 
    -0.004890254351683632, -0.0047366451435592004, -0.0045847175957878629, 
    -0.0044349869742913691, -0.0042879491034084711, -0.0041440769033595677, 
    -0.004003817307179169, -0.0038675845309823721, -0.0037357637367402951, 
    -0.0036087061012145564, -0.003486735632749813, -0.0033701526826578065, 
    -0.0032592399864186218, -0.0031542687600031338, -0.00305551146681354, 
    -0.0029632480569745366, -0.0028777750406767345, -0.0027994074005497581, 
    -0.0027284745621945715, -0.0026653129955248817, -0.0026102539305205498, 
    -0.0025636097011730108, -0.0025256622591551254, -0.0024966543384997925, 
    -0.0024767827950493309, -0.0024661976210305124, -0.0024650000947638506, 
    -0.0024732420750218195, -0.0024909246996103022, -0.0025180013383764967, 
    -0.0025543734415799206, -0.0025998934255172875, -0.0026543573290885485, 
    -0.0027175034986479584, -0.0027890114182175262, -0.0028684934226925573, 
    -0.0029554955152667891, -0.0030494918064472797, -0.0031498841154413097, 
    -0.0032560010970211898, -0.0033670991040483911, -0.0034823684387525165, 
    -0.003600938294090025, -0.0037218878275271212, -0.0038442594825900405, 
    -0.0039670721829869931, -0.0040893370099395207, -0.0042100729002417913, 
    -0.004328319571098603, -0.0044431493399645812, -0.0045536766354557666, 
    -0.0046590668480602374, -0.0047585387825284462, -0.004851377382090359, 
    -0.0049369350372164928, -0.0050146427880685797, -0.0050840158072125285, 
    -0.0051446589162160283, -0.0051962645909217307, -0.0052386109445999871, 
    -0.0052715562707134414, -0.0052950305427745467, -0.0053090266192400044, 
    -0.0053135917681843741, -0.0053088187664851591, -0.0052948444171860148, 
    -0.0052718382328414363, -0.0052399987044163543, -0.0051995494266784993, 
    -0.0051507245992560274, -0.0050937629015048074, -0.0050288952767678389, 
    -0.0049563407784090664, -0.0048762926361879122, -0.0047889187855275142, 
    -0.0046943563313163296, -0.0045927107478649105, -0.0044840619009824728, 
    -0.0043684717258716055, -0.0042459857583915777, -0.0041166444545553517, 
    -0.0039804907577906624, -0.0038375695807816405, -0.0036879303228011138, 
    -0.0035316252034157496, -0.0033687109868897453, -0.0031992441847402521, 
    -0.0030232851860538365, -0.0028408963586150559, -0.0026521526310888353, 
    -0.0024571435706375734, -0.0022559824519453255, -0.0020488160719821439, 
    -0.0018358291448895116, -0.0016172441225165959, -0.0013933241042782592, 
    -0.0011643659140160821, -0.00093069341317930621, -0.0006926533593291399, 
    -0.00045060734168397252, -0.00020493004403710158, 4.3990629113575407e-05, 
    0.00029575436899648833, 0.00054994716451040569, 0.00080613323292387832, 
    0.001063854343046521, 0.0013226210030661202, 0.0015819109154248693, 
    0.0018411674055511362, 0.0020997953705733999, 0.0023571742397308854, 
    0.00261265871552956, 0.0028655898981419328, 0.0031152982298185386, 
    0.0033611121541539967, 0.0036023578121083962, 0.0038383695963196277, 
    0.0040684973965736245, 0.0042921122131007773, 0.0045086200425846412, 
    0.0047174751470294074, 0.0049181899323192894, 0.0051103449992752218, 
    0.0052936002250474701, 0.0054676941594025029, 0.0056324510852807123, 
    0.0057877743978735864, 0.0059336397648536024, 0.0060700852341934773, 
    0.006197204147536035, 0.0063151279763869576, 0.0064240206410291481, 
    0.0065240735630986155, 0.0066154975328127676, 0.0066985269528084595, 
    0.0067734204025156116, 0.0068404702672053138, 0.006900002700814015, 
    0.0069523878174962157, 0.0069980413840607433, 0.0070374237526644005, 
    0.0070710330783364788, 0.0070993983651345847, 0.0071230693728068905, 
    0.0071426051217494619, 0.0071585653987759866, 0.007171507542367235, 
    0.0071819833087542551, 0.0071905369671505888, 0.0071977048739772318, 
    0.0072040204240096687, 0.0072100158734583648, 0.0072162282267437105, 
    0.0072232001276662898, 0.0072314863362856049, 0.0072416572776427242, 
    0.0072542958063400772, 0.0072699935705847216, 0.0072893455987310101, 
    0.0073129382190918243, 0.0073413330911944203, 0.0073750499578348486, 
    0.0074145539435302764, 0.0074602405696704921, 0.0075124252873651105, 
    0.0075713384278053427, 0.007637121634843552, 0.0077098304729108494, 
    0.0077894459276991951, 0.007875879133778102, 0.0079689853235647302, 
    0.0080685791989345227, 0.0081744477296365765, 0.0082863659626226036, 
    0.0084041125068297622, 0.0085274899346769843, 0.0086563385454884456, 
    0.008790551610669382, 0.0089300837385638716, 0.0090749502077772954, 
    0.0092252165974575032, 0.0093809783810771281, 0.0095423423324392451, 
    0.0097094078083141029, 0.0098822577658216511, 0.010060946787716737, 
    0.010245500751790707, 0.01043591551089757, 0.010632152483925905, 
    0.010834141103901693, 0.011041772269170899, 0.011254897700355903, 
    0.011473323834224888, 0.011696809165560129, 0.011925057259584428, 
    0.012157718414452498, 0.012394385749685871, 0.012634597554159478, 
    0.012877843572335113, 0.013123575881568943, 0.013371213119066741, 
    0.013620155449344593, 0.013869794555808624, 0.014119519518612622, 
    0.014368722906078579, 0.01461680465280423, 0.014863171258128935, 
    0.015107235672199576, 0.015348413415303486, 0.01558612740479892, 
    0.015819810055314902, 0.016048909336430398, 0.016272896425292106, 
    0.016491268670491211, 0.016703563247910256, 0.016909355315244345, 
    0.017108278993099964, 0.0173000338139962, 0.017484395496211797, 
    0.017661218637065948, 0.017830441752581201, 0.017992090368736099, 
    0.018146276076350491, 0.018293197374149375, 0.018433134183259769, 
    0.018566440775102628, 0.01869353954597365, 0.018814900170506306, 
    0.018931030691007451, 0.019042453282769628, 0.019149687429740388, 
    0.019253234749948233, 0.019353555915018843, 0.019451066908902959, 
    0.019546133784327929, 0.019639065144067179, 0.01973012077124283, 
    0.01981950258069003, 0.019907353412271411, 0.019993751966333111, 
    0.020078707844919493, 0.020162163904780896, 0.020243996073291186, 
    0.02032402627781563, 0.020402033324032356, 0.020477773376660159, 
    0.020550997600066716, 0.020621467338581854, 0.020688966722019718, 
    0.020753313895508649, 0.020814368305959334, 0.020872034914417321, 
    0.02092626803409256, 0.020977073326954157, 0.021024505178968363, 
    0.021068670445204777, 0.021109721671485192, 0.021147853002945537, 
    0.021183286858680067, 0.021216264751493109, 0.021247024809225981, 
    0.02127578782603708, 0.021302729062830865, 0.021327971347119969, 
    0.021351558942910284, 0.021373446605416308, 0.021393486627501793, 
    0.021411429735118361, 0.02142692627426665, 0.021439528605393193, 
    0.021448705166142581, 0.021453854503126601, 0.021454326294651424, 
    0.021449443644028288, 0.021438516693450704, 0.021420874551209189, 
    0.021395878839079174, 0.021362943535463096, 0.021321544933670066, 
    0.021271228137741186, 0.021211614772938907, 0.02114239921428061, 
    0.021063342500430876, 0.020974266466688547, 0.020875044309997766, 
    0.020765601089474939, 0.020645915338133473, 0.020516036893237461, 
    0.020376103453018872, 0.020226360279123747, 0.020067173594239682, 
    0.019899030971349846, 0.019722536323131402, 0.019538391082247933, 
    0.019347382477603241, 0.019150358164952145, 0.018948209047194787, 
    0.018741840279077087, 0.018532154224301073, 0.01832003482425755, 
    0.0181063276237746, 0.017891831551118131, 0.01767729447308929, 
    0.017463414455809966, 0.017250833240255004, 0.017040139779477458, 
    0.016831855232604959, 0.016626430414166775, 0.016424229911049928, 
    0.016225525523406614, 0.016030488916770558, 0.015839191124237189, 
    0.015651607571024791, 0.015467628054086864, 0.015287078297521975, 
    0.015109739077857913, 0.01493536955231, 0.014763729089107901, 
    0.014594596346549667, 0.014427780984482106, 0.014263131025412419, 
    0.014100538616610101, 0.013939938583434348, 0.01378130175446045, 
    0.013624636461166734, 0.013469990527251478, 0.013317449604778977, 
    0.01316714349760853, 0.0130192469966858, 0.01287397923974979, 
    0.012731596278300377, 0.012592384216384462, 0.012456645965195572, 
    0.012324685428227011, 0.012196795402260357, 0.012073239584579691, 
    0.011954246687583629, 0.011839995527919636, 0.011730620834390004, 
    0.011626208554434142, 0.011526800029222167, 0.011432397445650123, 
    0.0113429719942866, 0.011258469777429286, 0.011178827268986752, 
    0.011103970530029776, 0.011033824633315967, 0.010968291668990215, 
    0.010907228051463476, 0.010850416721617979, 0.010797550240470105, 
    0.010748221381784976, 0.010701936256045557, 0.010658124067845333, 
    0.01061615131419244, 0.01057533962833797, 0.010534976041564888, 
    0.010494333607715109, 0.010452683871830267, 0.010409315633371722, 
    0.010363546917651597, 0.010314730262360416, 0.010262259311895739, 
    0.010205565927997196, 0.010144114467959429, 0.010077395196571623, 
    0.010004929154207422, 0.0099262602778417749, 0.0098409659815772172, 
    0.0097486596462465318, 0.0096490085459474493, 0.009541750297497667, 
    0.0094267023232575721, 0.0093037756090312944, 0.0091729849710251755, 
    0.009034450384831973, 0.0088884057337237973, 0.0087351947151395534, 
    0.0085752781222681786, 0.0084092294837679934, 0.0082377365562595027, 
    0.0080615908461085378, 0.0078816704499127272, 0.0076989092663905479, 
    0.0075142683461556234, 0.0073287061197359008, 0.0071431588071980282, 
    0.0069585344431288944, 0.0067757126902951862, 0.0065955493266191319, 
    0.0064188790664944486, 0.0062465180706399101, 0.0060792636007892331, 
    0.0059178909726208375, 0.0057631414255313431, 0.005615717673792279, 
    0.0054762701571842171, 0.0053453848039366897, 0.0052235780927494604, 
    0.0051112969409537346, 0.005008909035331569, 0.0049167125491442736, 
    0.0048349373317004077, 0.0047637524565182906, 0.0047032716360240522, 
    0.0046535567796101478, 0.0046146329239353159, 0.0045864798068611838, 
    0.0045690371206874129, 0.0045622110717486453, 0.0045658701978377623, 
    0.0045798537419109945, 0.0046039717309354512, 0.004638012318278064, 
    0.0046817404242929551, 0.0047349046338392223, 0.0047972334981166058, 
    0.0048684370094054649, 0.0049482099578007626, 0.0050362315403107948, 
    0.0051321689412513454, 0.0052356910356139465, 0.0053464607585796131, 
    0.0054641547574629089, 0.0055884581002593747, 0.0057190865277501769, 
    0.0058557851267801104, 0.005998348568198213, 0.0061466297129636697, 
    0.0063005412746483464, 0.0064600537767178466, 0.0066251807970250966, 
    0.0067959746563719114, 0.0069725042422226317, 0.0071548263729237539, 
    0.0073429789726834139, 0.0075369458499640269, 0.0077366404586485431, 
    0.0079418966046465519, 0.0081524582014211103, 0.0083679724187520274, 
    0.0085879936234377393, 0.0088119844423156287, 0.0090393263457974188, 
    0.0092693216288194918, 0.009501215600025063, 0.0097342027019908031, 
    0.0099674521901374751, 0.010200125856628944, 0.01043141447468156, 
    0.010660555555250717, 0.010886864043965492, 0.011109743878972424, 
    0.011328710915375425, 0.011543395061608234, 0.011753549237773993, 
    0.011959053750270452, 0.012159928314369585, 0.012356324391050701, 
    0.012548537873816479, 0.012736993978130898, 0.012922242640789804, 
    0.013104946469053299, 0.013285859511941434, 0.013465821166094698, 
    0.013645732256136019, 0.013826555708779692, 0.014009281309897096, 
    0.014194944150678427, 0.014384597965449037, 0.014579302551283816, 
    0.01478012251798585, 0.014988121293532185, 0.015204348888537464, 
    0.015429841485517907, 0.015665608572895413, 0.015912628893664862, 
    0.016171827773642934, 0.01644405937063555, 0.016730088031960764, 
    0.017030556816015369, 0.01734597946187388, 0.017676711598485488, 
    0.018022940598258479, 0.018384666112423946, 0.018761704037270226, 
    0.019153661509244201, 0.019559927326739203, 0.019979665488951043, 
    0.0204118167422776, 0.020855092702115351, 0.021307988659078275, 
    0.021768799147131538, 0.022235653966640432, 0.022706540699499195, 
    0.023179346441238324, 0.023651891417278307, 0.024121955525522026, 
    0.024587312191924275, 0.025045750527752552, 0.025495090629417152, 
    0.025933198746745552, 0.026358001883482546, 0.026767507720649605, 
    0.02715979848624309, 0.027533047808433055, 0.027885526162447122, 
    0.028215615646096551, 0.028521814759202128, 0.028802748773176134, 
    0.029057191278174393, 0.029284072314319318, 0.029482497466171934, 
    0.029651767542630596, 0.029791394021270113, 0.02990111259031223, 
    0.029980896459395459, 0.030030963900177211, 0.030051765029315697, 
    0.030043978881116099, 0.030008491137171675, 0.029946367649670631, 
    0.029858811808694388, 0.029747137281396729, 0.029612739916922218, 
    0.02945706689239689, 0.029281604332084661, 0.02908785497443412, 
    0.02887733937046344, 0.028651589684562183, 0.028412131980711432, 
    0.028160492660383816, 0.027898185834501005, 0.027626712659181926, 
    0.027347554421927326, 0.027062178208704959, 0.026772026170276617, 
    0.026478511731529125, 0.026183006027267974, 0.025886830539994871, 
    0.025591232942835742, 0.025297374122745887, 0.025006301574691678, 
    0.024718938679395105, 0.024436045012831576, 0.024158191260913175, 
    0.023885730166116739, 0.023618773581457714, 0.023357190014581822, 
    0.023100585474653684, 0.022848332578604746, 0.022599587422175715, 
    0.022353327459193169, 0.022108401476303989, 0.021863577600937427, 
    0.021617599327888488, 0.021369248831219479, 0.021117374526473696, 
    0.020860944108441984, 0.020599059041056748, 0.020330996961166685, 
    0.020056223203857734, 0.019774402151592735, 0.01948541481568292, 
    0.019189382945279179, 0.018886679299747463, 0.018577959395939394, 
    0.018264170548255403, 0.017946518858692445, 0.01762645805312606, 
    0.017305610686860269, 0.016985681122585566, 0.016668371185031689, 
    0.016355311685816696, 0.016048015279451339, 0.015747834290025881, 
    0.015455943490260944, 0.015173309447033698, 0.014900667311212286, 
    0.01463850092536801, 0.014387028987464277, 0.014146217614162593, 
    0.013915785736807976, 0.01369525491390914, 0.013483968423665111, 
    0.013281159821509861, 0.013085979930719948, 0.012897539999125095, 
    0.012714938958580833, 0.012537304756939762, 0.01236380075349997, 
    0.012193655582229875, 0.012026175525149983, 0.01186077100886225, 
    0.011696944077333732, 0.011534328665747183, 0.011372672903892173, 
    0.011211843184993842, 0.011051810566943944, 0.010892662633172305, 
    0.010734586568445401, 0.010577849392301547, 0.01042279920660368, 
    0.010269841271852228, 0.010119410754375112, 0.0099719695550803001, 
    0.0098280007657852077, 0.0096880045004823778, 0.0095525139742985102, 
    0.0094220831938040712, 0.0092972752063718109, 0.0091786367570722421, 
    0.0090666706615178116, 0.0089618223127760112, 0.0088644457097763231, 
    0.0087747880879007738, 0.0086929866568735276, 0.0086190301809996716, 
    0.0085527830046602492, 0.0084939510071434885, 0.0084420802353248354, 
    0.0083965260762384128, 0.0083564835485908755, 0.0083209448698039756, 
    0.0082887232267904645, 0.0082584414349180669, 0.0082285546546545883, 
    0.0081973594790344349, 0.0081630406558653289, 0.0081236947818118278, 
    0.0080773928414783844, 0.008022239232725931, 0.0079564366488424545, 
    0.007878335382086871, 0.0077865269223703713, 0.0076798906168892263, 
    0.0075576347087296294, 0.0074193357840727538, 0.0072649480529973446, 
    0.0070948025879529085, 0.0069095823618509928, 0.0067102683205108342, 
    0.0064980833639351763, 0.0062743963241765005, 0.006040628758589235, 
    0.0057981708715705493, 0.0055483173046788998, 0.0052922241058142106, 
    0.0050309304250678484, 0.0047653886001411613, 0.0044964801352813683, 
    0.0042251082977841263, 0.0039522165445443251, 0.003678858558862476, 
    0.0034062121315482246, 0.0031356064544594787, 0.0028684918876759296, 
    0.0026064920757718269, 0.0023512950238864677, 0.0021046847773168857, 
    0.00186845839399233, 0.0016444425131055156, 0.0014344487778681495, 
    0.0012402635066770321, 0.0010636198382923245, 0.00090622071304341599, 
    0.00076969363705283421, 0.00065558651095725209, 0.00056538229254711058, 
    0.00050047054549221979, 0.0004622054940764566, 0.00045186380484233329, 
    0.00047073159856634699, 0.00052007825073185747, 0.0006012397492844466, 
    0.0007155710781464519, 0.00086449988484582673, 0.0010494834925417519, 
    0.0012719462619158401, 0.0015332471695110243, 0.001834544179564057, 
    0.0021766731241105106, 0.0025600684340081306, 0.0029846543723669439, 
    0.0034497657483520288, 0.003954132811248655, 0.0044958343968979231, 
    0.005072375668926851, 0.0056807134223120937, 0.0063173400905246861, 
    0.0069784005397946075, 0.0076597719556979072, 0.008357180682163453, 
    0.0090663048994643232, 0.0097828954345860388, 0.010502876146260741, 
    0.011222470523036581, 0.01193830850378938, 0.012647525943137922, 
    0.013347861591335705, 0.014037736071737536, 0.014716357353807113, 
    0.015383699531342629, 0.0160405199983659, 0.016688317629702965, 
    0.017329124940255475, 0.017965277469864479, 0.01859913740533186, 
    0.019232781757271812, 0.0198675781809074, 0.020504102966165453, 
    0.021141912704515393, 0.021779631102934911, 0.022415104409918944, 
    0.02304557029013406, 0.02366791755326229, 0.024278973157615812, 
    0.024875809740365091, 0.025455880732214737, 0.026017197846047224, 
    0.026558363547371892, 0.027078298596970359, 0.027576061152959314, 
    0.028050498145143047, 0.028499858806463829, 0.028921730945277425, 
    0.029312612282468484, 0.029667943063915472, 0.029982623563449377, 
    0.030250932555997156, 0.030466979253933154, 0.030625324567682452, 
    0.030720586222547655, 0.030747947133626347, 0.03070309698135,
  // Fqt-total(2, 0-1999)
    0.99999999999999956, 0.99912099397931353, 0.99649405232743093, 
    0.99214881327123461, 0.98613352705625135, 0.97851370627121459, 
    0.96937035196335053, 0.95879785977696375, 0.94690170494398629, 
    0.93379601344866914, 0.91960111874456385, 0.9044411839762464, 
    0.88844196230957884, 0.87172874990310045, 0.85442456576052128, 
    0.83664857997492093, 0.81851479760361456, 0.8001310044455231, 
    0.7815979434638155, 0.76300872685504972, 0.74444845204903387, 
    0.72599400504485856, 0.70771403327933446, 0.68966905577013859, 
    0.67191170098469288, 0.65448703200351754, 0.63743294454006572, 
    0.62078062017012092, 0.60455500973179566, 0.58877533849307839, 
    0.5734556327326451, 0.55860523471564849, 0.54422932673538049, 
    0.5303294251479308, 0.51690385548859519, 0.50394819395006341, 
    0.49145567558273162, 0.47941756789929457, 0.46782350512539045, 
    0.45666179656235767, 0.44591969387471259, 0.4355836398954529, 
    0.42563948419803604, 0.41607268051030988, 0.40686845575036512, 
    0.39801195894291685, 0.38948838685887854, 0.38128309422329171, 
    0.37338168335194855, 0.36577008032079633, 0.35843458827966196, 
    0.35136194043890884, 0.34453933095204359, 0.337954445004919, 
    0.33159547182468435, 0.32545111967762053, 0.31951061908314105, 
    0.31376371953944659, 0.30820068633649922, 0.30281229428504941, 
    0.29758980687235043, 0.29252496197616967, 0.28760995357664221, 
    0.28283740037787619, 0.27820032581659926, 0.27369212757138367, 
    0.26930654947065186, 0.26503765928549611, 0.26087982170272772, 
    0.25682767852577659, 0.25287613033853618, 0.24902031480194964, 
    0.24525559418648621, 0.24157753575556515, 0.2379819004935573, 
    0.23446463160187697, 0.2310218465644695, 0.22764983075836873, 
    0.22434503118069959, 0.22110406084065251, 0.21792369138076273, 
    0.21480086036280324, 0.2117326700595524, 0.20871639331585728, 
    0.20574947991332185, 0.20282956607405042, 0.19995448016853479, 
    0.197122255069513, 0.19433113744521255, 0.19157958491371954, 
    0.18886627173594006, 0.18619008509931995, 0.18355011914207556, 
    0.18094567127477112, 0.17837623571168951, 0.17584150106665383, 
    0.17334133597547441, 0.17087578021477631, 0.16844502368681771, 
    0.1660493888385409, 0.16368930585151426, 0.16136528984576101, 
    0.15907791523195691, 0.15682779332297286, 0.15461555382243913, 
    0.15244182530683142, 0.15030721782921774, 0.14821231097811047, 
    0.14615764795002681, 0.1441437254336394, 0.14217099402655645, 
    0.14023985528988744, 0.13835066705934254, 0.13650374192613396, 
    0.13469935101831787, 0.13293772146607244, 0.13121902727746851, 
    0.129543380927954, 0.12791082750504959, 0.12632133587251562, 
    0.12477479639029301, 0.12327102119631819, 0.12180974456732029, 
    0.12039062744274992, 0.11901325727061111, 0.1176771483561424, 
    0.11638174045971558, 0.11512639505828488, 0.1139103912202872, 
    0.1127329188667657, 0.11159307478943678, 0.11048986376922496, 
    0.10942219855412774, 0.10838889969833175, 0.10738869381582855, 
    0.10642021492260763, 0.1054820047482793, 0.10457251643990109, 
    0.1036901248350165, 0.10283314002812251, 0.10199982420536789, 
    0.10118841086353095, 0.10039712495655857, 0.099624198327049371, 
    0.09886788871535844, 0.098126486950358166, 0.09739833455594353, 
    0.096681826286769704, 0.095975418519373787, 0.095277632533710355, 
    0.094587058626892456, 0.093902357875661507, 0.093222265916762997, 
    0.092545591325854853, 0.091871218480311906, 0.091198111426458908, 
    0.090525311949964993, 0.089851946828740259, 0.089177230819411729, 
    0.08850047598426404, 0.087821094913377612, 0.087138608330085923, 
    0.086452642531750001, 0.085762926741322992, 0.085069281392312568, 
    0.084371606451204562, 0.083669862727168864, 0.082964055248844301, 
    0.082254219360764685, 0.081540405947167813, 0.080822680811637501, 
    0.080101123379354724, 0.079375835029622088, 0.078646941801442147, 
    0.077914603560352916, 0.07717901686684106, 0.076440422942531686, 
    0.075699110281213164, 0.074955417018522652, 0.074209734813132394, 
    0.073462507587551656, 0.072714231441016478, 0.07196545214320868, 
    0.071216761459120689, 0.070468784932428433, 0.069722178589655223, 
    0.06897761264830915, 0.068235766396200298, 0.067497317488385722, 
    0.066762938436157993, 0.066033289916227728, 0.065309025439432372, 
    0.06459078898545921, 0.063879212702443122, 0.063174916825229688, 
    0.062478503998832501, 0.061790551382569947, 0.061111603593910692, 
    0.060442156397233542, 0.059782645718051391, 0.059133429344880632, 
    0.058494785566891819, 0.057866896147402987, 0.057249850734714482, 
    0.056643643159806689, 0.056048180036571117, 0.055463283554337071, 
    0.054888707149373932, 0.054324145596931828, 0.053769248631657079, 
    0.053223639829400787, 0.05268692884234881, 0.052158730523459942, 
    0.051638680425107282, 0.051126448876054026, 0.050621755588260139, 
    0.050124377985376972, 0.049634157563403516, 0.04915100032860005, 
    0.048674874706278196, 0.048205803336463106, 0.047743856289618143, 
    0.047289139586394857, 0.046841785558009261, 0.046401942509131294, 
    0.045969767373906789, 0.045545413399838856, 0.045129026803973349, 
    0.044720736985696757, 0.044320646979374219, 0.043928833088775876, 
    0.043545330628258806, 0.043170133245799866, 0.042803186278818926, 
    0.042444381498990498, 0.042093549538346438, 0.041750453001524732, 
    0.04141478562173017, 0.041086163651287678, 0.040764127103295425, 
    0.040448150363460333, 0.040137648622428537, 0.039832002128162965, 
    0.039530572490477298, 0.039232736908277527, 0.038937904552063814, 
    0.038645542333379558, 0.038355188627027283, 0.038066465476961769, 
    0.03777908582555424, 0.03749285347484449, 0.037207666984659674, 
    0.03692351506068401, 0.036640472446659883, 0.036358697601407898, 
    0.036078433167390643, 0.03579999713594896, 0.03552378619882151, 
    0.035250263105804334, 0.03497994581754596, 0.034713390125317857, 
    0.03445116727940515, 0.034193841866422957, 0.033941940383307653, 
    0.033695928217542852, 0.033456189663048523, 0.033223004993569692, 
    0.032996547874240605, 0.032776879056148803, 0.032563952495081212, 
    0.032357628650050672, 0.032157684012892304, 0.031963830470167778, 
    0.031775728242819115, 0.031593004650796196, 0.031415268701296913, 
    0.031242125163116103, 0.031073187672653206, 0.030908090081480148, 
    0.03074649804818097, 0.03058811639479983, 0.030432696428036074, 
    0.030280038317863744, 0.030129992202508858, 0.029982459210820933, 
    0.029837386029182261, 0.029694763141050642, 0.029554615603284883, 
    0.029416998421773748, 0.029281987031053055, 0.029149665155582597, 
    0.029020118248418419, 0.028893420780232451, 0.028769627014661573, 
    0.028648770352201189, 0.028530856045216709, 0.028415864400641047, 
    0.028303748259812404, 0.028194434333751437, 0.028087819876769615, 
    0.027983766135434018, 0.027882091759784046, 0.027782562573113512, 
    0.027684886796079604, 0.027588706115053839, 0.027493596624844432, 
    0.0273990650637537, 0.027304553136862322, 0.027209437565939305, 
    0.027113040315641181, 0.027014631414958998, 0.026913443169558494, 
    0.026808683174558288, 0.026699553853814291, 0.026585270548239046, 
    0.026465086908657301, 0.026338317955694399, 0.026204361439810697, 
    0.026062720784757423, 0.025913024371580915, 0.025755038349190087, 
    0.025588680986274634, 0.025414032895437685, 0.02523134046257303, 
    0.025041018265190368, 0.024843642764520762, 0.024639941434989127, 
    0.024430779719599931, 0.024217138278417413, 0.024000095800147191, 
    0.023780806287393957, 0.023560484634445225, 0.023340389754259554, 
    0.023121812613332404, 0.022906067705893932, 0.022694479447823192, 
    0.022488370103524221, 0.022289041690657683, 0.022097757395242144, 
    0.021915716407938757, 0.02174402957212913, 0.021583692025784126, 
    0.021435558442266963, 0.02130032147381589, 0.021178488819370348, 
    0.021070369358026423, 0.020976057681466192, 0.020895426599224016, 
    0.020828127450836769, 0.020773589054947566, 0.020731032318324873, 
    0.020699484681404281, 0.020677800357436018, 0.020664686143440258, 
    0.020658727963719849, 0.020658418778034499, 0.020662186437381099, 
    0.020668420036063864, 0.020675497425648115, 0.020681812764980965, 
    0.020685801236138644, 0.02068596181591854, 0.020680881305902021, 
    0.020669258034221826, 0.020649924252318968, 0.020621863538168663, 
    0.020584225927548779, 0.02053633581472324, 0.020477694240228307, 
    0.020407976471527988, 0.020327022779520192, 0.020234826798822915, 
    0.020131521243957302, 0.020017362863270848, 0.019892715063521853, 
    0.019758031609084112, 0.019613844472120869, 0.019460750801017418, 
    0.019299403692875666, 0.019130507557428844, 0.01895481285335569, 
    0.01877311672685647, 0.018586261196707463, 0.01839513227162333, 
    0.018200657983743221, 0.018003799533190128, 0.017805548206655641, 
    0.017606907866113103, 0.01740888825574163, 0.017212490612021247, 
    0.017018701037702755, 0.016828483623933198, 0.016642773375234558, 
    0.0164624680347722, 0.016288415863429762, 0.016121402235769227, 
    0.015962135953873465, 0.015811236494473236, 0.015669226850337791, 
    0.015536528277099587, 0.015413457844344568, 0.015300233619358651, 
    0.015196975320684054, 0.015103705907774713, 0.015020353257482681, 
    0.014946747104520715, 0.014882618499476339, 0.01482760282665012, 
    0.014781245041233779, 0.014743006493256864, 0.014712275960446665, 
    0.014688377366006901, 0.014670583254210482, 0.014658126582561225, 
    0.014650209731290482, 0.014646018125589135, 0.014644732319434134, 
    0.014645540866227033, 0.014647655355543793, 0.014650322067857867, 
    0.01465283661445177, 0.014654552846179501, 0.014654892557013296, 
    0.014653355353322021, 0.014649525398146427, 0.014643076056013962, 
    0.014633777296070792, 0.014621496859212985, 0.014606203465805774, 
    0.014587966885009565, 0.014566953778873492, 0.014543422439519499, 
    0.014517713933888583, 0.014490245061024818, 0.014461499993052898, 
    0.014432016864372905, 0.014402372807180867, 0.014373171652169909, 
    0.014345023609977092, 0.014318523640942538, 0.014294230446097452, 
    0.014272648806337785, 0.014254209711521965, 0.014239261903467089, 
    0.014228064030170915, 0.014220779375704876, 0.014217480271227902, 
    0.014218147531061855, 0.014222678151519142, 0.014230887258035776, 
    0.014242511026282097, 0.014257212945238429, 0.01427458219041932, 
    0.014294140028179846, 0.01431534822709442, 0.014337619076487979, 
    0.01436032817784544, 0.014382827502683576, 0.014404459909716297, 
    0.014424568562556968, 0.01444251233115545, 0.014457671709336052, 
    0.014469456238002771, 0.014477312286582564, 0.014480731002818785, 
    0.014479251225510407, 0.014472469313430648, 0.014460042644465813, 
    0.014441692464197612, 0.014417206050977788, 0.014386434804860687, 
    0.014349293050717814, 0.014305748308347114, 0.014255819518211912, 
    0.014199572533149057, 0.014137114530585268, 0.014068594150273901, 
    0.013994201614362246, 0.013914169756406402, 0.013828775787627697, 
    0.013738346320293814, 0.013643256364968558, 0.013543931766847204, 
    0.013440847283120488, 0.013334524046288911, 0.013225519949092128, 
    0.013114422032293708, 0.013001833514864171, 0.012888357745515361, 
    0.012774586212920876, 0.012661081836984407, 0.012548372392016106, 
    0.012436941466482474, 0.012327226639954126, 0.012219621072355016, 
    0.012114478298359793, 0.012012110226368337, 0.011912787004261646, 
    0.011816730460290678, 0.011724104374555415, 0.011635008195371995, 
    0.011549462917706149, 0.011467410589200854, 0.011388711298177574, 
    0.011313143436259611, 0.011240411629303906, 0.011170157366736416, 
    0.011101971161166143, 0.011035407812751929, 0.010970001734394311, 
    0.010905282549611239, 0.010840794012640896, 0.010776106041735666, 
    0.010710831744860958, 0.01064463931345948, 0.010577258840474241, 
    0.010508486039775019, 0.010438182208410448, 0.010366269766617815, 
    0.010292724855212165, 0.010217564777738802, 0.010140839544290549, 
    0.010062615015971246, 0.0099829602601046886, 0.0099019407487678027, 
    0.0098196093084352669, 0.0097360093622215205, 0.0096511780986576947, 
    0.0095651504536288408, 0.0094779715371801718, 0.0093896966415089513, 
    0.0093004017250719693, 0.0092101805924428362, 0.0091191522193614961, 
    0.0090274565703384966, 0.0089352540307668822, 0.0088427194682341118, 
    0.0087500437536918892, 0.0086574276214323176, 0.0085650819956736377, 
    0.008473226292358577, 0.0083820920236672269, 0.0082919184177351491, 
    0.0082029530918723351, 0.0081154479038794726, 0.0080296551576893912, 
    0.0079458203774283604, 0.007864171890512894, 0.0077849154748854538, 
    0.0077082212780497823, 0.0076342148203033229, 0.0075629635692307491, 
    0.0074944652492898315, 0.0074286402054444039, 0.0073653233843067956, 
    0.0073042621744249282, 0.0072451205993921287, 0.007187481936544767, 
    0.0071308638239869181, 0.0070747297837245662, 0.0070185094109915577, 
    0.0069616123108290776, 0.0069034455219326414, 0.0068434254035286959, 
    0.0067809898351745288, 0.006715612126947706, 0.0066468154703011127, 
    0.00657418467429854, 0.0064973864116291543, 0.0064161790780665976, 
    0.0063304273331660889, 0.0062401075646337503, 0.0061453159757608646, 
    0.006046267344221385, 0.0059432983726852313, 0.0058368567933912785, 
    0.0057274989840351209, 0.0056158752282619391, 0.0055027166154192151, 
    0.0053888184661203473, 0.0052750221131399339, 0.0051621938989429295, 
    0.0050512094325640558, 0.0049429310733513938, 0.0048381934181095741, 
    0.0047377850261016343, 0.0046424319335595801, 0.0045527806491332187, 
    0.0044693819427020602, 0.0043926774084939585, 0.0043229858123074137, 
    0.0042604986683611639, 0.0042052704537758959, 0.0041572238700144466, 
    0.0041161553921520893, 0.0040817474374440733, 0.0040535873221612404, 
    0.0040311857080481735, 0.0040139999699635529, 0.004001455929293205, 
    0.0039929690228204043, 0.0039879654920511806, 0.0039859022429795561, 
    0.003986277762080946, 0.0039886469307222972, 0.0039926240443117602, 
    0.0039978824240439522, 0.0040041486183622615, 0.0040111949187621801, 
    0.0040188273100572091, 0.0040268743306729341, 0.0040351833014500051, 
    0.0040436066289991721, 0.0040519984372220704, 0.0040602092251827669, 
    0.004068078647925636, 0.0040754311001657976, 0.0040820697211750969, 
    0.0040877686702577055, 0.0040922638684713023, 0.0040952466951904966, 
    0.004096356277769924, 0.0040951731847794492, 0.0040912175623717103, 
    0.0040839477276084016, 0.0040727635963379921, 0.0040570146258778151, 
    0.0040360115938669712, 0.004009034121236362, 0.0039753449848443333, 
    0.0039342056098064385, 0.0038848892605147655, 0.0038266994357535476, 
    0.003758989976007585, 0.0036811843708057538, 0.003592794417828545, 
    0.0034934376315563669, 0.0033828486297093866, 0.0032608861091023471, 
    0.003127540492120539, 0.0029829295652242763, 0.0028272977454445684, 
    0.0026610058261204057, 0.0024845262776490911, 0.002298431934044724, 
    0.002103387523202153, 0.0019001426761919081, 0.0016895177183523715, 
    0.0014723999159041684, 0.0012497283298996203, 0.0010224886228375376, 
    0.00079170232353942792, 0.00055841899251945961, 0.00032370772898756824, 
    8.8647209433146478e-05, -0.00014568444934069311, -0.00037822430395474519, 
    -0.00060794275848550063, -0.00083386605723516848, -0.0010550997191439331, 
    -0.0012708611188976162, -0.001480498148228546, -0.0016835096809523912, 
    -0.0018795450079968142, -0.0020684012704097316, -0.0022500104585514032, 
    -0.0024244208942084127, -0.0025917825889533769, -0.0027523298310303626, 
    -0.0029063683734309401, -0.0030542655240336281, -0.0031964376258395771, 
    -0.0033333461439164001, -0.0034654869154826587, -0.0035933865579460922, 
    -0.0037175926911200475, -0.0038386781696211113, -0.0039572307029241147, 
    -0.0040738516591048565, -0.0041891575958202159, -0.0043037745996122225, 
    -0.0044183376372298501, -0.0045334875136912858, -0.004649864473623453, 
    -0.004768097668888545, -0.0048887882086709926, -0.0050124874761565122, 
    -0.005139672527845039, -0.0052707225871887692, -0.0054059003047349664, 
    -0.0055453415993905308, -0.0056890452037404856, -0.0058368722021283201, 
    -0.0059885597819829628, -0.0061437369068340396, -0.0063019593980235423, 
    -0.0064627447656937665, -0.0066256124654879194, -0.0067901208135983876, 
    -0.0069558909926301345, -0.0071226306291391379, -0.0072901485275213406, 
    -0.0074583641609443545, -0.0076273121505218379, -0.0077971422155983716, 
    -0.0079681124347578767, -0.0081405777704476392, -0.0083149759621321141, 
    -0.0084918063500320478, -0.0086716119105713155, -0.0088549550132320624, 
    -0.0090423929649276723, -0.009234462445393379, -0.0094316527773485141, 
    -0.0096343959654584983, -0.0098430481721508839, -0.010057878677303745, 
    -0.010279059594028752, -0.010506655956415322, -0.010740617410033121, 
    -0.010980773770344909, -0.011226827285964604, -0.011478352223705957, 
    -0.011734792892423811, -0.011995470680405665, -0.01225958807557811, 
    -0.012526243297888028, -0.012794446959621678, -0.013063141337968213, 
    -0.01333122685983225, -0.013597585274301003, -0.013861107986091676, 
    -0.014120713814647952, -0.01437537292801732, -0.014624127926854717, 
    -0.014866107720568055, -0.015100544187546612, -0.015326786939320457, 
    -0.015544313456521585, -0.015752739423142707, -0.015951821214004215, 
    -0.016141460703862867, -0.016321701593372189, -0.016492726642258256, 
    -0.016654856578829105, -0.016808542552355532, -0.01695435735528503, 
    -0.017092979627016596, -0.017225174137320675, -0.017351766548766794, 
    -0.017473613178711968, -0.017591576414358909, -0.017706489702170907, 
    -0.017819131670655519, -0.01793019222762969, -0.018040249617942171, 
    -0.018149743187109959, -0.018258955629895809, -0.018368000405686806, 
    -0.01847681491991511, -0.018585162089900614, -0.018692638098812709, 
    -0.018798687949372492, -0.01890262836116623, -0.019003673229754939, 
    -0.019100962878588274, -0.01919359481902785, -0.019280649398940402, 
    -0.01936121525363825, -0.01943441365463525, -0.019499416344898057, 
    -0.019555457643618376, -0.019601844159603015, -0.019637958637260495, 
    -0.019663262710301499, -0.019677297931443006, -0.019679681453085591, 
    -0.019670107520687003, -0.019648345959375618, -0.01961424526882008, 
    -0.019567733617753675, -0.019508817270075272, -0.019437582215875427, 
    -0.019354187367029936, -0.019258863566552865, -0.019151901507845764, 
    -0.019033646247964938, -0.018904487067706581, -0.018764842986789643, 
    -0.018615158547711879, -0.018455891664042264, -0.018287509298600478, 
    -0.018110480294598934, -0.01792527259173397, -0.017732357668057013, 
    -0.017532208541378679, -0.017325310170880737, -0.017112167079394652, 
    -0.01689331266716956, -0.016669315294310962, -0.016440783781965951, 
    -0.016208371379846206, -0.015972770354589223, -0.015734708621075805, 
    -0.015494945204019018, -0.015254263247769248, -0.015013464545931674, 
    -0.014773362785858168, -0.014534773106891706, -0.014298502193623176, 
    -0.01406533828799055, -0.013836033691683588, -0.0136112936844328, 
    -0.013391762812367, -0.013178010299348154, -0.012970518270132297, 
    -0.012769672184436035, -0.012575751957313343, -0.012388924335721299, 
    -0.012209240901017241, -0.012036632002062788, -0.011870905203306598, 
    -0.011711746135090661, -0.011558717887222143, -0.011411271034579798, 
    -0.011268748620263957, -0.011130402297467406, -0.010995408183437898, 
    -0.010862883699620055, -0.010731913525103403, -0.010601566055744001, 
    -0.010470917123829361, -0.010339068117064665, -0.010205166801665945, 
    -0.010068426345263976, -0.0099281409063561119, -0.0097836998259326242, 
    -0.0096346046272303941, -0.0094804755649557735, -0.0093210610745593676, 
    -0.0091562390867026763, -0.0089860173126738788, -0.008810530367167382, 
    -0.0086300350335965868, -0.0084449012241952313, -0.0082555997440601214, 
    -0.0080626923183493293, -0.0078668161880472744, -0.00766866988797, 
    -0.0074689961415542539, -0.0072685743947737483, -0.0070682086841617432, 
    -0.0068687169992666074, -0.0066709301557561209, -0.0064756805394930433, 
    -0.0062837997677366933, -0.006096106727924832, -0.0059133963513794243, 
    -0.005736422882796543, -0.0055658818511319444, -0.0054023905831334183, 
    -0.0052464699211580094, -0.0050985313242596173, -0.0049588640188079503, 
    -0.0048276280161655425, -0.0047048531042411298, -0.0045904391841594195, 
    -0.0044841630439300647, -0.0043856835571013343, -0.004294553999880716, 
    -0.0042102318612994355, -0.0041320940867896096, -0.0040594540604156548, 
    -0.003991577653664171, -0.0039277030681481011, -0.0038670613206599406, 
    -0.0038088926780298813, -0.0037524599818466301, -0.0036970606806778676, 
    -0.0036420326399094274, -0.0035867596366928188, -0.0035306728947890921, 
    -0.0034732509371184087, -0.0034140185111587659, -0.003352544887720767, 
    -0.003288442123581523, -0.0032213605519376427, -0.0031509928807584514, 
    -0.003077067847950202, -0.0029993544801559207, -0.0029176560194271259, 
    -0.0028318145340218326, -0.0027417103324999812, -0.002647262086990025, 
    -0.0025484327815347369, -0.0024452307206508351, -0.0023377188187508691, 
    -0.0022260149765194639, -0.0021102966704683833, -0.0019907997623266824, 
    -0.001867813677031017, -0.0017416733445601888, -0.0016127493801813288, 
    -0.0014814320485865475, -0.0013481171628804828, -0.001213188778467666, 
    -0.0010770049908089654, -0.00093988697075992657, -0.00080211328195242692, 
    -0.00066392429794077197, -0.00052553542616174472, 
    -0.00038715234592618698, -0.0002489891904890221, -0.00011128479466297468, 
    2.5688863650640569e-05, 0.00016162259958896557, 0.00029616995481122888, 
    0.0004289502946524352, 0.00055955229943116427, 0.00068753849841462372, 
    0.00081245099487753164, 0.00093381924783714448, 0.0010511668626668575, 
    0.0011640215475662745, 0.0012719264291590183, 0.0013744464678343473, 
    0.0014711801896274462, 0.0015617684194394895, 0.0016458990357751256, 
    0.001723317140066126, 0.0017938266426813702, 0.0018572968709219169, 
    0.0019136656266953952, 0.0019629394955312895, 0.0020051955981251744, 
    0.0020405809622102205, 0.0020693079001171582, 0.0020916488501946211, 
    0.0021079360518855717, 0.002118555451971117, 0.002123945028908896, 
    0.0021245863910149287, 0.0021210017739057983, 0.002113745658388763, 
    0.0021033922101389825, 0.0020905255311917449, 0.0020757278613792733, 
    0.0020595679344373478, 0.0020425918814033629, 0.0020253153456516759, 
    0.0020082161402774413, 0.0019917281778457029, 0.0019762358793007028, 
    0.0019620692089544838, 0.0019495012812224305, 0.0019387413727489089, 
    0.001929930977470703, 0.001923134180332109, 0.0019183339635840894, 
    0.0019154257390269817, 0.0019142137926847641, 0.001914417562181021, 
    0.0019156718889254375, 0.0019175375878570289, 0.0019195095802782072, 
    0.0019210272800434876, 0.0019214867975761193, 0.0019202499153214163, 
    0.0019166581722910984, 0.001910045823990266, 0.0018997544025395133, 
    0.0018851476040709319, 0.0018656241722357562, 0.0018406407116148894, 
    0.0018097194188302051, 0.0017724627033060495, 0.0017285614928093701, 
    0.0016778010121639758, 0.0016200554566623514, 0.0015552848426355166, 
    0.0014835204310623847, 0.0014048525231810513, 0.0013194120045652172, 
    0.0012273531937135678, 0.0011288399761797505, 0.0010240310664842583, 
    0.00091307249375348657, 0.00079609115864266256, 0.0006731889521410236, 
    0.00054444678141984525, 0.00040992543367928238, 0.00026967800926092609, 
    0.0001237608438435163, -2.7753828422592644e-05, -0.00018476157049098407, 
    -0.00034710987450480561, -0.00051458674117192574, 
    -0.00068690672598768646, -0.00086370039007065808, -0.0010445046146026989, 
    -0.0012287548653713012, -0.0014157803220436261, -0.0016048018773655722, 
    -0.0017949394072981268, -0.0019852210626991884, -0.0021746021815107707, 
    -0.0023619894661168778, -0.0025462704910281567, -0.0027263424320363161, 
    -0.0029011447142280739, -0.0030696809354157808, -0.0032310393722446329, 
    -0.0033844056746276225, -0.0035290747050899058, -0.0036644573669843937, 
    -0.0037900879651960192, -0.0039056194875758286, -0.0040108256309859761, 
    -0.004105589701974729, -0.0041898885403016707, -0.00426378069248736, 
    -0.0043273858097576832, -0.0043808655910939675, -0.0044244058943984027, 
    -0.0044582035793117114, -0.0044824518398956644, -0.0044973330042609345, 
    -0.0045030135632426306, -0.0044996398683814073, -0.0044873434105150425, 
    -0.0044662421454574955, -0.0044364468110227977, -0.0043980699193764605, 
    -0.0043512335930002144, -0.0042960794480010438, -0.0042327799025057671, 
    -0.0041615413636867235, -0.0040826125792786765, -0.0039962860558234439, 
    -0.0039029006368864545, -0.0038028369382835945, -0.0036965144343045621, 
    -0.003584386220012223, -0.0034669323897752349, -0.003344653127358085, 
    -0.0032180589615339568, -0.0030876632039488015, -0.0029539724575730233, 
    -0.0028174795070097318, -0.0026786592003390196, -0.0025379660108239407, 
    -0.0023958354799289796, -0.0022526897445897184, -0.0021089468287591264, 
    -0.0019650308889526693, -0.0018213832192395831, -0.0016784747955872149, 
    -0.0015368128311156462, -0.0013969419034624432, -0.0012594470827748563, 
    -0.0011249487432907909, -0.0009940990058520025, -0.0008675792251144433, 
    -0.00074609531739326792, -0.00063037241041656697, 
    -0.00052115025209803446, -0.00041916958946364526, 
    -0.00032516191394806721, -0.0002398325603018134, -0.00016384482945671551, 
    -9.7797858588891795e-05, -4.2209405579760493e-05, 2.5036574100066477e-06, 
    3.6040136718573237e-05, 5.8220428104934283e-05, 6.8994145278842406e-05, 
    6.843067896269357e-05, 5.6714011484322946e-05, 3.4123561026762697e-05, 
    1.0155602445907435e-06, -4.2196148497731846e-05, -9.5060742306907634e-05, 
    -0.00015710569670990279, -0.00022784844707845504, 
    -0.00030679913107000447, -0.00039346049192793626, 
    -0.00048732202070972592, -0.00058785224706303868, 
    -0.00069449347655050687, -0.00080665799052890305, -0.0009237257766683965, 
    -0.0010450429642951571, -0.0011699211730291637, -0.0012976323493971561, 
    -0.0014274013504657508, -0.0015584044670893175, -0.0016897647981762973, 
    -0.0018205489519941749, -0.0019497699742400125, -0.0020763860388386167, 
    -0.0021993037409851544, -0.0023173838277192149, -0.0024294496817939804, 
    -0.0025342982361631298, -0.002630714934409552, -0.0027174975509448632, 
    -0.0027934721142080766, -0.0028575223740240035, -0.0029086101354671473, 
    -0.002945800534428303, -0.0029682845784232714, -0.0029753976514009027, 
    -0.0029666407251130642, -0.0029416944638312628, -0.0029004371840617832, 
    -0.002842953465741318, -0.0027695442055414221, -0.0026807297745185255, 
    -0.0025772478575236905, -0.002460046747104695, -0.0023302739003147142, 
    -0.002189257880400293, -0.002038485100362827, -0.0018795755953329577, 
    -0.0017142502159558327, -0.0015443035499276313, -0.0013715696424108888, 
    -0.0011978959389594081, -0.0010251157920501365, -0.00085502268425537457, 
    -0.00068934722530628197, -0.00052973770792891705, 
    -0.00037774200811130132, -0.00023478840076427738, 
    -0.00010217661914428435, 1.8928780474494355e-05, 0.00012750851429293604, 
    0.00022268602308204728, 0.0003037281736419724, 0.00037004162170565548, 
    0.00042116881632638114, 0.00045677955422692763, 0.00047666788517115253, 
    0.00048074347839040834, 0.00046902753269669975, 0.00044165074485083588, 
    0.00039884723123995332, 0.00034095156848285436, 0.00026839362351649897, 
    0.00018168875543088191, 8.1432691595028928e-05, -3.1711870377865215e-05, 
    -0.00015702359233797709, -0.00029373015292769164, 
    -0.00044101378168255525, -0.00059801674987421409, 
    -0.00076384344379285907, -0.00093756543322396128, -0.0011182232848675334, 
    -0.0013048303278778033, -0.0014963773149925513, -0.0016918455073377078, 
    -0.0018902151739085536, -0.0020904789644817694, -0.0022916606197935429, 
    -0.0024928274667795278, -0.0026931086545571906, -0.0028917110343239399, 
    -0.0030879292044115347, -0.0032811568029526058, -0.0034708965797853007, 
    -0.0036567589584750909, -0.0038384626104625993, -0.0040158281710501696, 
    -0.0041887723717987171, -0.0043572915426640466, -0.0045214521168724644, 
    -0.0046813805487501779, -0.0048372504211083153, -0.0049892774109299024, 
    -0.0051377128271769901, -0.0052828332773152608, -0.0054249317172741984, 
    -0.0055643063148526992, -0.0057012486887765643, -0.0058360266351461442, 
    -0.0059688726578072766, -0.0060999730843168546, -0.0062294594780748103, 
    -0.0063574020369867616, -0.0064838072933398258, -0.0066086197417695395, 
    -0.0067317205275683762, -0.0068529297107962394, -0.0069720006086005657, 
    -0.0070886214418350519, -0.0072024085697744633, -0.0073129115347707859, 
    -0.0074196101321375657, -0.0075219235288910211, -0.0076192200019409946, 
    -0.007710833733091697, -0.0077960834701791739, -0.007874292348274501, 
    -0.0079448105350181947, -0.008007028148127782, -0.0080603896104440142, 
    -0.0081044024243898463, -0.0081386411336740079, -0.0081627522806910074, 
    -0.0081764530668117039, -0.0081795329702799638, -0.0081718507138631123, 
    -0.0081533336323127148, -0.0081239754050430359, -0.0080838348115779505, 
    -0.0080330328453118195, -0.00797174840338764, -0.0079002144945400817, 
    -0.0078187071688343643, -0.00772753905373939, -0.0076270531903377551, 
    -0.0075176110072927042, -0.007399587667559368, -0.0072733683377930293, 
    -0.0071393397675636018, -0.006997894633237859, -0.0068494198384088049, 
    -0.006694302109584614, -0.0065329198461069023, -0.0063656476507294993, 
    -0.0061928510860798387, -0.0060148946409939548, -0.0058321437157119408, 
    -0.0056449709557063743, -0.0054537644221627039, -0.0052589321110434514, 
    -0.0050609099170804955, -0.0048601600056612576, -0.0046571720882164006, 
    -0.0044524593649858182, -0.0042465490110086745, -0.0040399727820330964, 
    -0.0038332547646355614, -0.0036269019925457965, -0.00342138872903311, 
    -0.003217147384122859, -0.0030145560850958599, -0.0028139320081797627, 
    -0.0026155263339874032, -0.0024195189076470932, -0.0022260294252257526, 
    -0.0020351230256636104, -0.0018468387057018021, -0.0016611964191365035, 
    -0.0014782246119624568, -0.001297971435680555, -0.0011204999458636368, 
    -0.00094588497457191679, -0.00077419565645075474, 
    -0.00060547239095241976, -0.00043970772671891325, 
    -0.00027683418161375718, -0.00011671727647226541, 4.0837972304151724e-05, 
    0.00019607857804977428, 0.00034928340675290928, 0.00050074286542568509, 
    0.00065073958032730423, 0.00079953330135843111, 0.0009473458534166319, 
    0.0010943525074486101, 0.0012406784413006632, 0.0013863948730632283, 
    0.0015315220928100019, 0.0016760297335966388, 0.0018198422936938083, 
    0.0019628359246062952, 0.0021048493807773691, 0.0022456812654167179, 
    0.0023850981145933487, 0.0025228354073004518, 0.0026586010556696278, 
    0.0027920778978282441, 0.0029229252880456731, 0.0030507845586103008, 
    0.0031752819931976572, 0.0032960372303342269, 0.0034126697537320725, 
    0.0035248051712776863, 0.0036320763104482679, 0.0037341290018683797, 
    0.0038306259544536418, 0.0039212471916366867, 0.0040056982652933188, 
    0.0040837147609180946, 0.004155065641909002, 0.0042195700557951755, 
    0.0042771019372481274, 0.0043275986000864642, 0.0043710684774624286, 
    0.0044075899990075069, 0.0044373146214910066, 0.0044604548528100725, 
    0.0044772774740241281, 0.0044880911983547402, 0.0044932329559413528, 
    0.0044930576165317223, 0.0044879311912164486, 0.0044782217142657942, 
    0.00446430255534394, 0.0044465526597016088, 0.0044253566297035394, 
    0.0044011130249733089, 0.0043742333210082538, 0.0043451392590103163, 
    0.0043142560284664469, 0.0042820012940887478, 0.00424876602158947, 
    0.0042149057551986212, 0.0041807263641675677, 0.0041464826408067566, 
    0.0041123753304840313, 0.0040785661887983559, 0.0040451862087354526, 
    0.004012349844196959, 0.0039801709210482037, 0.0039487762791905294, 
    0.003918316547204783, 0.0038889741473721903, 0.0038609620303719366, 
    0.0038345269021458702, 0.0038099407681798634, 0.0037874919787091324, 
    0.0037674856331036855, 0.0037502294487603669, 0.0037360247571710504, 
    0.0037251524120091306, 0.0037178590058389409, 0.0037143390449368161, 
    0.0037147190055935447, 0.0037190499640268218, 0.0037272944058686446, 
    0.0037393279463459727, 0.00375494355917189, 0.0037738511810445656, 
    0.0037956945333846126, 0.0038200446176099071, 0.0038464164876867986, 
    0.0038742639950870889, 0.0039029898309708121, 0.0039319454609440425, 
    0.0039604428660859016, 0.0039877582806480986, 0.0040131459271979253, 
    0.0040358501985102956, 0.004055122712198391, 0.0040702330663619753, 
    0.004080483369329437, 0.0040852152335846079, 0.0040838219176646331, 
    0.0040757490983588844, 0.0040605014866022153, 0.0040376381842317189, 
    0.0040067719959613977, 0.00396756478518591, 0.0039197195239074334, 
    0.0038629789387660731, 0.0037971198490605582, 0.0037219557812887783, 
    0.0036373427797761304, 0.0035431844202776751, 0.0034394471736546562, 
    0.0033261664119436187, 0.0032034557961851551, 0.003071512692798495, 
    0.002930616492746996, 0.0027811256479655399, 0.0026234624589734218, 
    0.0024581034922777608, 0.0022855543752910695, 0.0021063488142154954, 
    0.0019210360827941544, 0.0017301893998960412, 0.0015344123076196196, 
    0.0013343461861481964, 0.0011306816437266427, 0.00092415561351572809, 
    0.00071555207051048942, 0.00050569205313015129, 0.00029542035955438498, 
    8.559382731352184e-05, -0.00012293336827353706, -0.00032932566679984418, 
    -0.00053277262305728745, -0.00073250582293919698, 
    -0.00092780067506216426, -0.0011179829730188775, -0.001302436165518174, 
    -0.001480594898473541, -0.0016519480205799755, -0.0018160198686299998, 
    -0.001972369101703187, -0.0021205775507368834, -0.002260239206258995, 
    -0.0023909633509741684, -0.002512377132065393, -0.0026241398344195033, 
    -0.0027259609613360801, -0.0028176096737512627, -0.0028989310233596467, 
    -0.0029698467489355745, -0.0030303639658708342, -0.0030805678128784197, 
    -0.00312061603440424, -0.0031507361462297543, -0.0031712214274945412, 
    -0.0031824253349596243, -0.0031847693714925729, -0.0031787357406879739, 
    -0.0031648655208618018, -0.0031437557542179982, -0.0031160364355551922, 
    -0.0030823692669223451, -0.0030434202802970267, -0.0029998557672586733, 
    -0.0029523254596934383, -0.0029014677949731008, -0.0028478934641860097, 
    -0.0027921915854267681, -0.0027349240045124903, -0.0026766251000631919, 
    -0.002617789008661481, -0.002558867046312046, -0.0025002502033374782, 
    -0.0024422664638866307, -0.0023851615504441766, -0.0023290864263966404, 
    -0.0022740861476987185, -0.0022200881057517327, -0.0021668920043081308, 
    -0.0021141726978446827, -0.002061484051168504, -0.0020082784325859936, 
    -0.0019539416140096203, -0.0018978366727996571, -0.0018393508509953189, 
    -0.0017779448817770945, -0.0017131802497914084, -0.0016447389452902391, 
    -0.0015724287561045423, -0.0014961859886958103, -0.0014160692561372853, 
    -0.0013322543468502247, -0.0012450236295881408, -0.0011547543493907562, 
    -0.0010619040108255356, -0.00096699445435115261, -0.00087059283539779023, 
    -0.00077330149155578436, -0.00067574349992802229, 
    -0.00057855832471833562, -0.0004823981325794312, -0.00038792142534406558, 
    -0.00029578654688844146, -0.0002066416558092242, -0.00012110704870232312, 
    -3.9753667151645421e-05, 3.6912334571660878e-05, 0.0001084661605626068, 
    0.00017456974798761248, 0.00023496988253102582, 0.00028948453412737976, 
    0.00033798889963434885, 0.00038040605441906991, 0.00041669747426044558, 
    0.00044686694036923769, 0.00047097405949672209, 0.00048914417135188218, 
    0.00050158403547551024, 0.00050858550238314819, 0.00051051342194642884, 
    0.00050778937002477072, 0.00050086526021942118, 0.00049019363767509978, 
    0.00047620759268703864, 0.00045931411563920242, 0.00043987639281692657, 
    0.00041821685128852698, 0.00039461580234639458, 0.00036930774610563347, 
    0.00034248078003580102, 0.00031427178870970619, 0.00028476956640661815, 
    0.00025400860353435743, 0.00022197643808005693, 0.00018861781156893304, 
    0.00015383365025591926, 0.00011749543433286035, 7.9450905777221775e-05, 
    3.9527660711496395e-05, -2.4562180137546889e-06, -4.6685778079105104e-05, 
    -9.3349787327655942e-05, -0.00014262878797506283, 
    -0.00019469211994690692, -0.00024969266372850356, 
    -0.00030775674897370371, -0.00036898354234366735, 
    -0.00043345302502139721, -0.00050123189419482982, 
    -0.00057238283282192175, -0.00064698299116277582, 
    -0.00072512953167896011, -0.00080694914159520101, 
    -0.00089260094155284026, -0.00098226670068270162, -0.0010761452937273371, 
    -0.0011744394462885317, -0.0012773349243830237, -0.0013849775862201639, 
    -0.0014974548674133662, -0.0016147758603151199, -0.001736848203955803, 
    -0.00186347439033703, -0.0019943442814775877, -0.0021290393637255589, 
    -0.0022670440273637724, -0.0024077615687361198, -0.0025505398367277232, 
    -0.0026946878325747243, -0.0028395046062533536, -0.0029842971518042691, 
    -0.0031284009472615092, -0.0032712032640760821, -0.0034121572322367991, 
    -0.0035507980727201714, -0.003686754558654672, -0.003819748597478299, 
    -0.0039495895564950088, -0.0040761541524652932, -0.0041993605844429429, 
    -0.0043191307291727552, -0.0044353620395608754, -0.0045478910100204724, 
    -0.0046564777183096357, -0.00476078469570765, -0.0048603947410947044, 
    -0.004954823610746781, -0.0050435569784385388, -0.005126094525499475, 
    -0.0052019886020184831, -0.0052708739568695304, -0.0053324918559831628, 
    -0.005386698729462759, -0.005433472525080623, -0.0054729308379085307, 
    -0.0055053363250070772, -0.0055310976983338938, -0.005550771101909097, 
    -0.0055650457284653516, -0.00557471259958212, -0.0055806430102933874, 
    -0.0055837404846079365, -0.0055849016022637976, -0.0055849716570578719, 
    -0.0055847121546381898, -0.005584762666403743, -0.0055856236206277823, 
    -0.0055876381254051132, -0.0055909820121395771, -0.0055956588201904215, 
    -0.0056015171327606162, -0.0056082658009660976, -0.0056155053037614195, 
    -0.0056227614478005063, -0.0056295222409627329, -0.0056352566850588473, 
    -0.005639435871315897, -0.0056415409681416758, -0.0056410573842493863, 
    -0.0056374838401017334, -0.0056303341243174156, -0.0056191455835424304, 
    -0.0056034910190968495, -0.0055829937505591631, -0.0055573514459435263, 
    -0.0055263495545657274, -0.0054898936870143803, -0.0054480275440186941, 
    -0.0054009507400422313, -0.0053490216208663312, -0.0052927551829404628, 
    -0.0052327951934690847, -0.0051698881523485661, -0.0051048462083988682, 
    -0.0050385012575466723, -0.0049716716801032398, -0.0049051294021439165, 
    -0.0048395694281406307, -0.0047755957649791188, -0.0047137188577015604, 
    -0.0046543552584128785, -0.0045978377728676445, -0.0045444308703391154, 
    -0.0044943352351357081, -0.0044477060394498861, -0.0044046442872100328, 
    -0.0043652095351175519, -0.004329423332264078, -0.0042972867618988296, 
    -0.0042687951399536716, -0.0042439635347728943, -0.0042228504364994974, 
    -0.0042055771675884599, -0.0041923416084258614, -0.0041834206740651797, 
    -0.0041791681098313875, -0.0041800034978151969, -0.0041864026787119916, 
    -0.0041988731928743629, -0.0042179414216205703, -0.0042441207046795435, 
    -0.0042778891530857264, -0.0043196721148752847, -0.0043698024196904741, 
    -0.0044285112860156005, -0.0044959019540451303, -0.0045719382128471238, 
    -0.0046564428590511846, -0.0047491024941679642, -0.0048494673713729269, 
    -0.0049569770461072096, -0.0050709630305618156, -0.0051906802122452037, 
    -0.0053153137148713586, -0.0054439950187445138, -0.0055758202087294352, 
    -0.0057098628973414212, -0.0058451840237794192, -0.0059808499986549425, 
    -0.0061159436989149992, -0.0062495829148403676, -0.0063809383757161484, 
    -0.0065092454390810886, -0.0066338268714537449, -0.0067540949156884638, 
    -0.0068695478458416434, -0.006979762452573474, -0.0070843602479678195, 
    -0.0071829882525451102, -0.0072753000688645496, -0.007360940125800069, 
    -0.0074395442567579276, -0.0075107422749151956, -0.0075741784320781831, 
    -0.0076295198322520524, -0.0076764887717599905, -0.0077148780498525575, 
    -0.0077445828981421673, -0.0077655989989679434, -0.007778029816917313, 
    -0.0077820767462238151, -0.0077780217746025154, -0.0077662035829890808, 
    -0.007746998247988233, -0.0077208042404292533, -0.0076880294501200019, 
    -0.0076490999515861175, -0.0076044533288523626, -0.0075545660194421922, 
    -0.0074999622304758786, -0.0074412396677727118, -0.0073790728261073774, 
    -0.0073142216117296254, -0.0072475085071983733, -0.0071798066891356474, 
    -0.0071120124303877385, -0.0070450030016103865, -0.0069796168666496575, 
    -0.0069166070997579328, -0.0068566240073393257, -0.0068001800844231866, 
    -0.0067476403972244114, -0.0066992157762543218, -0.0066549656655340564, 
    -0.0066148069316448758, -0.0065785378787466906, -0.0065458533605195933, 
    -0.0065163734755072289, -0.0064896615398164371, -0.0064652489328912129, 
    -0.0064426627521155227, -0.006421462152558793, -0.0064012793697782256, 
    -0.006381856711709326, -0.0063630734276536524, -0.0063449557309378807, 
    -0.0063276467500365148, -0.0063113717038045429, -0.0062963806086388492, 
    -0.0062829002614985191, -0.0062710918697342103, -0.0062610104281376417, 
    -0.006252592794316808, -0.0062456457758365757, -0.0062398507063128657, 
    -0.0062347769746675767, -0.0062299019805712617, -0.0062246305419427737, 
    -0.0062183178779686458, -0.0062103037773494907, -0.0061999215087914627, 
    -0.0061865180016444851, -0.0061694604100857205, -0.0061481472774450605, 
    -0.0061220097593425874, -0.0060905215769363353, -0.0060532086311457815, 
    -0.0060096726362066054, -0.0059596108089445656, -0.0059028382699003439, 
    -0.005839303338437565, -0.0057690887803789051, -0.0056924113415476336, 
    -0.0056096080641093119, -0.0055211133723811227, -0.0054274435672868413, 
    -0.0053291734961899402, -0.0052269304398009165, -0.0051213970604733249, 
    -0.0050133098037506733, -0.0049034715096618721, -0.0047927584894112878, 
    -0.0046821193797281814, -0.0045725545626153011, -0.0044650878076456547, 
    -0.0043607275741864406, -0.0042604289021275256, -0.0041650510635349736, 
    -0.0040753228085913208, -0.0039918164458476986, -0.0039149382146204349, 
    -0.0038449242182842587, -0.0037818605357112602, -0.0037256940121931175, 
    -0.0036762658375587513, -0.0036333271097784342, -0.003596559453982115, 
    -0.0035655900954203587, -0.0035399857994207642, -0.0035192503537639455, 
    -0.0035028241375646986, -0.0034900718207806422, -0.0034802832783462369, 
    -0.0034726873404955882, -0.0034664460996750319, -0.003460668192832386, 
    -0.0034544137135939139, -0.003446694822234119, -0.0034364787319679049, 
    -0.0034227102681860253, -0.0034043184548840991, -0.0033802282675950289, 
    -0.0033493817546248281, -0.0033107410525857559, -0.0032632986584582775, 
    -0.0032060899639826156, -0.0031382115017502738, -0.0030588633683871352, 
    -0.0029673731538247738, -0.0028632480779994464, -0.0027462023166045526, 
    -0.0026161834261469652, -0.0024733921661638895, -0.0023182787919533102, 
    -0.0021515265982971336, -0.0019740386074518349, -0.00178688948101749, 
    -0.0015913044531008836, -0.0013886038696273671, -0.0011801590101909835, 
    -0.00096735310152934993, -0.00075153374732379462, 
    -0.00053399654510378244, -0.00031596495789124816, 
    -9.8592267189960553e-05, 0.00011702563550826905, 0.00032984316918919089, 
    0.00053883896635118726, 0.00074302689791922057, 0.00094144691869657213, 
    0.0011331785733697231, 0.0013173602897694234, 0.001493201775493771, 
    0.0016600008705708127, 0.0018171503805489942, 0.0019641622884492916, 
    0.0021006656073217804, 0.0022264143348256051, 0.0023413052397847777, 
    0.0024453500723951587, 0.0025386784048091618, 0.002621523104293119, 
    0.0026941791025306585, 0.0027569695745470468, 0.0028102067638573832, 
    0.0028541531656176536, 0.0028889785998076757, 0.0029147270979695541, 
    0.0029313004840315461, 0.0029384224169857311, 0.0029356465836755073, 
    0.0029223478889558612, 0.0028977411749302067, 0.0028609032262972029, 
    0.0028108146262474736, 0.0027464103572194111, 0.0026666293389617443, 
    0.0025704706420638392, 0.0024570611781946773, 0.0023256970793060056, 
    0.0021758734575498496, 0.0020073468269258738, 0.001820147823141179, 
    0.0016146331606187079, 0.0013915171017589657, 0.001151890147453485, 
    0.00089726305764357614, 0.00062957665032340447, 0.00035122077547204239, 
    6.5034862483573738e-05, -0.00022572320512856853, -0.00051748525947806819, 
    -0.0008064883490562564, -0.0010890125709743345, -0.001361578309343579, 
    -0.0016211175820376163, -0.0018650825859581064, -0.0020914808043635824, 
    -0.0022988498446575622, -0.002486212388416707, -0.0026530125899640036, 
    -0.0027990580665571488, -0.0029244492642165245, -0.0030295329361500934, 
    -0.0031148457314433956, -0.0031811090096982085, -0.0032291774392542195, 
    -0.0032600621944146066, -0.0032749017005988036, -0.0032749528490050046, 
    -0.0032615501471323872, -0.0032360691029938906, -0.0031998814311061255, 
    -0.0031543068238727491, -0.0031006164510304483, -0.0030400178098902936, 
    -0.0029736899325892236, -0.0029028232856334558, -0.0028286456234055952, 
    -0.0027524504668946384, -0.0026755970724323818, -0.0025994865997258443, 
    -0.0025255530936961904, -0.0024552162355821784, -0.002389877326729851, 
    -0.0023308794419889508, -0.0022794667349735499, -0.00223677519358274, 
    -0.002203785759289058, -0.0021813125608273628, -0.0021699691624794525, 
    -0.0021701659920335893, -0.0021821252167637823, -0.002205879821531964, 
    -0.0022413197143141563, -0.0022882272074249577, -0.0023463326115078435, 
    -0.0024153683232340348, -0.0024951161447894906, -0.0025854555267390837, 
    -0.002686357832590316, -0.002797856386438429, -0.0029200362568122108, 
    -0.003052948304655041, -0.0031966058551569894, -0.0033509261316540181, 
    -0.0035157460457713816, -0.0036907929700039253, -0.0038757012079890843, 
    -0.0040700429796309799, -0.0042733267141552593, -0.0044850424918146444, 
    -0.0047046604948382644, -0.0049316680072005424, -0.0051655686128915523, 
    -0.0054058965831086086, -0.0056522037251031778, -0.0059040236494848249, 
    -0.0061608202319815321, -0.0064219592996619711, -0.0066866367924155266, 
    -0.0069538285051150422, -0.0072222587403417164, -0.0074904002128834708, 
    -0.0077564948117512271, -0.0080185985344801702, -0.0082746439789812103, 
    -0.0085224882314131091, -0.008759933821711606, -0.0089847498902939985, 
    -0.009194663480748386, -0.0093873229814311586, -0.0095603084264740835, 
    -0.0097111373995451417, -0.0098372974565541834, -0.0099362980838789, 
    -0.010005744943399756, -0.010043410447896776, -0.010047334670078038, 
    -0.010015870146870026, -0.0099477578158651044, -0.009842207207173775, 
    -0.0096989220748527356, -0.0095182025402135682, -0.0093009691345691068, 
    -0.0090488385212220308, -0.0087641492182017992, -0.0084500010764535696, 
    -0.0081102770758707983, -0.0077495728845335997, -0.0073731853415049398, 
    -0.0069869783705991985, -0.0065972637869026888, -0.006210629640542178, 
    -0.0058337742626566515, -0.0054733940158547927, -0.0051359990164084922, 
    -0.0048277804592283613, -0.0045545047617789897, -0.004321376772171653, 
    -0.0041329340420059721, -0.003992983598519022, -0.0039044751326352909, 
    -0.0038695015403942628, -0.003889208089434036, -0.0039638172012008768, 
    -0.0040925957506474661, -0.0042739027524403067, -0.0045051681912251671, 
    -0.004782921819674402, -0.0051027841352744444, -0.0054595502380941682, 
    -0.0058472056324644969, -0.006258985299173239, -0.0066874896345896166, 
    -0.0071247570991937962, -0.0075625115376217762, -0.0079923080733199873, 
    -0.0084058348326171133, -0.0087950967890585898, -0.00915276283176388, 
    -0.0094723005623328586, -0.0097482709228610114, -0.0099763935831529548, 
    -0.010153724706199085, -0.010278768247257316, -0.010351480427525187, 
    -0.010373260156513128, -0.010346869573274855, -0.010276325046414295, 
    -0.010166781208946343, -0.010024203589391214, -0.0098551866679940092, 
    -0.009666584659982937, -0.0094651533043203888, -0.0092572819516039701, 
    -0.0090489245787799891, -0.0088455215634346863, -0.008652023467146483, 
    -0.0084729653905379464, -0.008312133629443906, -0.008172578949352206, 
    -0.0080561719320758635, -0.0079636970461046987, -0.0078946115732303011, 
    -0.0078472405208973098, -0.0078189747536673918, -0.0078063659586341495, 
    -0.0078055328635840346, -0.0078122614184040554, -0.0078228430439056772, 
    -0.0078337780594672918, -0.007842903389293325, -0.00784912989995999, 
    -0.0078531915497903563, -0.0078572172502032432, -0.0078660499872288975, 
    -0.0078858072068214158,
  // Fqt-total(3, 0-1999)
    0.99999999999999956, 0.99846471136867121, 0.99388228071062956, 
    0.98632198318067488, 0.97589643545085514, 0.96275773808925313, 
    0.94709243731803305, 0.92911562745031151, 0.90906451741142158, 
    0.88719179554963268, 0.86375909890267621, 0.83903083601554285, 
    0.81326856968153916, 0.78672610539847321, 0.7596453651214351, 
    0.73225308450442717, 0.70475832163725716, 0.67735074811606066, 
    0.65019962908098861, 0.62345344148796278, 0.59724001968879081, 
    0.57166714772281224, 0.54682350664363599, 0.52277987699723216, 
    0.49959053721017632, 0.47729475702796265, 0.45591835062583752, 
    0.43547523805130911, 0.41596897220462675, 0.39739420695839395, 
    0.3797380942104247, 0.36298157032716249, 0.34710054826546999, 
    0.33206698154784198, 0.31784981164390869, 0.30441579102813537, 
    0.29173019241680409, 0.27975741054899178, 0.26846146259479503, 
    0.25780641166497409, 0.24775670851630111, 0.2382774823783454, 
    0.22933477057842044, 0.22089571622359197, 0.21292871310634068, 
    0.20540352452186122, 0.19829136430488692, 0.19156495325052122, 
    0.18519854709494216, 0.17916794701110483, 0.17345047958969362, 
    0.16802497478512698, 0.1628717215478786, 0.15797242117843485, 
    0.15331012618460388, 0.1488691805575893, 0.14463515420566841, 
    0.14059477134996928, 0.136735842274432, 0.1330471992920291, 
    0.12951861900248127, 0.12614075384217235, 0.12290506375472317, 
    0.11980373253168346, 0.1168295868877068, 0.11397600380081811, 
    0.11123681124425085, 0.10860619790693213, 0.10607862027336556, 
    0.1036487326259531, 0.10131133633603057, 0.099061342792124765, 
    0.096893759629758769, 0.094803684115552428, 0.092786312148650449, 
    0.090836951005573874, 0.088951033159677909, 0.087124134680374304, 
    0.085351988125956013, 0.083630504674963413, 0.081955781206930839, 
    0.080324120913139008, 0.078732044126837097, 0.077176307617527182, 
    0.07565391931804534, 0.074162157715102053, 0.072698588095861605, 
    0.071261081582787184, 0.069847826423772671, 0.068457327391284614, 
    0.067088413513842093, 0.065740230134832697, 0.064412234438603569, 
    0.063104188757404922, 0.061816148588768369, 0.060548452995417695, 
    0.059301696559651812, 0.058076699523705998, 0.056874460656925516, 
    0.055696113095392616, 0.054542873004593817, 0.05341599177394276, 
    0.052316711497325807, 0.051246226407662111, 0.050205654338327563, 
    0.049196009189050635, 0.048218184556804655, 0.047272937772284064, 
    0.046360888252812725, 0.045482511698167846, 0.044638144198861321, 
    0.043827987302746133, 0.043052116856717941, 0.042310485944003336, 
    0.041602933633186595, 0.040929187187494158, 0.040288859678734544, 
    0.039681447949271163, 0.039106332981364671, 0.038562785098849438, 
    0.038049965897003567, 0.037566940822465332, 0.037112684010157486, 
    0.036686093900896617, 0.036285995294101835, 0.035911145128052283, 
    0.035560233192581031, 0.035231877458673816, 0.034924622789838058, 
    0.034636935066129852, 0.034367199424613193, 0.03411373145458968, 
    0.033874779780582377, 0.033648536083474401, 0.033433144696301799, 
    0.033226717837570793, 0.033027347741206345, 0.032833129835697895, 
    0.03264218802582524, 0.032452706192231499, 0.032262960338337962, 
    0.032071353775461081, 0.031876445281988623, 0.031676973376976655, 
    0.031471872332775756, 0.031260274711793025, 0.03104151593586273, 
    0.030815121783469339, 0.030580797171688712, 0.030338411043198718, 
    0.030087980483253594, 0.029829647128341061, 0.029563665772020381, 
    0.02929037783753391, 0.02901019605549273, 0.028723586188478905, 
    0.028431046074084042, 0.028133095163653438, 0.027830263533501765, 
    0.027523094685116146, 0.02721214701619417, 0.026898011204384262, 
    0.02658131950548227, 0.026262758520128947, 0.025943071065776466, 
    0.02562305574335114, 0.025303548387685889, 0.024985397571874974, 
    0.024669439064886476, 0.024356461248850405, 0.024047182830245772, 
    0.02374223528073453, 0.023442152809706053, 0.02314736038303962, 
    0.022858170313044518, 0.022574778608509562, 0.022297265779634971, 
    0.02202559737542974, 0.021759625426920868, 0.021499094852441589, 
    0.021243645828939336, 0.020992826506305202, 0.020746100170089234, 
    0.020502874023312228, 0.020262514205487039, 0.020024383059142302, 
    0.019787866943691921, 0.019552409432734775, 0.019317546100813716, 
    0.01908293725954777, 0.018848396740351429, 0.018613921271524274, 
    0.018379707135918029, 0.018146155193751949, 0.017913864231214983, 
    0.017683607380441339, 0.017456300328722942, 0.017232963085139542, 
    0.017014670007747264, 0.016802505104283997, 0.016597512074615343, 
    0.016400654797374389, 0.016212772538617692, 0.016034550684001815, 
    0.015866493488501922, 0.015708907127156998, 0.015561889569531168, 
    0.015425329765918476, 0.015298913134056355, 0.015182133172408829, 
    0.01507430810595198, 0.014974601676807826, 0.014882050303974331, 
    0.014795588966167563, 0.014714078594931047, 0.014636337867493219, 
    0.014561169156323849, 0.014487386866463352, 0.014413836297063899, 
    0.014339415131816158, 0.014263084980529993, 0.01418388702676949, 
    0.014100949640075891, 0.014013499758767797, 0.013920871304586828, 
    0.013822515675117632, 0.013718005297135212, 0.01360704560658987, 
    0.013489473682137916, 0.013365258474994949, 0.013234506402745727, 
    0.013097449142523193, 0.01295444031651229, 0.012805946343431846, 
    0.012652532595725284, 0.012494849628602651, 0.012333613040673224, 
    0.01216958870641548, 0.012003569199016264, 0.011836355937855109, 
    0.011668740322580405, 0.01150148663880857, 0.011335317679909217, 
    0.011170905324830853, 0.011008867007808013, 0.010849759740877825, 
    0.010694080946970205, 0.010542266451040739, 0.010394690763272237, 
    0.010251670220596967, 0.010113460506895749, 0.0099802665782005653, 
    0.0098522494739180233, 0.0097295306107907948, 0.0096122098911357867, 
    0.0095003784465771887, 0.009394133737821336, 0.0092936053450024762, 
    0.0091989704902652059, 0.009110467043098083, 0.0090284052286568415, 
    0.0089531674866865103, 0.0088852027308601797, 0.0088250079672444314, 
    0.0087731044246419244, 0.0087300153038504698, 0.0086962330688563523, 
    0.008672202256468562, 0.0086582926876445972, 0.0086547909269173717, 
    0.0086618904869649616, 0.0086796864381326402, 0.008708179763461988, 
    0.0087472777220496852, 0.0087968089295718584, 0.0088565334072790557, 
    0.0089261589569958697, 0.0090053585099810832, 0.0090937845266525867, 
    0.0091910828926995234, 0.009296903167258468, 0.0094109002595177283, 
    0.0095327347208127595, 0.0096620671515618654, 0.0097985523843153784, 
    0.0099418289857134447, 0.010091505786484264, 0.010247148935134284, 
    0.010408263937857917, 0.010574283948159067, 0.010744542531418924, 
    0.010918266067281881, 0.011094549309519102, 0.011272352982592172, 
    0.011450499522555261, 0.011627676915955615, 0.011802450814672256, 
    0.011973282011387264, 0.012138545944763927, 0.012296555674000783, 
    0.012445581950080465, 0.012583871666988152, 0.012709665237776863, 
    0.012821217912122309, 0.01291681358009527, 0.012994784420576099, 
    0.013053524816465519, 0.013091507850844215, 0.013107293631322398, 
    0.01309954393859797, 0.013067026726919109, 0.013008626984982527, 
    0.012923359445982172, 0.012810388910099287, 0.012669053660128509, 
    0.012498902956482533, 0.012299734426789161, 0.012071630097855545, 
    0.011814989171256193, 0.011530553668918697, 0.011219411607876775, 
    0.010882996196330529, 0.010523064018159039, 0.010141663524391496, 
    0.0097410901279126674, 0.0093238345235630033, 0.0088925296573898003, 
    0.0084498992551745762, 0.0079987062137321201, 0.0075417132188859747, 
    0.0070816480216326838, 0.0066211832694480482, 0.0061629223302575647, 
    0.0057093932849970235, 0.0052630490733847832, 0.0048262678048786182, 
    0.0044013459058670889, 0.0039904843175977908, 0.0035957771328612564, 
    0.0032191830917732223, 0.0028625022132838396, 0.0025273512592190891, 
    0.0022151428617254885, 0.0019270739577930164, 0.0016641097971757267, 
    0.0014269780473637743, 0.001216158841358549, 0.001031873960950459, 
    0.00087408059599229225, 0.00074246121356316317, 0.00063642333310559042, 
    0.00055509870973600333, 0.00049736259946018364, 0.00046185593041699378, 
    0.00044702772674860402, 0.00045117933666797736, 0.00047252014445419278, 
    0.00050921858023447221, 0.00055945010974861684, 0.00062143625479697145, 
    0.00069347672999880614, 0.00077397006915054967, 0.00086142988286290326, 
    0.00095448956698815477, 0.0010519095139032671, 0.0011525747117504983, 
    0.0012554976640155729, 0.0013598202822351776, 0.0014648168156448816, 
    0.0015698988516884731, 0.0016746174584812957, 0.0017786673928847604, 
    0.0018818832615564358, 0.0019842397516749693, 0.0020858419332923164, 
    0.0021869115932002304, 0.002287776871372126, 0.0023888538933339045, 
    0.0024906305597489622, 0.0025936543984064293, 0.002698517271094564, 
    0.0028058388348080345, 0.0029162542107228086, 0.0030303865482418802, 
    0.0031488327719398261, 0.0032721373530722651, 0.0034007718086114915, 
    0.0035351139765957603, 0.0036754314832697617, 0.0038218680498895846, 
    0.0039744372657786889, 0.0041330178178059238, 0.0042973501533598449, 
    0.0044670419985794151, 0.0046415681444436216, 0.0048202772652734972, 
    0.0050024013494744408, 0.0051870641791556564, 0.0053733007829200388, 
    0.0055600653342760169, 0.0057462488280990908, 0.0059306958055601253, 
    0.0061122162459593468, 0.006289597022899363, 0.0064616123902726209, 
    0.0066270327037391908, 0.0067846291551377164, 0.0069331800910943748, 
    0.0070714809473810388, 0.0071983542119208746, 0.0073126598807074844, 
    0.007413314620513145, 0.0074993118654917926, 0.007569748039871713, 
    0.0076238475934317018, 0.0076609865063816578, 0.0076807056685373933, 
    0.0076827248878735509, 0.0076669386022057209, 0.0076334114113128099, 
    0.0075823698183585383, 0.007514193468902192, 0.007429414102209965, 
    0.0073287139734180126, 0.0072129299432219752, 0.0070830600141567994, 
    0.0069402699893341899, 0.006785899057052909, 0.006621456666645366, 
    0.006448616251684006, 0.006269201933442459, 0.0060851658771697683, 
    0.0058985663571595928, 0.0057115405446570558, 0.0055262716978489263, 
    0.0053449490464590604, 0.0051697264997505711, 0.0050026750900390646, 
    0.0048457383282339648, 0.0047006871539596864, 0.0045690849745753303, 
    0.0044522619701064352, 0.0043512944475329988, 0.0042669954347343648, 
    0.0041999172208827462, 0.0041503511009093859, 0.0041183422324161259, 
    0.0041037008598999595, 0.0041060184676747838, 0.0041246821976086145, 
    0.0041588928259679277, 0.004207679034110165, 0.0042699106804242343, 
    0.00434431472320363, 0.0044294985972955095, 0.0045239783004993577, 
    0.0046262128718239379, 0.0047346443757256447, 0.004847738625325203, 
    0.0049640142257196028, 0.0050820759424608586, 0.0052006328934758057, 
    0.0053185089847464723, 0.0054346511214126052, 0.005548129115853207, 
    0.0056581372055166373, 0.0057639918788929207, 0.0058651282687230827, 
    0.0059610966706896322, 0.0060515544114383294, 0.006136259797508945, 
    0.0062150633785825393, 0.006287899623249233, 0.0063547778253691288, 
    0.0064157778363140199, 0.006471051347774974, 0.0065208143721403045, 
    0.0065653537449030155, 0.0066050221320138576, 0.0066402349539179395, 
    0.0066714634719351575, 0.006699229738356809, 0.0067240892701084919, 
    0.006746617511372126, 0.0067673901841371082, 0.0067869592806146803, 
    0.0068058212840923799, 0.0068243895996686092, 0.0068429616383282738, 
    0.0068616894803774572, 0.006880559523913571, 0.0068993788273135331, 
    0.0069177744399889886, 0.0069352113253622208, 0.0069510145459039229, 
    0.0069644048301603628, 0.0069745284445929465, 0.0069804902444173325, 
    0.0069813792083140364, 0.006976288980824012, 0.0069643328004361394, 
    0.0069446590740898581, 0.0069164652844137166, 0.0068790220093613557, 
    0.0068316911250784259, 0.0067739593866366641, 0.0067054642920621058, 
    0.0066260205556435423, 0.0065356394656076889, 0.0064345437428218986, 
    0.0063231774676107298, 0.0062022127963694551, 0.0060725512032233182, 
    0.0059353195432902319, 0.0057918640405916844, 0.0056437314036168829, 
    0.0054926464653177664, 0.005340476898564068, 0.0051892001609587651, 
    0.0050408591649677191, 0.0048975181378765912, 0.0047612219466459027, 
    0.0046339491718667214, 0.0045175704057761274, 0.0044138086285387991, 
    0.004324205204706901, 0.0042500917873299566, 0.0041925734706042212, 
    0.0041525102646028655, 0.0041305127043785627, 0.0041269322794571647, 
    0.0041418543258980676, 0.0041750944050639848, 0.0042261963866920922, 
    0.0042944339166349809, 0.0043788142730223131, 0.0044780855272371564, 
    0.0045907495981618333, 0.0047150792993543534, 0.0048491497673965062, 
    0.0049908781026428966, 0.0051380801699293698, 0.0052885290877263966, 
    0.0054400254527426093, 0.0055904634502781216, 0.005737892244255095, 
    0.0058805656346621682, 0.0060169797672137929, 0.0061458988247455968, 
    0.0062663655085063857, 0.0063777052598185842, 0.0064795156907828753, 
    0.0065716529813641565, 0.0066542153311602101, 0.0067275178698761639, 
    0.0067920659389047533, 0.0068485255321783121, 0.0068976879724733271, 
    0.0069404322602815661, 0.0069776881999248424, 0.0070104011094010406, 
    0.0070394977833436994, 0.0070658613601724454, 0.0070903058565588281, 
    0.0071135566001686362, 0.0071362385324294005, 0.0071588700374049319, 
    0.0071818605707353825, 0.0072055209995889888, 0.0072300635681112344, 
    0.0072556141451275346, 0.0072822215429589826, 0.0073098712767089595, 
    0.007338498373651337, 0.0073680031523510898, 0.0073982648592465106, 
    0.0074291607849465442, 0.0074605768412393083, 0.0074924209903021342, 
    0.0075246286190495254, 0.0075571764986755831, 0.0075900813996574636, 
    0.0076233994892315384, 0.0076572176803826851, 0.0076916459738299199, 
    0.0077267967780872164, 0.007762764198762327, 0.0077995950020566919, 
    0.007837269619525019, 0.0078756813100876021, 0.0079146141128523719, 
    0.0079537450470291496, 0.007992636464315056, 0.0080307489522308123, 
    0.0080674560523369739, 0.0081020716250569912, 0.0081338761749218686, 
    0.0081621479636303645, 0.0081861891132931335, 0.0082053432343390555, 
    0.0082190079657316045, 0.0082266384249998614, 0.0082277480388170121, 
    0.0082219011492365487, 0.0082087063313786585, 0.0081878100173157758, 
    0.0081588899403825573, 0.0081216537478976513, 0.0080758403110265994, 
    0.0080212261875706042, 0.0079576375358166775, 0.00788496314458461, 
    0.0078031708516335613, 0.0077123259384448547, 0.0076126024820579244, 
    0.0075042983500816811, 0.0073878374826570415, 0.0072637683804858445, 
    0.007132757608785568, 0.006995568673599138, 0.0068530429559239669, 
    0.0067060750078384015, 0.0065555854424342993, 0.0064024963448486433, 
    0.0062477067867866961, 0.0060920729916775626, 0.0059363906007368203, 
    0.0057813846866751843, 0.0056276969974530253, 0.0054758883709369148, 
    0.0053264407089604372, 0.0051797621205227455, 0.0050362012681031722, 
    0.0048960590695582267, 0.0047596076973317651, 0.0046271078267146552, 
    0.0044988267159128056, 0.0043750544644080369, 0.004256110746696626, 
    0.0041423488453378871, 0.0040341462214639624, 0.0039318949788877287, 
    0.003835975289861317, 0.0037467379716392508, 0.0036644822121371739, 
    0.0035894429318666971, 0.0035217865329548277, 0.0034616088247080494, 
    0.0034089447117184989, 0.0033637745021446127, 0.0033260339985258904, 
    0.0032956209637042696, 0.0032724052015790442, 0.0032562286540876676, 
    0.0032469116350820216, 0.0032442514269105877, 0.003248017133427485, 
    0.0032579459082919169, 0.0032737336258687657, 0.0032950184714112402, 
    0.0033213656327708077, 0.0033522545143688976, 0.0033870724782462543, 
    0.0034251216701142733, 0.0034656392170378178, 0.003507826267715185, 
    0.0035508904580980436, 0.0035940839805579487, 0.0036367412040168596, 
    0.0036783095209671065, 0.0037183622553933686, 0.0037566062693921865, 
    0.0037928663057391955, 0.0038270757472110965, 0.0038592462962860207, 
    0.0038894467021565286, 0.0039177743030061746, 0.0039443342944638403, 
    0.0039692156745422978, 0.0039924728253627091, 0.004014106754147046, 
    0.0040340572871373614, 0.0040521924147297024, 0.0040683214735365179, 
    0.0040822029821131062, 0.0040935661563891619, 0.0041021367234438553, 
    0.0041076606911478377, 0.0041099218892206146, 0.0041087548791350409, 
    0.0041040435178594185, 0.0040957220030008691, 0.0040837639075198126, 
    0.0040681682215293249, 0.0040489486002608108, 0.0040261154934153583, 
    0.003999660738677864, 0.0039695331059089517, 0.0039356098495775642, 
    0.0038976814285964041, 0.0038554267944439476, 0.0038084087728713291, 
    0.0037560817955867723, 0.0036978035495926673, 0.0036328648216733821, 
    0.0035605159869199093, 0.0034800050069434376, 0.0033906096481845331, 
    0.0032916712587683621, 0.0031826197630073602, 0.0030630005934878649, 
    0.002932491627225837, 0.0027909115948227051, 0.0026382334895831867, 
    0.0024745764291215981, 0.0023002079004064324, 0.002115528079607471, 
    0.0019210597523635275, 0.0017174311659497756, 0.0015053588459975399, 
    0.0012856294566997864, 0.0010590833761694057, 0.00082659977342198121, 
    0.00058908488717597507, 0.00034746736708435603, 0.00010269826889464181, 
    -0.00014424537913421937, -0.00039234955167458677, 
    -0.00064055434057486843, -0.00088774382277982645, -0.0011327430247031554, 
    -0.0013743166590671539, -0.0016111740963740257, -0.0018419859895054071, 
    -0.0020654013042154936, -0.0022800684346470329, -0.0024846554949353328, 
    -0.0026778718771853262, -0.0028584880755187364, -0.0030253537674447381, 
    -0.0031774182387287694, -0.0033137559580187336, -0.0034335925663912647, 
    -0.0035363311395629872, -0.0036215842684363692, -0.003689193795184691, 
    -0.0037392474506273672, -0.0037720783654301843, -0.0037882562683447655, 
    -0.0037885573955426903, -0.0037739376029143831, -0.0037454933158791114, 
    -0.00370442582247942, -0.0036520120824829107, -0.0035895720775206241, 
    -0.0035184552936824011, -0.0034400149649242498, -0.0033555967562604702, 
    -0.003266525630057417, -0.0031740904569231522, -0.0030795357588082406, 
    -0.0029840495153820169, -0.002888760674360653, -0.0027947297505094963, 
    -0.0027029510927569981, -0.0026143436295030234, -0.0025297533090648098, 
    -0.0024499461043109676, -0.0023756064630687667, -0.0023073336365247365, 
    -0.0022456409799768476, -0.0021909492262254067, -0.002143587951619251, 
    -0.0021037975037151114, -0.0020717298370118362, -0.0020474606493243461, 
    -0.0020309944774935724, -0.0020222790819432969, -0.0020212107579266037, 
    -0.0020276455190114838, -0.0020414041643634921, -0.0020622800528483612, 
    -0.0020900361372535249, -0.0021244079649353114, -0.0021651028082503468, 
    -0.0022117963159701726, -0.0022641327909092108, -0.0023217220051105231, 
    -0.0023841358521863283, -0.0024509145802502027, -0.0025215594339112308, 
    -0.0025955389093473362, -0.0026722850436508307, -0.0027512021182941539, 
    -0.0028316643489808809, -0.0029130296291770283, -0.0029946434675376167, 
    -0.0030758514466781117, -0.0031560076039285588, -0.0032344840733673883, 
    -0.0033106786945646173, -0.0033840250679654051, -0.0034540015973096808, 
    -0.0035201460990975982, -0.0035820643776281243, -0.0036394457969172148, 
    -0.0036920714303308962, -0.0037398200023042879, -0.0037826727953523534, 
    -0.0038207105881541731, -0.0038541068260607462, -0.0038831175146415951, 
    -0.0039080729370916346, -0.00392936682828216, -0.0039474474187304867, 
    -0.0039628099518874546, -0.0039759873734451267, -0.0039875408843256729, 
    -0.0039980462656503176, -0.0040080863042271792, -0.0040182261204060902, 
    -0.0040289996053314465, -0.004040890076823519, -0.0040543057689635424, 
    -0.0040695599983214641, -0.0040868516963245101, -0.0041062494385104885, 
    -0.0041276835630986138, -0.004150941359162592, -0.004175666596780152, 
    -0.004201371556849666, -0.0042274406793330792, -0.0042531483986576616, 
    -0.0042776702458733997, -0.0043000989668153973, -0.0043194571423378555, 
    -0.0043347159897621987, -0.0043448132646107356, -0.0043486783231536427, 
    -0.0043452594787873828, -0.0043335555150927083, -0.0043126502038496406, 
    -0.0042817488268178279, -0.004240210268574701, -0.0041875821908351363, 
    -0.0041236205494745706, -0.0040483115948199448, -0.0039618839277990358, 
    -0.0038648071792194314, -0.0037577873950676534, -0.0036417527031406324, 
    -0.0035178324434458836, -0.0033873329219514412, -0.0032517054870710724, 
    -0.003112511111073718, -0.0029713939804556417, -0.002830038313433654, 
    -0.0026901321927978957, -0.0025533279805270283, -0.0024211931943875472, 
    -0.0022951698077421207, -0.0021765259810915326, -0.0020663147470763215, 
    -0.0019653374140746025, -0.0018741120061231736, -0.0017928544578623604, 
    -0.0017214779505824768, -0.0016595947017948275, -0.0016065405972877428, 
    -0.0015614053266386797, -0.0015230755007465571, -0.0014902872657407257, 
    -0.0014616756145056713, -0.0014358240374294248, -0.0014113117567864555, 
    -0.0013867508462096906, -0.0013608134467323642, -0.0013322519746758056, 
    -0.0012999095592293515, -0.001262724058971428, -0.0012197280173628765, 
    -0.0011700428025665014, -0.0011128736663537347, -0.0010475042788738709, 
    -0.00097329210628933189, -0.00088967058730368047, 
    -0.00079614877054649173, -0.00069231674950793239, 
    -0.00057785594256552612, -0.00045254566002755458, 
    -0.00031627104246755684, -0.00016903400662525829, 
    -1.0958702804288822e-05, 0.00015770290157687499, 0.0003365678873178002, 
    0.00052512366045182589, 0.00072272887899632891, 0.00092862215092107733, 
    0.0011419229716444184, 0.0013616461292857368, 0.0015867065765512642, 
    0.0018159283806437547, 0.0020480520833280409, 0.0022817435341752914, 
    0.0025156026827111793, 0.0027481837434343683, 0.0029780123046231656, 
    0.0032036125206911675, 0.0034235345388449303, 0.0036363775460505204, 
    0.0038408127326552493, 0.004035595928610405, 0.004219574701251649, 
    0.0043916911839687323, 0.0045509840980366536, 0.0046965808989456251, 
    0.0048276925213300926, 0.0049435990695292312, 0.0050436355743796214, 
    0.0051271828772369186, 0.0051936568999224296, 0.0052425054043773109, 
    0.0052732097511113477, 0.005285293679764839, 0.0052783311369826802, 
    0.0052519550792017016, 0.0052058678063345749, 0.0051398439504739026, 
    0.0050537313983049321, 0.0049474478309962091, 0.0048209826909337405, 
    0.0046743963435475653, 0.0045078295223207124, 0.0043215087876773391, 
    0.0041157658164269247, 0.0038910480810400785, 0.0036479418463670997, 
    0.0033871830558361957, 0.003109671941906784, 0.0028164775888556313, 
    0.0025088460927445645, 0.0021881952527977471, 0.0018561101937728177, 
    0.0015143350264417601, 0.0011647638129714567, 0.00080942354521561775, 
    0.00045045902452504313, 9.010467491057166e-05, -0.00026934530918064023, 
    -0.00062557262268302647, -0.00097627969240734341, -0.001319226633064883, 
    -0.001652270921141026, -0.0019733986456662118, -0.0022807611054258005, 
    -0.0025726870632536924, -0.0028477028237205567, -0.0031045349082024104, 
    -0.0033421125519009589, -0.0035595576285158853, -0.0037561780814292555, 
    -0.0039314545152591331, -0.0040850172459846864, -0.0042166335386741496, 
    -0.004326185400481076, -0.0044136482053355117, -0.004479076912385146, 
    -0.0045225896731120414, -0.0045443627753823579, -0.0045446221577415662, 
    -0.0045236441636642578, -0.004481755554156237, -0.0044193347195538865, 
    -0.0043368221257609084, -0.0042347313592526522, -0.0041136607854922709, 
    -0.0039743111296033414, -0.0038175045370855, -0.0036441952621334216, 
    -0.0034554883817250227, -0.0032526512504392831, -0.0030371148746713454, 
    -0.0028104810411510284, -0.0025745106256794786, -0.0023311108444316617, 
    -0.002082314334834683, -0.0018302581451163772, -0.0015771550685539002, 
    -0.0013252641860515898, -0.0010768566355826127, -0.0008341821646780681, 
    -0.00059942973261338278, -0.00037469208847478223, 
    -0.00016192617823543968, 3.7087453730953836e-05, 0.0002207746413588383, 
    0.00038779906937129119, 0.00053708204678850984, 0.00066781432163811195, 
    0.00077946032723962575, 0.00087174848057135852, 0.00094465956683112504, 
    0.00099840693966827469, 0.0010334111012130771, 0.0010502791013853421, 
    0.0010497789912362868, 0.0010328207407903044, 0.0010004431416678939, 
    0.00095379603464699017, 0.0008941236091026594, 0.00082273271999584263, 
    0.00074096235810346047, 0.00065013631501416303, 0.00055151911919060399, 
    0.00044628085474327612, 0.00033546842468265569, 0.00021999191818803591, 
    0.00010062213968727311, -2.1999559718085154e-05, -0.00014734564646752717, 
    -0.00027498096870465515, -0.00040454202862848134, 
    -0.00053571460595010548, -0.00066821051911385696, 
    -0.00080174964757592467, -0.00093603695076864329, -0.0010707451672381317, 
    -0.0012054900257626544, -0.0013398173754256232, -0.0014731837008367856, 
    -0.0016049482183099625, -0.0017343678531289469, -0.0018605947427892567, 
    -0.0019826828495269266, -0.0020995984115921846, -0.0022102377073564806, 
    -0.0023134546462927254, -0.0024080855960626458, -0.0024929826885530747, 
    -0.0025670446934924307, -0.0026292430501069601, -0.0026786458574935591, 
    -0.0027144377267142839, -0.0027359343096398812, -0.0027425944760653626, 
    -0.0027340344634968748, -0.002710036055819568, -0.0026705590054927524, 
    -0.002615756131518686, -0.0025459738607349945, -0.0024617600934732789, 
    -0.0023638603636590605, -0.0022532067451752585, -0.0021309029177814108, 
    -0.001998201061467769, -0.0018564697320301781, -0.0017071628890720631, 
    -0.0015517844514280632, -0.0013918569875997909, -0.001228893123462201, 
    -0.0010643745547453008, -0.00089974019200928304, -0.00073637353353698024, 
    -0.00057559884387150379, -0.00041867480903045023, 
    -0.00026679441712836049, -0.00012107449978450676, 1.7449503190901363e-05, 
    0.00014783268680016283, 0.00026922878714884978, 0.00038089919490948051, 
    0.00048222053525720689, 0.00057268924270069725, 0.00065192732217595709, 
    0.00071968895040561045, 0.0007758619410231294, 0.00082047164419651777, 
    0.00085368309639142961, 0.00087579655772953722, 0.00088724616016426343, 
    0.00088859285205047001, 0.00088051711361348997, 0.00086380475749101384, 
    0.00083933252298543841, 0.00080805463295343109, 0.00077097042504596744, 
    0.00072910258508045395, 0.0006834685709392437, 0.00063505047446401383, 
    0.00058477499455936968, 0.00053349236173290578, 0.00048196945907565499, 
    0.0004308820291138558, 0.00038081319634508388, 0.00033226257495829457, 
    0.00028565310220388047, 0.00024134659336332216, 0.00019966456481369227, 
    0.00016091182241127793, 0.0001254003075712409, 9.3467227929707841e-05, 
    6.5486875663117337e-05, 4.1869245072755656e-05, 2.3057006247652494e-05, 
    9.5016058785770058e-06, 1.6406891670571201e-06, -1.3368742988484568e-07, 
    4.4929625046181354e-06, 1.5723728608491129e-05, 3.3621194513569662e-05, 
    5.809071845090077e-05, 8.8863949292598799e-05, 0.00012550258183546877, 
    0.00016740612278212281, 0.00021382465330667925, 0.0002638828992382429, 
    0.00031660886944334974, 0.00037096340113125997, 0.00042587416143794946, 
    0.00048027417851105646, 0.00053313611156256087, 0.00058350899201175057, 
    0.00063054730727543651, 0.000673533451921667, 0.00071190561431234902, 
    0.00074526514821904777, 0.00077339117154960331, 0.00079624310459968208, 
    0.00081396474987391213, 0.00082688150513372902, 0.00083549734910818598, 
    0.00084048854525742127, 0.00084269336123018405, 0.00084309235451229879, 
    0.00084278159557901516, 0.00084294029740102821, 0.00084479227207628004, 
    0.0008495603872025971, 0.00085841810033045033, 0.00087244330172687545, 
    0.00089256726718738456, 0.00091953179104805173, 0.00095385534235889946, 
    0.00099580428859994785, 0.001045380865376784, 0.0011023133989238021, 
    0.001166060199684095, 0.0012358189532544602, 0.0013105424339417231, 
    0.0013889596906555095, 0.0014695972202735277, 0.0015508122519050723, 
    0.0016308270919064684, 0.0017077667500776316, 0.0017797086283950065, 
    0.0018447258603289242, 0.0019009358359114573, 0.0019465486302663285, 
    0.0019799104316007175, 0.0019995414943050965, 0.0020041723716301709, 
    0.001992771445613252, 0.0019645648484612464, 0.0019190555966558664, 
    0.0018560307288496732, 0.0017755579111652941, 0.0016779808061148207, 
    0.0015638993251734107, 0.0014341468194568744, 0.0012897581794158017, 
    0.0011319365035194577, 0.00096202069789394636, 0.00078144601865996353, 
    0.0005917084354997074, 0.0003943245099700815, 0.00019079817140958634, 
    -1.7418233038808236e-05, -0.0002289538411299029, -0.00044254006444980205, 
    -0.00065702885596979812, -0.00087139305397255682, -0.0010847261860695739, 
    -0.0012962283131496221, -0.0015051931663243626, -0.0017109852967048971, 
    -0.0019130271836018621, -0.0021107886154850455, -0.0023037808078561249, 
    -0.0024915611617043029, -0.0026737373260979375, -0.0028499780971413752, 
    -0.0030200225424441437, -0.0031836902173704809, -0.0033408796948973239, 
    -0.0034915732841808511, -0.0036358321872368288, -0.0037737943971915774, 
    -0.0039056752338701229, -0.0040317589271952111, -0.0041524030934923335, 
    -0.0042680372081795783, -0.0043791590441064282, -0.0044863357509455741, 
    -0.0045901946363782172, -0.0046914146780186348, -0.0047907057874286701, 
    -0.0048887920788268438, -0.0049863831485733034, -0.0050841531234048394, 
    -0.0051827171141955852, -0.0052826156011464278, -0.005384304163047143, 
    -0.0054881472141291984, -0.0055944187236853142, -0.005703301879680444, 
    -0.0058148933780438243, -0.0059291988048920021, -0.006046134692821452, 
    -0.0061655195631279925, -0.0062870761471226447, -0.0064104211948891989, 
    -0.0065350699059544574, -0.0066604404402328191, -0.0067858620857606591, 
    -0.0069105904981425536, -0.0070338303551630054, -0.0071547558132253868, 
    -0.0072725368120647718, -0.0073863643017906292, -0.0074954759693079461, 
    -0.0075991699573233753, -0.0076968274481260838, -0.0077879257098225968, 
    -0.0078720551270149187, -0.0079489304823916491, -0.0080184084688708981, 
    -0.0080804877140990376, -0.0081353187051760277, -0.008183193487402091, 
    -0.0082245321808198536, -0.0082598565457875171, -0.0082897624300518353, 
    -0.008314885803658037, -0.0083358686678659671, -0.00835332877055627, 
    -0.0083678332332883364, -0.0083798801531684546, -0.0083898839411355175, 
    -0.0083981746866612864, -0.0084050062868446518, -0.0084105826111559954, 
    -0.00841509204036495, -0.0084187403184368872, -0.0084217838933289789, 
    -0.0084245575332874169, -0.0084274878867502921, -0.008431100917905443, 
    -0.0084360133303717031, -0.0084429144753381587, -0.0084525283437701625, 
    -0.0084655759641402775, -0.0084827266764546608, -0.0085045616600610847, 
    -0.0085315318172045802, -0.00856393167001465, -0.0086018799004538449, 
    -0.0086453100034907613, -0.008693960568671763, -0.0087473806682144672, 
    -0.0088049334056448259, -0.0088658004502723646, -0.0089290065549364975, 
    -0.0089934355957522333, -0.0090578675623550556, -0.0091210161858186287, 
    -0.0091815786065331216, -0.00923828222878453, -0.0092899349871321327, 
    -0.0093354600853268275, -0.0093739288496664901, -0.0094045768813909424, 
    -0.0094268083142188541, -0.0094401966849064281, -0.0094444744591628341, 
    -0.0094395122830734177, -0.009425305919866251, -0.0094019474848710434, 
    -0.0093695993749968003, -0.0093284528182917843, -0.0092787022984960003, 
    -0.0092205119618038508, -0.0091539852300151943, -0.0090791505877976242, 
    -0.0089959433088023406, -0.0089042027080238444, -0.0088036796363250448, 
    -0.0086940536096930063, -0.0085749539219898384, -0.008445991575887539, 
    -0.0083067925351292555, -0.0081570286227185158, -0.0079964527279071402, 
    -0.0078249159666146494, -0.007642389240946736, -0.0074489749679417195, 
    -0.0072449036791173036, -0.0070305300787928257, -0.0068063340114769043, 
    -0.0065729049383376316, -0.0063309496551957768, -0.0060812572021511063, 
    -0.0058246791340046946, -0.0055620805936539468, -0.005294291853645279, 
    -0.0050220680689231269, -0.0047460606645115941, -0.0044668039170800587, 
    -0.0041847125927285591, -0.0039001054902177614, -0.0036132215463881533, 
    -0.0033242413024662043, -0.0030333129039026908, -0.0027405721873918149, 
    -0.0024461675242502699, -0.0021502770108916863, -0.001853142015801031, 
    -0.0015550837477009373, -0.0012565347343116238, -0.00095805182452863961, 
    -0.00066033644448838639, -0.00036424340680914463, 
    -7.0790025405220928e-05, 0.00021885493570983125, 0.00050338049642967547, 
    0.00078135738529545049, 0.0010512654719950403, 0.0013115341986688707, 
    0.0015605728073279253, 0.0017968048476428781, 0.0020186857467418334, 
    0.0022247232974388765, 0.0024134805703470716, 0.0025835831843112052, 
    0.0027337148047421982, 0.0028626264296074183, 0.0029691448959822428, 
    0.0030521868911900238, 0.0031107740106094475, 0.0031440375773983424, 
    0.0031512324745030696, 0.0031317401773645554, 0.003085069574544917, 
    0.0030108649766486511, 0.0029089201039271761, 0.002779182622539381, 
    0.0026217787247123652, 0.0024370231982755179, 0.0022254316540988098, 
    0.0019877264741843723, 0.0017248293867819996, 0.0014378577811349521, 
    0.0011280940188045955, 0.00079697058919803512, 0.00044604948605598161, 
    7.6999008229561495e-05, -0.00030842767623391685, -0.00070841283094285246, 
    -0.0011210837580532993, -0.0015445412810696497, -0.0019768787100911244, 
    -0.0024162033822540509, -0.0028606602539060356, -0.0033084461357592047, 
    -0.003757830921359403, -0.0042071629146368163, -0.0046548787608879849, 
    -0.0050994986173735716, -0.005539617258590394, -0.0059738953511549375, 
    -0.006401037056018727, -0.0068197822039229418, -0.00722889785971361, 
    -0.0076271766426747566, -0.0080134441966282829, -0.0083865687182028449, 
    -0.0087454713992441944, -0.0090891333603251561, -0.0094166084994175576, 
    -0.0097270290417337951, -0.010019609382829321, -0.010293649310281799, 
    -0.010548534362178143, -0.010783736734750898, -0.010998814546856212, 
    -0.011193415701572295, -0.011367275611530335, -0.011520223945370885, 
    -0.011652184708293052, -0.01176318674660856, -0.011853363937866429, 
    -0.011922963458582235, -0.011972344897664779, -0.012001982953887413, 
    -0.0120124611142397, -0.012004461382830291, -0.011978744158347104, 
    -0.011936121316386668, -0.01187742369382932, -0.011803467411258029, 
    -0.011715020018730723, -0.011612778040049582, -0.01149734427396459, 
    -0.011369213702869354, -0.011228772676985488, -0.011076297323451693, 
    -0.010911966052498929, -0.010735865754815355, -0.010548020171916715, 
    -0.010348408050482627, -0.010136988818318902, -0.0099137342666293267, 
    -0.0096786585074254364, -0.0094318377675287213, -0.0091734443763131623, 
    -0.0089037698233690975, -0.00862324844473061, -0.0083324782676875223, 
    -0.0080322297338571158, -0.0077234611917339699, -0.0074073204945476418, 
    -0.0070851390476886775, -0.0067584298484641816, -0.0064288714545823328, 
    -0.0060982874167660808, -0.0057686259377211216, -0.0054419252889376215, 
    -0.0051202838770973676, -0.0048058240651338499, -0.0045006495746346574, 
    -0.0042068199215273983, -0.0039263162050671698, -0.0036610240378765232, 
    -0.0034127163916826287, -0.0031830479531263392, -0.0029735553923707866, 
    -0.0027856501016693077, -0.0026206222734276793, -0.0024796233053959189, 
    -0.0023636570892141846, -0.0022735531454323664, -0.0022099463487823736, 
    -0.0021732529056287266, -0.0021636446879613014, -0.0021810320001238244, 
    -0.0022250493684767927, -0.0022950588007754555, -0.0023901534908238641, 
    -0.0025091827756116357, -0.0026507726657756386, -0.0028133631019384899, 
    -0.002995247609471458, -0.0031946063177534572, -0.0034095444521089965, 
    -0.0036381402906065087, -0.0038784775488317556, -0.0041287004180658154, 
    -0.0043870617260896496, -0.0046519622334521508, -0.0049219758171505229, 
    -0.0051958648479264085, -0.0054725655022107101, -0.005751164394941841, 
    -0.0060308606207400764, -0.0063109338645055543, -0.0065907086670648042, 
    -0.0068695234608426806, -0.007146712327567235, -0.0074215752630494717, 
    -0.0076933890836013959, -0.0079613886739410295, -0.008224775323599413, 
    -0.0084827270871005132, -0.0087344069092456789, -0.0089789854743043598, 
    -0.0092156586230445949, -0.0094436802802068415, -0.0096623820724784926, 
    -0.0098712134565589905, -0.010069770973488318, -0.010257823968485796, 
    -0.010435349648914233, -0.010602547428280529, -0.010759839184202711, 
    -0.010907858671871383, -0.011047413477794704, -0.011179440887194076, 
    -0.011304938864894221, -0.011424905241518164, -0.011540279190584564, 
    -0.011651876368142076, -0.01176036544758499, -0.011866242457558809, 
    -0.011969822384031346, -0.012071258713644208, -0.012170561147980525, 
    -0.012267617459486707, -0.012362236690077241, -0.012454149337467097, 
    -0.012543021521698566, -0.012628434962172416, -0.012709866918908691, 
    -0.012786663431877489, -0.012858027991227898, -0.012923003716812429, 
    -0.01298049159172498, -0.013029257737306984, -0.013067952914810645, 
    -0.013095139946184794, -0.013109309038078972, -0.013108900283425358, 
    -0.013092319656364546, -0.013057971022659532, -0.013004291536473211, 
    -0.012929779459622081, -0.012833048076183018, -0.01271287684303346, 
    -0.012568252096217232, -0.012398433068968932, -0.012202983667464806, 
    -0.011981817026397111, -0.011735220543833283, -0.011463877257597543, 
    -0.011168871434216462, -0.010851689315972029, -0.01051419752458854, 
    -0.010158619688466618, -0.0097874940212178078, -0.0094036319115062758, 
    -0.0090100568379720327, -0.0086099276136146277, -0.0082064646208426881, 
    -0.0078028359933601452, -0.0074020403062543781, -0.0070067814743106716, 
    -0.0066193451401205909, -0.0062415023709101614, -0.0058744417582075924, 
    -0.0055187716540916988, -0.0051745618032970099, -0.0048414501005902173, 
    -0.0045187890856907501, -0.0042057779916367223, -0.0039015998213895245, 
    -0.0036054802917614213, -0.0033167182801888727, -0.0030346745438544669, 
    -0.002758761153221741, -0.002488408107019442, -0.0022230477565909064, 
    -0.0019621018260215081, -0.0017049910006660303, -0.0014511481285864806, 
    -0.001200063725281753, -0.00095132309823782533, -0.00070468646360941393, 
    -0.00046012818500195041, -0.00021789919628973891, 2.1467886489441149e-05, 
    0.00025715716280206116, 0.00048810587409882437, 0.00071306686814598104, 
    0.00093067676159736814, 0.001139533013014032, 0.0013382691485763726, 
    0.0015256236348135973, 0.0017004909779584295, 0.0018619675666090582, 
    0.0020093899400306214, 0.0021423509374771501, 0.0022607117335715181, 
    0.0023645990040357758, 0.0024543888987894101, 0.0025306847914967215, 
    0.002594281938579383, 0.0026461266645272158, 0.0026872638062840691, 
    0.0027187998078278272, 0.0027418569749454308, 0.0027575278004847068, 
    0.0027668571123902492, 0.0027708228626635843, 0.0027703291474187063, 
    0.0027661959018411334, 0.0027591656875670468, 0.0027498925583956703, 
    0.002738938555156307, 0.0027267805338370044, 0.0027138039830954786, 
    0.0027003064011056131, 0.0026865105899231958, 0.0026725589793656222, 
    0.0026585169064607911, 0.0026443686177521782, 0.0026300112062152639, 
    0.0026152454709035514, 0.0025997705080311848, 0.002583175019114228, 
    0.0025649271024971326, 0.002544371160758477, 0.0025207179629125761, 
    0.0024930539281332355, 0.0024603719244311486, 0.0024216405439922615, 
    0.0023758917635079389, 0.0023223097561878626, 0.0022603049062152503, 
    0.002189568861828437, 0.0021100795993894209, 0.0020221066141420051, 
    0.0019261919506422432, 0.0018231349121210214, 0.0017139631092049675, 
    0.0015998984157570314, 0.0014823376508820451, 0.0013627962962111588, 
    0.0012428789925182687, 0.0011242235518679619, 0.0010084716492849408, 
    0.00089721904013811114, 0.00079199347019258751, 0.00069424052888548114, 
    0.00060531203671026059, 0.00052645931955753707, 0.00045883786375527447, 
    0.0004034872977409614, 0.00036131896369564977, 0.00033309984045919459, 
    0.00031943737917987603, 0.0003207684522201175, 0.00033737674690393195, 
    0.00036940034875278737, 0.00041687475851182639, 0.00047975622785620159, 
    0.00055795386390292069, 0.00065136780193498893, 0.00075989951340372402, 
    0.00088344625500097614, 0.0010219012566862924, 0.0011750980953684105, 
    0.0013427591992273781, 0.0015244414285528814, 0.0017194849202417234, 
    0.0019269829473857792, 0.0021457767666907658, 0.0023744710446790373, 
    0.0026114772926639539, 0.0028550631628126775, 0.0031034159037019397, 
    0.0033547127781629257, 0.003607179887081995, 0.0038591502156889467, 
    0.0041090903628893619, 0.0043556112563544478, 0.0045974654275971662, 
    0.0048335052684761633, 0.0050626592912544899, 0.0052839032678324432, 
    0.0054962080091216113, 0.0056985441687606711, 0.0058898741126344745, 
    0.0060691628212168934, 0.0062353964455876074, 0.0063875956940126488, 
    0.0065248312073465497, 0.0066462202251457115, 0.0067509330194471971, 
    0.0068382007157141763, 0.0069073025279249353, 0.0069575932995422666, 
    0.0069885195196739188, 0.006999655772648424, 0.0069907327237782079, 
    0.0069616797229374089, 0.0069126364763807888, 0.0068439646043934495, 
    0.0067562408164781396, 0.0066502403670976118, 0.0065269140088309047, 
    0.0063873355872971936, 0.0062326877431367377, 0.0060642133480161564, 
    0.0058831819085041594, 0.005690852224745929, 0.0054884197744253715, 
    0.0052769927695312611, 0.0050575679311109564, 0.0048310338583642401, 
    0.0045981689102491874, 0.0043596447406616971, 0.0041160586232289664, 
    0.0038679421205198841, 0.0036158218233951424, 0.0033602615318339656, 
    0.003101926250916463, 0.0028416607515647277, 0.0025805236543294994, 
    0.0023198531976935111, 0.0020612781438624286, 0.0018067490987875628, 
    0.0015585224008837226, 0.0013191465603017449, 0.0010914103752158871, 
    0.00087827684983586823, 0.00068279405378095519, 0.00050798826020939073, 
    0.00035676011299978582, 0.00023175653200978037, 0.00013527319256763354, 
    6.915999090864952e-05, 3.4749224514981099e-05, 3.2801352311967482e-05, 
    6.3482651882239364e-05, 0.00012634204195100486, 0.00022034118194561332, 
    0.00034386924988949377, 0.00049480383416877511, 0.00067056857389549696, 
    0.00086820447442816594, 0.0010844506541646147, 0.0013158353319107311, 
    0.0015587530784715524, 0.0018095682923404931, 0.0020647168315941124, 
    0.0023207891432257409, 0.0025746106546681159, 0.0028233133628794657, 
    0.0030643732257138647, 0.003295618511041736, 0.0035152127832765003, 
    0.0037216019441987267, 0.0039134681574187835, 0.0040896552038622736, 
    0.0042491227626736171, 0.0043909106488660768, 0.0045141128368975077, 
    0.0046178663057264892, 0.004701372604699704, 0.0047638898574302348, 
    0.0048047288450038649, 0.0048232510787658174, 0.0048188457179652927, 
    0.0047909150085589857, 0.0047388729598922992, 0.0046621146470765045, 
    0.0045600138276726048, 0.004431928926079267, 0.0042772034237058805, 
    0.0040951922366329243, 0.0038853052453988123, 0.0036470677442462279, 
    0.0033801941233866212, 0.0030846530445545108, 0.0027607209466652726, 
    0.0024090287806629047, 0.0020305906980382293, 0.001626833599914592, 
    0.0011996066508771924, 0.00075123250174224672, 0.00028450950290276957, 
    -0.00019726598936214201, -0.00069028990425792349, -0.001190268645364422, 
    -0.0016924571716264009, -0.0021917449208869125, -0.0026827245671800777, 
    -0.0031598433251303812, -0.0036175129118864277, -0.0040502433563254572, 
    -0.0044527818197378395, -0.0048202208045835136, -0.005148096419208441, 
    -0.005432456351181305, -0.0056699177093525299, -0.0058577114339996832, 
    -0.0059936813725858544, -0.006076318312747628, -0.0061047492914576536, 
    -0.0060787337131226167, -0.0059986753500415367, -0.0058656257972024752, 
    -0.0056812880367485379, -0.0054480299624936786, -0.0051688615994320286, 
    -0.0048474384741999032, -0.0044880388682208916, -0.0040955020349269832, 
    -0.0036751729492128411, -0.0032328207712354769, -0.0027745405547106275, 
    -0.0023066376265908927, -0.0018355102789661692, -0.0013675246742507303, 
    -0.00090889278144211817, -0.00046554505095655954, 
    -4.3048683046410921e-05, 0.00035346533039701348, 0.0007193702033693423, 
    0.0010505505494720596, 0.0013434250570258683, 0.001594945652453531, 
    0.0018025933468983051, 0.0019644014838287585, 0.002078972093630416, 
    0.0021454719268708092, 0.0021636287379454226, 0.0021337311771760419, 
    0.0020565910180133646, 0.0019335080844082213, 0.0017662354737564452, 
    0.0015569317731710325, 0.0013080925992942369, 0.0010224619483925376, 
    0.0007029516379731455, 0.00035252763848164879, -2.5905465892944897e-05, 
    -0.00042955408904270622, -0.00085574670405342461, -0.0013018677473103342, 
    -0.0017652505376974032, -0.0022430310902162411, -0.0027319994461259146, 
    -0.0032284962633866653, -0.0037283668279749294, -0.0042270693510727177, 
    -0.0047198127150535193, -0.0052018640123512134, -0.005668781069103024, 
    -0.0061166323685723804, -0.0065420581222128127, -0.0069422909758306379, 
    -0.0073151194388965017, -0.0076588446757558642, -0.0079722590990484715, 
    -0.0082546688584256636, -0.0085058581944733383, -0.0087261024545718709, 
    -0.0089161041477292032, -0.0090769671753376489, -0.0092100862202363597, 
    -0.009317071066490306, -0.0093996471880870552, -0.0094595659257328078, 
    -0.0094985269460017268, -0.0095181398469364638, -0.0095198558878291269, 
    -0.009504987820652901, -0.0094747210190518471, -0.0094301273160511869, 
    -0.0093721942583418327, -0.0093018882395227657, -0.0092201818163475946, 
    -0.0091280831055510873, -0.0090266965476320377, -0.0089172025032160773, 
    -0.008800906478470906, -0.0086792070191466699, -0.008553629374203375, 
    -0.0084257858970383601, -0.0082973806478734043, -0.0081702281363942204, 
    -0.0080462380159685258, -0.0079273525459726702, -0.0078154916146856504, 
    -0.0077124497137940617, -0.0076198248685081186, -0.0075389843304684142, 
    -0.0074710716375678459, -0.007417066937505136, -0.0073778713813718718, 
    -0.0073544577859121652, -0.0073479812266827203, -0.0073598922272905534, 
    -0.007392009886702436, -0.0074465081940113149, -0.0075258818729040432, 
    -0.0076327977730639585, -0.0077699234107578268, -0.0079396632459250577, 
    -0.0081439020464234638, -0.0083837297055343388, -0.0086592487707981766, 
    -0.0089694586109978318, -0.0093121769827898479, -0.0096841269294670827, 
    -0.010081003592430002, -0.010497637411083687, -0.010928170607281318, 
    -0.011366249281229257, -0.011805243882802441, -0.012238451732504018, 
    -0.012659288388339865, -0.013061422735326449, -0.013438945926971077, 
    -0.013786405254067274, -0.014098880027932581, -0.014371950610721515, 
    -0.014601725167251662, -0.014784821686812371, -0.014918431403585331, 
    -0.015000390407310634, -0.015029310643611564, -0.015004654053014941, 
    -0.014926750777099288, -0.014796785708837698, -0.014616677497619357, 
    -0.014388920134675976, -0.014116424389743776, -0.013802403157419442, 
    -0.013450181505375802, -0.013063125306221741, -0.012644563414757599, 
    -0.012197770497393685, -0.011725928844186552, -0.011232172223060829, 
    -0.010719623415784498, -0.010191477554057275, -0.0096510737249684096, 
    -0.009101950149762424, -0.0085478439798397764, -0.00799265627741573, 
    -0.0074403146154043412, -0.0068946091441891531, -0.006358963741152036, 
    -0.0058361780405384572, -0.0053282003219599847, -0.0048359507420658605, 
    -0.0043592003652411929, -0.0038965550866570764, -0.0034455956644547066, 
    -0.0030030152140732864, -0.0025648406840527507, -0.0021266620554633484, 
    -0.0016839122611922398, -0.0012320367197869177, -0.00076671537193430275, 
    -0.00028401946134783802, 0.00021939395738283129, 0.00074622704125438838, 
    0.0012983564882515048, 0.0018766933885496192, 0.0024811172916693099, 
    0.0031102632738388316, 0.0037614252969290804, 0.004430467533311418, 
    0.0051117412744247949, 0.0057980704206473752, 0.0064808705408774623, 
    0.0071502870742619412, 0.0077954730970536991, 0.0084051327783959077, 
    0.0089679655241572866, 0.0094733608142816596, 0.0099120450014633255, 
    0.010276685240349573, 0.0105623690668492, 0.010766897787446838, 
    0.010890967898207073, 0.010937870542452707, 0.010913390507744905, 
    0.010825253979522498, 0.010682586536458691, 0.010495328353942101, 
    0.010273434819783401, 0.010026112830279739, 0.0097610878717177465, 
    0.009483720521540567, 0.0091964744440220444, 0.0088983774206857491, 
    0.0085849753052975319, 0.0082485813792186041, 0.0078789919329605353, 
    0.0074641464012479659, 0.006991428533884291, 0.0064488453526089715, 
    0.0058262352016912738, 0.00511625054987133, 0.0043151123816067066, 
    0.0034231492363946381, 0.0024447393983066429, 0.0013880642743215488, 
    0.00026425136752998357, -0.00091323434778068876, -0.0021297738254266903, 
    -0.0033700729235580174, -0.004619392064335686, -0.0058636262518346792, 
    -0.0070904277901963457, -0.0082885825766951509, -0.0094483174857871461, 
    -0.010560815869373028,
  // Fqt-total(4, 0-1999)
    0.99999999999999956, 0.9975779806166567, 0.99036171835243547, 
    0.97849809459360826, 0.9622245338768598, 0.94185885765112731, 
    0.91778619381303317, 0.89044389227843601, 0.86030542365024598, 
    0.8278642226847166, 0.79361832559580303, 0.75805646768911306, 
    0.72164613547370293, 0.68482387190415361, 0.64798793111543296, 
    0.61149325375952002, 0.57564859351694031, 0.54071556756306882, 
    0.50690930564548875, 0.47440042097723401, 0.44331796097632764, 
    0.41375306101852055, 0.38576302540572077, 0.35937559712028722, 
    0.3345932490439536, 0.31139732528895558, 0.28975194434307, 
    0.26960758903124338, 0.25090432728787626, 0.23357465443647574, 
    0.21754595170832725, 0.20274256430726276, 0.18908753849063153, 
    0.17650402909155496, 0.16491641664847181, 0.15425115922895785, 
    0.1444374271199555, 0.13540755005570163, 0.12709731408953565, 
    0.11944615936142229, 0.11239728288721379, 0.10589770228832183, 
    0.099898255392163682, 0.094353584776664806, 0.089222070681518509, 
    0.084465740183586782, 0.080050140823778163, 0.07594418478093154, 
    0.072119966145743133, 0.06855255661469252, 0.065219777750338478, 
    0.06210197052796966, 0.059181750121124255, 0.056443767762762782, 
    0.053874473527794751, 0.05146189151478768, 0.049195404167224802, 
    0.047065552608568276, 0.045063854876058199, 0.043182652165725581, 
    0.041414960412811945, 0.039754353579282017, 0.038194862906895333, 
    0.036730880786082443, 0.035357082509409311, 0.034068353500447214, 
    0.032859721915622621, 0.031726315440419872, 0.030663320088021119, 
    0.029665959804301301, 0.028729493090546541, 0.027849206949090776, 
    0.027020422455289836, 0.026238489402027915, 0.025498789119883389, 
    0.024796733929459368, 0.024127764109605113, 0.023487358063755234, 
    0.022871048134172178, 0.022274447597174819, 0.021693284553124755, 
    0.021123454384311555, 0.020561069706851585, 0.020002524482937857, 
    0.01944455423326534, 0.018884291690342035, 0.018319321530041194, 
    0.01774771750260995, 0.017168068100433, 0.016579477138166109, 
    0.015981562573313259, 0.015374426529850212, 0.014758628978033782, 
    0.014135150870331457, 0.013505350854239163, 0.012870924342508829, 
    0.012233857606538645, 0.011596375978573681, 0.01096088308139459, 
    0.010329905503820137, 0.0097060240734535494, 0.0090918040516946731, 
    0.0084897288911174682, 0.0079021367874169499, 0.0073311693664574931, 
    0.0067787306401680481, 0.0062464638611460579, 0.0057357462949418035, 
    0.0052476978434250468, 0.0047832104571809368, 0.004342989266439474, 
    0.0039276015789136099, 0.0035375394406545204, 0.0031732643135156343, 
    0.0028352591796026025, 0.0025240569165703858, 0.0022402556289705037, 
    0.0019845119379857815, 0.0017575266638072886, 0.0015600214406612353, 
    0.0013927066150579512, 0.0012562552520976929, 0.0011512737487798829, 
    0.0010782842609559158, 0.0010376984989270374, 0.001029804999446636, 
    0.0010547505497611387, 0.001112522691976708, 0.0012029293855421808, 
    0.0013255746690346109, 0.0014798293801904555, 0.001664803362269121, 
    0.0018793104033158145, 0.0021218376831444409, 0.0023905275842385759, 
    0.0026831650961244473, 0.0029971920942563606, 0.0033297292112082892, 
    0.0036776202001631226, 0.0040374871227061796, 0.0044057944826301912, 
    0.0047789186306138954, 0.005153213035570931, 0.0055250744864557937, 
    0.0058909957830098093, 0.0062476078711642151, 0.0065917164312356401, 
    0.0069203205861267103, 0.00723062839270509, 0.0075200646608063254, 
    0.0077862790377503177, 0.0080271397931866561, 0.0082407529470792697, 
    0.0084254637330995266, 0.0085798732150221615, 0.0087028575902567372, 
    0.0087935795718132714, 0.0088515169348713264, 0.0088764737092268398, 
    0.008868607066218127, 0.0088284446494099628, 0.0087569081263918006, 
    0.0086553251729089963, 0.0085254357952088602, 0.0083693843546800845, 
    0.0081896925647447459, 0.0079892165123865259, 0.0077710786634451086, 
    0.0075385976775943489, 0.007295199994095088, 0.0070443459551441032, 
    0.0067894597477128728, 0.0065338703743518462, 0.0062807539554561673, 
    0.0060330892693131717, 0.0057936108291665143, 0.0055647749978074536, 
    0.005348724590417301, 0.005147264106000771, 0.004961840129518536, 
    0.0047935232103263354, 0.0046430054494949243, 0.0045105938783986336, 
    0.0043962226151058985, 0.0042994650539880681, 0.0042195681454542952, 
    0.0041554826900584299, 0.0041059113747965283, 0.0040693577656392924, 
    0.004044183665000858, 0.0040286628282048481, 0.0040210389441368488, 
    0.0040195791925913792, 0.0040226220637042355, 0.0040286203888568279, 
    0.0040361733826852373, 0.0040440545001025029, 0.0040512331231627331, 
    0.0040568788240260643, 0.0040603598098885767, 0.004061228724486869, 
    0.0040592018432179461, 0.004054124946947282, 0.0040459435613931921, 
    0.0040346681340947474, 0.004020342105866952, 0.0040030152275385518, 
    0.003982724390111464, 0.003959481605180221, 0.00393327578366175, 
    0.0039040753105662267, 0.0038718504463498764, 0.0038365966626612369, 
    0.0037983651319514256, 0.003757292346137673, 0.0037136317575701804, 
    0.0036677695674929554, 0.0036202410273357389, 0.0035717140816201023, 
    0.0035229763609125452, 0.0034748889541298547, 0.0034283371801164227, 
    0.0033841687924427359, 0.0033431310010469096, 0.0033058073903345065, 
    0.003272560614500453, 0.0032434874102459685, 0.0032183856192591264, 
    0.0031967411567472071, 0.0031777274369908476, 0.0031602349308761934, 
    0.0031429077890213282, 0.0031242018614119856, 0.0031024566281361637, 
    0.0030759704366754843, 0.00304308260891292, 0.0030022487437440263, 
    0.0029521110169057679, 0.0028915538104959874, 0.002819741768760417, 
    0.0027361423814863338, 0.002640526299106407, 0.0025329467237320061, 
    0.0024137098354152838, 0.0022833249409454481, 0.0021424542408358589, 
    0.0019918497924224453, 0.0018323000117723893, 0.0016645759281008663, 
    0.0014893914910689096, 0.0013073675584150844, 0.0011190198159035107, 
    0.00092475570104163347, 0.00072488456907941344, 0.000519643649571521, 
    0.00030923597877552834, 9.3883253671020911e-05, -0.00012611303559943691, 
    -0.00035030605294319019, -0.00057804406589495225, 
    -0.00080841964898736309, -0.0010402368337488629, -0.0012720048707205594, 
    -0.0015019580354126559, -0.0017280900847783519, -0.0019482050680743434, 
    -0.0021599715240790329, -0.0023609808923928536, -0.0025488016651592678, 
    -0.0027210214924849136, -0.00287529508044431, -0.0030093803538972057, 
    -0.0031211719982435254, -0.0032087370172296289, -0.0032703345577684041, 
    -0.0033044401701138306, -0.0033097576757843842, -0.003285227266825706, 
    -0.0032300329761696749, -0.0031435953146854195, -0.0030255772446035833, 
    -0.002875881285208421, -0.0026946577623685576, -0.0024823075637130515, 
    -0.0022394945756503662, -0.0019671581573483797, -0.0016665266064960053, 
    -0.0013391263814972116, -0.00098679488112740849, -0.00061168595888044244, 
    -0.00021627938305573228, 0.0001966193422643718, 0.00062387686518969819, 
    0.0010620399114772594, 0.0015073484745523728, 0.0019557605088514848, 
    0.0024029832486212673, 0.0028445221132409057, 0.0032757390466333957, 
    0.003691925051903563, 0.0040883838238433929, 0.0044605213886668915, 
    0.0048039446592492013, 0.0051145582297631555, 0.0053886611313829977, 
    0.0056230324809688377, 0.0058150055078933106, 0.005962521810935352, 
    0.0060641676146774952, 0.0061191827279788742, 0.0061274554982066569, 
    0.0060894991299687779, 0.0060064160316073058, 0.0058798533214135217, 
    0.005711943842306136, 0.0055052513684824781, 0.0052627057736959184, 
    0.0049875400540240825, 0.0046832284421293681, 0.0043534242615150039, 
    0.0040018903662160151, 0.0036324277141958363, 0.0032487972691896982, 
    0.0028546336160748384, 0.0024533563577959325, 0.0020480849626010223, 
    0.0016415538338603931, 0.001236057568728571, 0.00083340406194792329, 
    0.00043491567146168022, 4.1458845422395388e-05, -0.00034647728646490674, 
    -0.00072867291186637221, -0.0011050396054491862, -0.001475471950775053, 
    -0.0018397079686453888, -0.0021972207080712502, -0.002547142817359912, 
    -0.0028882263183566451, -0.0032188501181788136, -0.0035370535853197116, 
    -0.0038405985667579754, -0.0041270463057115373, -0.0043938479766608349, 
    -0.0046384451179691802, -0.0048583658456791577, -0.0050513225416358044, 
    -0.0052153002379576284, -0.0053486328357071414, -0.0054500582854411757, 
    -0.0055187657256464571, -0.0055544147597892286, -0.0055571394904628882, 
    -0.0055275365562122911, -0.0054666387666157338, -0.0053758778195913811, 
    -0.0052570352896663458, -0.0051121798990057601, -0.004943600422625944, 
    -0.0047537293772164932, -0.0045450626037627237, -0.0043200829398410247, 
    -0.0040811877942530652, -0.003830626313389741, -0.003570446702876737, 
    -0.0033024549805859009, -0.0030281904851211421, -0.0027489112679198327, 
    -0.0024655918711972255, -0.0021789414377244134, -0.0018894277819061752, 
    -0.0015973166960485906, -0.0013027174371870284, -0.0010056347396763989, 
    -0.00070601549107578555, -0.00040379596609043734, 
    -9.8935575252133811e-05, 0.0002085540115408849, 0.00051858885652667993, 
    0.0008310002939645294, 0.0011455247799185308, 0.0014617997918183745, 
    0.0017793565009482837, 0.0020976161786055107, 0.0024158846564822536, 
    0.002733348181762811, 0.0030490718791858699, 0.0033620022840583621, 
    0.0036709796868372685, 0.0039747487415124341, 0.0042719776643357537, 
    0.0045612771827121187, 0.0048412210851986144, 0.0051103831310642034, 
    0.0053673664972390877, 0.0056108519908449062, 0.0058396369831704795, 
    0.0060526724154802798, 0.0062490948220312965, 0.006428252226539, 
    0.0065897212952787301, 0.0067333193381966137, 0.0068590930800571858, 
    0.0069673091336825022, 0.0070584212486650491, 0.0071330271441442054, 
    0.0071918205415037071, 0.0072355398168469911, 0.0072649152026841787, 
    0.0072806243242782747, 0.0072832546952143751, 0.0072732752636488138, 
    0.007251021591062029, 0.0072166952583636347, 0.0071703627846752861, 
    0.0071119722999368673, 0.0070413662626106072, 0.0069583014297470835, 
    0.0068624704023909373, 0.0067535294129650956, 0.0066311321163683781, 
    0.0064949721597854053, 0.0063448248558183786, 0.006180592889037829, 
    0.006002346381487369, 0.0058103619108953669, 0.0056051505611357461, 
    0.0053874846047722658, 0.0051584089523190645, 0.0049192431030957865, 
    0.0046715731821981221, 0.0044172222245173736, 0.0041582082510231424, 
    0.0038966840974800367, 0.0036348640686504449, 0.0033749544322340197, 
    0.0031190807100455746, 0.0028692290728592816, 0.0026271961267885524, 
    0.0023945604183267075, 0.0021726612069542283, 0.0019626009899024947, 
    0.0017652541925378277, 0.0015812887785815433, 0.0014111908985475854, 
    0.0012552911734666267, 0.001113790150880754, 0.00098677500515616527, 
    0.00087423673951735775, 0.00077607236746839484, 0.00069208369627381066, 
    0.00062196110601156376, 0.00056526342096243276, 0.00052138511734551186, 
    0.00048952579748868413, 0.00046866087563480889, 0.00045752866795340587, 
    0.00045463643696805209, 0.00045828186385225617, 0.00046660344787797836, 
    0.00047763973276336867, 0.00048939789692756892, 0.00049992892831869596, 
    0.00050739493089858563, 0.00051013774308959477, 0.00050673484286316663, 
    0.00049604901839160739, 0.0004772605831197669, 0.00044989500975777923, 
    0.00041382844901188094, 0.000369280340603703, 0.00031679127197851834, 
    0.00025718723574260456, 0.00019153552049546601, 0.00012109099174847847, 
    4.7241538724543142e-05, -2.8545220847143059e-05, -0.00010478114794467702, 
    -0.00018000718845107876, -0.00025284802742357769, 
    -0.00032205743924764471, -0.00038656099363925051, 
    -0.00044549043405036715, -0.00049821580477057525, 
    -0.00054436216026702627, -0.00058383164318591874, 
    -0.00061680173082995671, -0.00064372894317989366, 
    -0.00066533616022090782, -0.00068258066515137703, 
    -0.00069662647268701073, -0.0007087845483623017, -0.00072045778371995436, 
    -0.00073307242562252125, -0.00074801791276835918, 
    -0.00076658775435799209, -0.00078993953711577669, 
    -0.00081906159630991643, -0.00085475324097837872, 
    -0.00089761418969428223, -0.00094804458654436136, -0.001006243649419364, 
    -0.001072220423256503, -0.0011458002095181415, -0.0012266371052851921, 
    -0.0013142276637871299, -0.0014079364424167346, -0.0015070235496384607, 
    -0.0016106723448071983, -0.001718021567353085, -0.001828181239914512, 
    -0.0019402398830226225, -0.0020532621149873236, -0.0021662800587580969, 
    -0.0022782814414050011, -0.002388204078332231, -0.0024949349412385757, 
    -0.0025973132788895026, -0.0026941469537721543, -0.0027842268884455588, 
    -0.0028663424393123847, -0.0029392996489318634, -0.003001934403094075, 
    -0.0030531251658796328, -0.0030918065334942769, -0.0031169737029176771, 
    -0.0031276974638935252, -0.0031231456708991478, -0.0031026204289633348, 
    -0.0030656006274165765, -0.0030117985688585844, -0.002941207561419652, 
    -0.0028541355395880069, -0.0027512292766414025, -0.0026334785725628624, 
    -0.002502202445373294, -0.0023590175546822551, -0.0022057878060391368, 
    -0.0020445561531072889, -0.0018774637108757313, -0.0017066552166380619, 
    -0.0015341831555029874, -0.0013619146301665024, -0.0011914423217324708, 
    -0.0010240048018782403, -0.0008604258267274885, -0.00070106523185308443, 
    -0.00054579765746267078, -0.00039400696142093361, 
    -0.00024461324607107115, -9.6111387343225936e-05, 5.336329479956737e-05, 
    0.00020595437457279458, 0.00036399672928248727, 0.00052991354979833665, 
    0.00070610996463677965, 0.00089486629117845181, 0.0010982289987310988, 
    0.0013179116085030493, 0.0015552026050839277, 0.0018108908594257477, 
    0.0020852074738081502, 0.002377786290054282, 0.0026876457790348759, 
    0.0030131918737304904, 0.003352239915985569, 0.0037020534449578447, 
    0.0040594114371940871, 0.0044206908063500637, 0.0047819592853902641, 
    0.0051390917844757068, 0.0054878850016510453, 0.0058241781451111438, 
    0.006143968647813869, 0.0064435125178086503, 0.0067194173411235314, 
    0.0069687157883513316, 0.0071889184236849169, 0.0073780527676874383, 
    0.0075346770763401972, 0.0076578860606333551, 0.0077472889601596781, 
    0.0078029777157915528, 0.0078254826543238103, 0.0078157235063302972, 
    0.0077749445174062305, 0.0077046608234144906, 0.0076065886704330182, 
    0.0074825923243383493, 0.0073346242267217166, 0.0071646784486557652, 
    0.0069747540061612214, 0.0067668261417772385, 0.0065428354320117054, 
    0.0063046864462295033, 0.0060542625683008573, 0.0057934433674998445, 
    0.0055241287753558434, 0.0052482617097497986, 0.0049678452293590728, 
    0.0046849520909266222, 0.0044017244328260451, 0.0041203678737047845, 
    0.0038431330772745308, 0.0035722956261830911, 0.0033101237480517654, 
    0.003058848154041254, 0.00282062497241482, 0.0025974991461968143, 
    0.0023913682468450124, 0.0022039473866126234, 0.0020367375995343075, 
    0.0018909983336015967, 0.0017677270151194989, 0.001667640218000474, 
    0.0015911670584131819, 0.0015384396788148365, 0.0015092909041352096, 
    0.0015032553678427903, 0.0015195708963569793, 0.0015571855683606901, 
    0.0016147600109083745, 0.0016906769753519053, 0.0017830531364907657, 
    0.0018897505847375157, 0.0020083966417880831, 0.0021364124473335615, 
    0.0022710430646054607, 0.0024093960774252284, 0.0025484805300625764, 
    0.0026852509887221976, 0.0028166475483428649, 0.0029396490395887653, 
    0.0030513137084721103, 0.0031488374944755111, 0.0032296003512341676, 
    0.0032912264678278962, 0.0033316417867623447, 0.0033491301495925337, 
    0.0033423860914320886, 0.0033105567778240331, 0.0032532736411533679, 
    0.0031706647417553777, 0.0030633528027943107, 0.0029324291959520149, 
    0.0027794167382665515, 0.0026062266986531224, 0.0024151000764166481, 
    0.0022085590058347556, 0.001989347569551192, 0.0017603812742607616, 
    0.0015246879092226709, 0.0012853530424645073, 0.0010454593365986406, 
    0.000808028015454621, 0.00057595642945547582, 0.00035195530668794927, 
    0.00013849163295367103, -6.2266144776349698e-05, -0.00024849998356729972, 
    -0.0004187767859758225, -0.00057207446347320133, -0.00070778735722472059, 
    -0.00082571210162854384, -0.0009260172651266754, -0.0010091887079076891, 
    -0.0010759706711933879, -0.0011272909071889754, -0.0011641890034816095, 
    -0.0011877512912303999, -0.0011990628696809341, -0.0011991747283661553, 
    -0.0011890994570922012, -0.0011698203279349201, -0.001142325880514409, 
    -0.0011076463552872004, -0.0010669020977047221, -0.0010213458469777201, 
    -0.00097240366179726753, -0.00092170438577587606, 
    -0.00087108584844718172, -0.00082259074656831606, 
    -0.00077843226472997765, -0.00074093348570506128, 
    -0.00071245099875425746, -0.00069528627025656163, 
    -0.00069159197210191987, -0.00070327791988695706, 
    -0.00073193612038739057, -0.00077877214694246747, 
    -0.00084455866270893984, -0.00092959633841842564, -0.0010337051441545399, 
    -0.0011562176699797375, -0.0012959975355102465, -0.001451461583675857, 
    -0.0016206315451431463, -0.0018011912450953439, -0.0019905705596963484, 
    -0.0021860319429652351, -0.0023847629382870825, -0.0025839570094446829, 
    -0.0027808835910868622, -0.0029729488421646202, -0.0031577316031390127, 
    -0.0033330241077485193, -0.0034968373101176928, -0.0036474211246780401, 
    -0.0037832593828551198, -0.0039030751549748825, -0.0040058270669543631, 
    -0.0040907003585958874, -0.004157108799051722, -0.0042046779669472484, 
    -0.0042332355679876128, -0.0042427948025871463, -0.0042335329818983291, 
    -0.004205770853399131, -0.0041599465586440489, -0.0040966036828333696, 
    -0.0040163721989338787, -0.0039199663362782817, -0.0038081854071242882, 
    -0.0036819191229232342, -0.0035421579082167364, -0.0033900057196603831, 
    -0.0032266937177426536, -0.0030535813140068536, -0.0028721679257412537, 
    -0.002684093362500699, -0.0024911318948398643, -0.0022951849797086402, 
    -0.002098261639390888, -0.0019024574818312843, -0.0017099147165733394, 
    -0.0015227819333105538, -0.0013431609505636904, -0.0011730508527565192, 
    -0.00101429382183437, -0.00086852858767779751, -0.00073715452134108809, 
    -0.00062131264817347296, -0.00052188201284518486, 
    -0.00043950065800164314, -0.0003745955318675483, -0.00032742555670680907, 
    -0.0002981264668399138, -0.000286751475866002, -0.00029329803853576474, 
    -0.00031772463362414813, -0.00035995976920947024, -0.0004198971805240919, 
    -0.00049738016220973312, -0.00059217527151825874, 
    -0.00070393919379121972, -0.00083218820081700027, 
    -0.00097626537601716362, -0.0011353259712938977, -0.0013083281994378548, 
    -0.0014940325044212402, -0.0016910127753523901, -0.0018976733643028844, 
    -0.0021122743224408626, -0.0023329645275600047, -0.0025578131583002222, 
    -0.0027848481033401471, -0.0030120833789153484, -0.0032375490783270733, 
    -0.0034593090181028732, -0.0036754686852724181, -0.0038841788391333837, 
    -0.0040836191855493286, -0.0042719916101718082, -0.0044474994832639876, 
    -0.0046083412526938374, -0.0047527058901822962, -0.004878777419894142, 
    -0.004984746144747876, -0.0050688267917824046, -0.0051292832163411838, 
    -0.0051644543398458457, -0.005172788426256532, -0.0051528791000708474, 
    -0.0051035083952520044, -0.0050236905676928796, -0.0049127244099106699, 
    -0.0047702378874348791, -0.0045962348284438086, -0.0043911284915289671, 
    -0.0041557688124013873, -0.0038914513395395451, -0.0035999092536844993, 
    -0.0032833028380595047, -0.0029441860942269562, -0.0025854778411573396, 
    -0.0022104217814688729, -0.0018225529044411503, -0.0014256553651429212, 
    -0.001023717857879348, -0.00062088751787392656, -0.0002214106920760022, 
    0.00017043042351921512, 0.00055037990185785113, 0.0009142889470896352, 
    0.0012581918787874069, 0.0015783856124696335, 0.0018715153365192901, 
    0.0021346521343863995, 0.0023653585171984452, 0.0025617427931373901, 
    0.0027224930118394828, 0.0028468823636303197, 0.0029347514246667733, 
    0.0029864739258097781, 0.0030029077700659363, 0.0029853408908151599, 
    0.0029354294702614047, 0.0028551406860198676, 0.0027466946424476711, 
    0.0026125017162083037, 0.0024551081368456261, 0.0022771376745966037, 
    0.0020812345513101745, 0.0018700097712849844, 0.0016459950396812233, 
    0.0014115954187526279, 0.001169057196080722, 0.00092043850917555468, 
    0.00066759407220485752, 0.00041216851792983333, 0.00015559225321187052, 
    -0.00010090985288170252, -0.00035631154237464747, 
    -0.00060976213694311648, -0.00086057283732310049, -0.0011081887415335665, 
    -0.0013521654101922185, -0.0015921449479204864, -0.0018278331615579956, 
    -0.0020589836902251209, -0.0022853809562089523, -0.0025068370827240087, 
    -0.0027231881665854404, -0.0029342978029565634, -0.0031400675269688083, 
    -0.0033404399342802787, -0.0035354077763583578, -0.0037250163044607733, 
    -0.0039093604567260144, -0.0040885709763933522, -0.0042628008512322554, 
    -0.0044321988753559822, -0.0045968844100461696, -0.0047569124650955899, 
    -0.0049122428424702288, -0.0050627075627335677, -0.0052079821949810121, 
    -0.00534756157101082, -0.005480754521956779, -0.0056066817119468371, 
    -0.0057242989957366408, -0.0058324263957890291, -0.0059297886919101482, 
    -0.0060150612537209361, -0.0060869168588933735, -0.0061440712380814366, 
    -0.0061853307968805565, -0.0062096351599627937, -0.0062161020374132143, 
    -0.006204071919647689, -0.0061731466822192013, -0.0061232304866109541, 
    -0.0060545597484023559, -0.0059677259139542423, -0.0058636836010670362, 
    -0.0057437389174063349, -0.0056095221289125703, -0.0054629501340779296, 
    -0.0053061699656181882, -0.0051415049376063561, -0.0049713924949661295, 
    -0.0047983237890354405, -0.0046247883434491835, -0.0044532139714265574, 
    -0.0042859149342387671, -0.0041250316882525005, -0.0039724777262800685, 
    -0.0038298968486590586, -0.0036986245719702214, -0.0035796702206426418, 
    -0.0034737131240577504, -0.0033811128833172092, -0.0033019352891219115, 
    -0.0032359833625171513, -0.0031828344255047801, -0.0031418746077291359, 
    -0.003112323473112463, -0.003093260211339894, -0.0030836324245039951, 
    -0.0030822635262980833, -0.0030878542710698368, -0.0030989865597402908, 
    -0.0031141365395966924, -0.0031317023723623372, -0.0031500463021206272, 
    -0.0031675494239375057, -0.0031826746386977773, -0.003194023132588414, 
    -0.0032003838800926656, -0.003200760807068203, -0.003194384902207921, 
    -0.0031807116400377989, -0.0031594205104211273, -0.0031304101901548191, 
    -0.0030937946897335476, -0.0030499032872327021, -0.0029992597009027623, 
    -0.0029425586263951841, -0.0028806241716175744, -0.0028143663618792167, 
    -0.0027447312570605129, -0.002672654052663515, -0.0025990216863357508, 
    -0.0025246463817380138, -0.0024502500494261547, -0.0023764615449680523, 
    -0.0023038226095710864, -0.0022328004005884223, -0.0021637962854462209, 
    -0.002097157731606319, -0.0020331867822393273, -0.0019721377068072639, 
    -0.0019142177267011994, -0.0018595863480638129, -0.0018083527312529198, 
    -0.0017605766055806898, -0.0017162762167216615, -0.0016754452813838498, 
    -0.0016380754620442428, -0.001604185701941264, -0.0015738500172326423, 
    -0.0015472185118724619, -0.0015245296519812426, -0.0015061103607512123, 
    -0.00149236359597778, -0.0014837446777163836, -0.0014807325408149666, 
    -0.0014837956659450883, -0.0014933614319241775, -0.0015097897508374836, 
    -0.0015333448459753003, -0.001564180354394648, -0.0016023163298482408, 
    -0.001647628776837074, -0.0016998403898019203, -0.0017585166974224253, 
    -0.0018230675804698517, -0.0018927569894662552, -0.001966716290018398, 
    -0.0020439635419918453, -0.0021234283720685332, -0.0022039758750983505, 
    -0.0022844313856678548, -0.0023636010939857535, -0.0024402851220732607, 
    -0.0025132868774818762, -0.0025814196528019511, -0.0026435100251269964, 
    -0.0026984045629112386, -0.0027449795541439289, -0.0027821596045182291, 
    -0.0028089412128225514, -0.0028244227524790028, -0.002827836231365143, 
    -0.0028185710307111278, -0.0027962042249858954, -0.0027605152090398976, 
    -0.0027114901587614341, -0.0026493316480192021, -0.0025744470650019623, 
    -0.0024874531782041729, -0.0023891701030346012, -0.0022806211824240958, 
    -0.0021630337224173607, -0.0020378392004766241, -0.0019066712958899293, 
    -0.0017713590375558965, -0.0016339132613432418, -0.0014965042404638056, 
    -0.0013614297466604543, -0.001231061401076556, -0.0011077901671998913, 
    -0.00099394753399070085, -0.00089171740325280332, 
    -0.00080305829950506923, -0.00072962438151895847, -0.0006727093391679232, 
    -0.00063320436498998491, -0.00061157863591235261, -0.00060787381235361427, 
    -0.00062171335154745377, -0.00065232687317184391, 
    -0.00069858595735387634, -0.0007590479508630709, -0.00083201660199558531, 
    -0.00091559955095585691, -0.0010077683053426227, -0.0011064071497404549, 
    -0.0012093499789583861, -0.0013144103263312676, -0.0014193945720493335, 
    -0.0015221220544159098, -0.0016204439411687942, -0.0017122854284309028, 
    -0.0017956898455250725, -0.0018688749019288994, -0.0019302841298292611, 
    -0.001978626832283763, -0.0020129135400806879, -0.002032480063789993, 
    -0.00203700104667121, -0.0020265124172771654, -0.0020014183623279038, 
    -0.0019625022649246283, -0.001910924716546493, -0.0018482120822403618, 
    -0.0017762278903479651, -0.0016971261009239554, -0.0016132897447802249, 
    -0.0015272597106665653, -0.0014416548772734784, -0.0013590885237427699, 
    -0.0012820956578665037, -0.0012130567934645511, -0.0011541391362568506, 
    -0.0011072466501977729, -0.0010739816662111296, -0.0010556189156340589, 
    -0.0010530952878991938, -0.0010670051283388413, -0.0010976183588988497, 
    -0.0011448922453102005, -0.0012085002309566992, -0.0012878489083229451, 
    -0.0013820996664598228, -0.0014901727902315648, -0.0016107493678393298, 
    -0.0017422645242860439, -0.0018828974232235601, -0.0020305716524721073, 
    -0.0021829635287203605, -0.0023375282765554666, -0.0024915501870353771, 
    -0.0026422046319447032, -0.0027866296237040399, -0.0029220092550541373, 
    -0.0030456548273925989, -0.0031550768580486934, -0.0032480565657784558, 
    -0.0033227008724415171, -0.0033774897444984386, -0.0034113103137093357, 
    -0.003423482444515822, -0.0034137625889278868, -0.003382336076912637, 
    -0.0033297743367487896, -0.0032569867698558795, -0.0031651471539483013, 
    -0.0030556088960005641, -0.002929819741998436, -0.0027892310031705468, 
    -0.0026352205857259623, -0.002469016957717592, -0.0022916450772078887, 
    -0.0021038873984721451, -0.001906270469114895, -0.0016990820878332116, 
    -0.0014824057229860708, -0.0012561897246162982, -0.0010203235704884126, 
    -0.00077472516615808684, -0.00051942299428167573, 
    -0.00025462483321963089, 1.9231509120698344e-05, 0.00030144814878224824, 
    0.00059105619726375997, 0.00088681698762928891, 0.0011872322166478079, 
    0.0014905677292526758, 0.0017948759267071258, 0.0020980285630402429, 
    0.0023977463622042276, 0.0026916258160032719, 0.0029771669481773104, 
    0.0032517984224969807, 0.0035129093292095371, 0.0037578763671433603, 
    0.0039841069813886017, 0.0041890829571799371, 0.0043704064923250352, 
    0.0045258502881558279, 0.0046534123270580352, 0.0047513692063568432, 
    0.0048183307648428427, 0.0048532925280434114, 0.0048556839930067371, 
    0.0048254038447590932, 0.004762842564869944, 0.0046688908922679177, 
    0.0045449321524141393, 0.0043928134007883406, 0.0042148064331800064, 
    0.0040135471187720626, 0.0037919717896612508, 0.0035532350162402644, 
    0.0033006252326061567, 0.0030374768609298781, 0.002767092884255219, 
    0.0024926837288070549, 0.0022173203512172628, 0.0019439172203594393, 
    0.0016752348377767356, 0.0014138967112930399, 0.0011624113632783999, 
    0.00092319253136385231, 0.00069856746028165424, 0.00049077379548353452, 
    0.00030193932620316527, 0.00013405717568163908, -1.104310712851013e-05, 
    -0.0001317249538453531, -0.00022657113485806014, -0.00029441068930445493, 
    -0.00033433335377331292, -0.00034571214783052432, 
    -0.00032821522428017259, -0.00028181637766248521, 
    -0.00020680123026386001, -0.00010377360476507524, 2.6337678670283087e-05, 
    0.0001822819257287701, 0.00036248405696273151, 0.00056505141329252727, 
    0.00078777494919281287, 0.0010281392706939416, 0.0012833356548673507, 
    0.0015502637769260884, 0.0018255580043959338, 0.0021056098781010802, 
    0.0023865977756128824, 0.0026645411643071637, 0.0029353548383227097, 
    0.0031949184091414427, 0.0034391613992149211, 0.0036641546471362571, 
    0.0038662040525307109, 0.0040419443498751727, 0.0041884277622446309, 
    0.0043031940802822312, 0.0043843306070461691, 0.0044305106830262106, 
    0.0044410179914551916, 0.0044157521184164349, 0.0043552232376257924, 
    0.0042605338008305056, 0.004133344471482169, 0.0039758307201381909, 
    0.0037906194428001185, 0.0035807216553523547, 0.0033494546621946151, 
    0.003100354825234733, 0.0028370880084282895, 0.0025633630724509996, 
    0.0022828436562859714, 0.0019990773061488408, 0.0017154210822905456, 
    0.0014349908733669215, 0.0011606201498296791, 0.00089483454298604941, 
    0.00063984902486911854, 0.00039756786663603473, 0.00016960214715073036, 
    -4.270384594263622e-05, -0.00023825031066106338, -0.00041615143905332947, 
    -0.00057571008576005769, -0.00071640383886283586, 
    -0.00083786765157313188, -0.00093989234502070938, -0.0010224233843350828, 
    -0.0010855699421759531, -0.0011296127506326701, -0.001155009709208239, 
    -0.0011624012319522972, -0.0011526062356121203, -0.0011266144539239396, 
    -0.0010855691096228746, -0.0010307452885337724, -0.00096352305014840267, 
    -0.00088535144842227624, -0.00079771402977511221, 
    -0.00070208398939986558, -0.00059987916148704823, 
    -0.00049241022924856814, -0.00038083851008210941, 
    -0.00026613807510840573, -0.0001490705646978428, -3.0176645983763335e-05, 
    9.0219667478599435e-05, 0.00021198734683381399, 0.00033516552299248667, 
    0.00045992186094637562, 0.00058653134705348355, 0.00071532703611956348, 
    0.00084667217345069643, 0.00098091383989814575, 0.0011183363512592718, 
    0.0012591124353070751, 0.0014032543667633097, 0.0015505740621212401, 
    0.0017006534822684577, 0.0018528251660545904, 0.0020061764265802344, 
    0.0021595594607487605, 0.0023116206132797463, 0.002460830848032378, 
    0.0026055252389208922, 0.0027439387524438009, 0.0028742412601402366, 
    0.0029945621797293166, 0.0031030251264886474, 0.0031977743712807184, 
    0.0032770059700726268, 0.0033390045751348833, 0.003382186926686381, 
    0.003405143074469456, 0.0034066919876711435, 0.0033859202363848285, 
    0.0033422296104464052, 0.0032753736185697074, 0.003185484742263418, 
    0.0030730951300907963, 0.0029391410609015921, 0.0027849610899091009, 
    0.0026122769271132418, 0.0024231735393551784, 0.0022200658574750153, 
    0.0020056524772852436, 0.0017828638445348891, 0.0015548108594277779, 
    0.0013247175897556547, 0.0010958426017487265, 0.0008714064767506494, 
    0.00065449796403934876, 0.00044797797178240591, 0.00025437867924535558, 
    7.5802563670205431e-05, -8.614416822932093e-05, -0.00023040557877703871, 
    -0.00035647880305450958, -0.00046439692875521445, 
    -0.00055468061465681589, -0.0006282911994556149, -0.00068658085923499154, 
    -0.00073124509280410018, -0.00076428918317848283, 
    -0.00078798259818141066, -0.00080479847870135971, 
    -0.00081733561339740934, -0.00082821770531906196, 
    -0.00083998296230019967, -0.00085498064522355653, 
    -0.00087527342769667276, -0.0009025710077222713, -0.00093818482242791635, 
    -0.00098301041972071574, -0.001037528126672662, -0.001101833430860152, 
    -0.0011756611733842258, -0.001258426375287749, -0.0013492625932485926, 
    -0.0014470580323380313, -0.0015505111116339912, -0.0016581736727248695, 
    -0.0017685102579417622, -0.0018799637903758226, -0.0019910080548115462, 
    -0.0021002093571320947, -0.0022062604661899775, -0.0023080126721006346, 
    -0.0024044833478977694, -0.0024948569425843111, -0.0025784704628394168, 
    -0.0026548006825379356, -0.0027234468457603056, -0.0027841162596980427, 
    -0.0028366179019988658, -0.002880861599747125, -0.0029168642713054112, 
    -0.0029447527184105499, -0.002964778692433878, -0.0029773369857270318, 
    -0.0029829791805616899, -0.0029824377387523927, -0.0029766433737211436, 
    -0.0029667467652911093, -0.0029541218226404819, -0.0029403641909112564, 
    -0.0029272666214824467, -0.0029167785037006785, -0.0029109569737794652, 
    -0.0029119059582989959, -0.002921730343347632, -0.0029424744988278328, 
    -0.0029760726093907394, -0.0030242955915474592, -0.0030887155000102165, 
    -0.0031706548911053967, -0.0032711582939977469, -0.0033909459621446411, 
    -0.003530385737112608, -0.0036894579226515972, -0.0038677304219834853, 
    -0.004064357005712684, -0.0042780948873627081, -0.0045073384874584638, 
    -0.00475017236498708, -0.0050044305695893417, -0.0052677550521505545, 
    -0.0055376476152911407, -0.0058115061704013459, -0.0060866512479669579, 
    -0.0063603542668783679, -0.006629857034896533, -0.0068924091297675209, 
    -0.007145305705095477, -0.0073859416530451874, -0.0076118660994109284, 
    -0.0078208533506448526, -0.0080109609328116779, -0.0081805927989486247, 
    -0.0083285639693974709, -0.008454149429735271, -0.0085571429900657119, 
    -0.0086378850211710212, -0.0086972796657011544, -0.0087367803243083141, 
    -0.0087583394962064132, -0.0087643271203353412, -0.0087574100646849763, 
    -0.0087404182870624587, -0.0087161930066998756, -0.0086874497205854505, 
    -0.0086566581084839365, -0.0086259323962533455, -0.0085969792363066923, 
    -0.0085710543328102479, -0.0085489634794399232, -0.0085310802573192821, 
    -0.008517387203255896, -0.008507535294956417, -0.0085009090696298705, 
    -0.0084967093479285504, -0.0084940393478102148, -0.008491993227528612, 
    -0.0084897415081180583, -0.0084866083839042535, -0.0084821371544694327, 
    -0.0084761288319742875, -0.0084686637407868966, -0.0084600964128194595, 
    -0.0084510136626136743, -0.0084421807442622964, -0.0084344685945029526, 
    -0.0084287799141515834, -0.008425991112083888, -0.0084269009177604191, 
    -0.0084321732428379349, -0.0084422786223070281, -0.0084574060716801347, 
    -0.0084773681961400459, -0.0085015144458307282, -0.0085286773519908151, 
    -0.0085571629937999539, -0.00858479675031186, -0.0086090263957588446, 
    -0.008627056125618442, -0.0086360063948420288, -0.0086330711588598272, 
    -0.0086156510870980148, -0.0085814666860563622, -0.0085286215511725782, 
    -0.0084556463248347986, -0.0083614921101323059, -0.0082455125061700121, 
    -0.0081074131568069883, -0.0079471971331658859, -0.0077651178223727794, 
    -0.0075616154893234557, -0.0073372826741330442, -0.0070928334236615414, 
    -0.0068291010809962182, -0.006547037070716008, -0.0062477289554833349, 
    -0.0059324267843223148, -0.0056025640921235865, -0.0052597862770230319, 
    -0.0049059686737998841, -0.0045432235430476718, -0.004173908559064683, 
    -0.0038006079767781528, -0.0034261033824623749, -0.0030533131934217046, 
    -0.0026852335176890162, -0.0023248467857071506, -0.0019750387839092237, 
    -0.0016385331759603266, -0.0013178234657075503, -0.0010151240338508, 
    -0.00073234068935192846, -0.00047105319723553165, 
    -0.00023251097355707324, -1.7633821644973744e-05, 0.00017297835136538675, 
    0.00033902543588093265, 0.00048049954977376385, 0.00059766850361695888, 
    0.00069104865055286374, 0.00076138130648555904, 0.00080960138949901156, 
    0.00083680085777950743, 0.00084420385281404689, 0.0008331349811676233, 
    0.00080499943261064407, 0.00076126690712353799, 0.00070345702175801921, 
    0.00063313807768163933, 0.00055191289453594976, 0.00046140352915726584, 
    0.00036324309262590951, 0.00025904495420724441, 0.00015039785573066496, 
    3.8820551991276944e-05, -7.4253927088119553e-05, -0.00018750481925684564, 
    -0.00029973507258563176, -0.00040986018911628509, 
    -0.00051689028257261265, -0.00061989191429113381, 
    -0.00071796092771416191, -0.00081021594529006788, 
    -0.00089579723172914861, -0.00097389332336821402, -0.0010437844930655867, 
    -0.001104869375310559, -0.001156716505323006, -0.0011990966425681629, 
    -0.0012319888513584909, -0.0012555958988231621, -0.0012703089560259651, 
    -0.0012766723966252543, -0.0012753370529568278, -0.0012669909035953623, 
    -0.0012522987746136785, -0.0012318502221350634, -0.0012061319624465674, 
    -0.0011755105261596493, -0.0011402437391737268, -0.0011005017143711588, 
    -0.0010564064472065042, -0.0010080616710625347, -0.00095559253790390762, 
    -0.00089917888182018538, -0.00083907864562081185, 
    -0.00077564812492878518, -0.00070935093788172213, 
    -0.00064076237159871698, -0.00057056477224606806, -0.0004995226787539264, 
    -0.00042846422005333404, -0.00035823562606749113, 
    -0.00028967385478944745, -0.00022355952117150192, 
    -0.00016059979515704723, -0.00010140384347231168, 
    -4.6478387992045811e-05, 3.7764211181738782e-06, 4.9069426972634184e-05, 
    8.9235363751964173e-05, 0.00012425797621580799, 0.0001543132991801169, 
    0.0001798078594284009, 0.0002014123540217973, 0.00022009345002240013, 
    0.00023710906320566376, 0.00025397831219945815, 0.00027242542842297502, 
    0.00029429971185127501, 0.00032148858701252294, 0.00035583082654624813, 
    0.00039903287750182241, 0.00045260307083570784, 0.00051780305319522118, 
    0.0005955940362556136, 0.00068661449251107261, 0.00079114791168667078, 
    0.00090911203593270473, 0.0010400491394893384, 0.0011831373328945482, 
    0.0013371945262506159, 0.0015007153998783437, 0.0016719096868916608, 
    0.0018487625468949901, 0.0020290993596479515, 0.0022106525568186693, 
    0.0023911324735481584, 0.0025682850639929928, 0.0027399568294817303, 
    0.0029041316952408735, 0.0030589833301010137, 0.0032028991819557104, 
    0.0033345063039622899, 0.0034526819476199365, 0.0035565599487879488, 
    0.0036455278043179581, 0.0037192333788420105, 0.0037775795319747946, 
    0.0038207358024711898, 0.0038491178578957883, 0.0038633927083895109, 
    0.0038644357651097445, 0.0038532994324440685, 0.0038311672014847489, 
    0.0037993043672876208, 0.0037590124325679029, 0.0037115921079148195, 
    0.0036583131732088516, 0.0036003672142090964, 0.0035388324343963271, 
    0.0034746278535177145, 0.0034084559312009453, 0.0033407655316640195, 
    0.0032717223411447755, 0.0032012184090943092, 0.0031289007299075667, 
    0.0030542383424842696, 0.0029765863058828458, 0.002895265529006145, 
    0.0028095851228953318, 0.0027188463252236202, 0.0026223137511983095, 
    0.0025191684229010866, 0.002408475919833614, 0.0022891688778539599, 
    0.002160049425738675, 0.0020198024757893504, 0.0018670073064537313, 
    0.0017001816654271527, 0.0015178264041356608, 0.0013184947087066955, 
    0.001100864083579473, 0.00086381773281020207, 0.00060651817678625025, 
    0.00032846408578864566, 2.9514560735649288e-05, -0.00029010117114290987, 
    -0.00062981178873225386, -0.00098872870492222056, -0.0013656992216426263, 
    -0.0017593191163803622, -0.0021679556573052719, -0.0025897395599700822, 
    -0.0030225621859046774, -0.0034640562612227501, -0.0039115914409360176, 
    -0.0043622583208819451, -0.0048128684951614896, -0.0052599567167190631, 
    -0.0056998143159014076, -0.0061285067556077315, -0.0065419364862920864, 
    -0.0069358996683428599, -0.0073061623709721815, -0.007648551932587096, 
    -0.0079590556981256385, -0.008233929369322086, -0.0084698013667661685, 
    -0.0086637652313493324, -0.0088134639379733662, -0.0089171356967337728, 
    -0.0089736470001386664, -0.008982508118293285, -0.0089438629463665011, 
    -0.0088584872665425727, -0.0087277435590791316, -0.0085535405158315998, 
    -0.0083382698080989148, -0.0080847408875853888, -0.0077961030638675584, 
    -0.0074757640969392554, -0.0071273133022379618, -0.0067544755097308853, 
    -0.0063610766634951124, -0.0059510246140656335, -0.0055283082157801628, 
    -0.0050969848456153535, -0.0046611633316395642, -0.0042249661432482198, 
    -0.003792486169903405, -0.0033677131540643603, -0.002954474947137633, 
    -0.0025563577020777822, -0.0021766482110836946, -0.0018182743337489243, 
    -0.0014837581301572653, -0.001175210536463317, -0.00089433737323096462, 
    -0.00064249774698836115, -0.00042077024012884666, 
    -0.00023002139287265258, -7.0946930618795968e-05, 5.5921785584648218e-05, 
    0.00015026535458524871, 0.0002120540366416402, 0.00024164616967816763, 
    0.0002398750286227935, 0.00020809526514056157, 0.00014818565716492903, 
    6.2504614507032766e-05, -4.6199202940346632e-05, -0.00017489614268956837, 
    -0.00032038388117559103, -0.0004793629007904161, -0.00064849049064778981, 
    -0.00082438288237716702, -0.0010036123834890596, -0.001182675114523528, 
    -0.0013579612631445931, -0.0015257569138393706, -0.0016822402216778013, 
    -0.0018235317639682383, -0.0019457751354851954, -0.0020452256908565199, 
    -0.0021183802249759953, -0.0021621079221279976, -0.0021737930147056449, 
    -0.0021514385748049362, -0.0020937611736562014, -0.0020002280643437119, 
    -0.0018710512409361854, -0.0017071872280323107, -0.0015103063053275511, 
    -0.001282784894189735, -0.0010276765887863835, -0.00074868191703301621, 
    -0.0004500893737016113, -0.00013669025870165254, 0.00018631896063237577, 
    0.00051344551970504198, 0.00083902009630597752, 0.0011572960204554686, 
    0.0014625909324807742, 0.0017494030591953013, 0.0020125274812393427, 
    0.0022472044939478783, 0.0024492139625191525, 0.0026149726210268473, 
    0.0027416147474665065, 0.0028270121248708487, 0.00286979284197878, 
    0.00286932702186361, 0.0028256962379797274, 0.0027396638054999318, 
    0.0026126309470230723, 0.0024465941100229767, 0.0022441034351041774, 
    0.0020082318125838354, 0.0017424981044335199, 0.0014508203004498068, 
    0.0011374493918817838, 0.00080689129153045365, 0.00046384947670140644, 
    0.00011315469321695254, -0.00024029403008618197, -0.00059158780411618659, 
    -0.00093588587602770395, -0.0012684868215465405, -0.0015849184960731587, 
    -0.0018810415424646378, -0.0021531582308572405, -0.0023981395244637646, 
    -0.0026135452848050403, -0.00279775022844664, -0.0029500558655967879, 
    -0.0030707484273261006, -0.0031611156735744301, -0.0032234151848076513, 
    -0.0032607783613305156, -0.0032770848011628825, -0.003276778464980441, 
    -0.0032646885676114231, -0.0032458425726364423, -0.0032252703930260632, 
    -0.0032078502613327275, -0.0031981600445629746, -0.0032003923467768826, 
    -0.0032182495020155939, -0.0032549086980760331, -0.0033129725902317384, 
    -0.003394426545337705, -0.0035006262327778297, -0.0036322757020795858, 
    -0.0037894359137581463, -0.0039715034125158378, -0.0041772402597126676, 
    -0.0044048077512720179, -0.0046518121216389584, -0.0049153671585064626, 
    -0.005192191328795389, -0.0054787179033651172, -0.0057712268086856488, 
    -0.0060659747954527141, -0.0063593534162045906, -0.0066480163320918797, 
    -0.0069290077151845115, -0.0071998271699284079, -0.0074584754862384263, 
    -0.007703459075088106, -0.0079337409346052767, -0.008148717144894525, 
    -0.0083481627837765169, -0.0085321932265145211, -0.0087012231422277757, 
    -0.0088559314291755328, -0.0089972135232619464, -0.0091261366194104587, 
    -0.0092438761939934617, -0.0093516857985729458, -0.0094508202126613507, 
    -0.0095424791654560651, -0.0096277758911135769, -0.0097076596552281794, 
    -0.0097828853355127407, -0.0098539838727388449, -0.0099212415319163538, 
    -0.0099847178162467791, -0.010044257265925503, -0.010099510212846068, 
    -0.010149942484082986, -0.010194854667042428, -0.010233419847838005, 
    -0.010264701185089639, -0.010287667856747994, -0.010301236836050786, 
    -0.010304292037519034, -0.010295723365772103, -0.010274456860983001, 
    -0.010239519649814403, -0.010190109991384462, -0.010125665798676154, 
    -0.010045932899699688, -0.0099510090801053063, -0.0098413387870364081, 
    -0.0097176998408826758, -0.0095811343619709444, -0.0094329137421909851, 
    -0.0092744768583828251, -0.009107397990567638, -0.0089333628950562169, 
    -0.0087541325287457169, -0.0085715125389569796, -0.0083873204559413699, 
    -0.0082032852792731752, -0.0080209980520470105, -0.0078418336474053666, 
    -0.0076668802585797028, -0.0074968989263127402, -0.0073323205298596967, 
    -0.0071732359466060098, -0.0070194643179789908, -0.0068706162127588144, 
    -0.0067261619961945223, -0.0065855434556017015, -0.0064482239055622904, 
    -0.0063137317601380935, -0.0061816672965067775, -0.0060516578179310686, 
    -0.0059232830614727779, -0.0057960195395409557, -0.0056691257594196085, 
    -0.0055415927395665518, -0.0054120865300087435, -0.0052789611315688335, 
    -0.0051402820749646286, -0.0049939220162219296, -0.0048376544284886858, 
    -0.0046692906652113699, -0.0044867899416565667, -0.0042883941013927623, 
    -0.0040727381545086032, -0.0038389160287203784, -0.003586546291795108, 
    -0.0033157781763335577, -0.003027280769085153, -0.0027221708579516102, 
    -0.0024019412250145438, -0.0020683404296877273, -0.0017232622188862942, 
    -0.0013686375922103739, -0.0010063450569819253, -0.00063818451350251284, 
    -0.00026585662198897023, 0.00010899545574723271, 0.00048477164279491321, 
    0.0008598396424055085, 0.0012324971737363508, 0.0016009197785272688, 
    0.0019631542629891677, 0.0023171063724527893, 0.0026605394459447282, 
    0.0029911473312638948, 0.0033065910040120487, 0.0036046147999124162, 
    0.0038831128016063024, 0.0041402095896659842, 0.0043743762966525438, 
    0.0045845351239614703, 0.0047701362818392502, 0.0049312916254097934, 
    0.0050688551085946287, 0.0051845058506167089, 0.0052807486078933555, 
    0.0053607746620029113, 0.0054281503281822883, 0.005486267088143643, 
    0.0055377382349676568, 0.0055838634706973905, 0.0056243865232509732, 
    0.0056575040722934107, 0.005680160211666928, 0.0056884579149307146, 
    0.0056780882694164765, 0.0056447364020837682, 0.0055844624046600174, 
    0.0054939331343449522, 0.0053706513552879073, 0.0052129806994493065, 
    0.0050202275398543092, 0.0047925206118485915, 0.0045308239518684649, 
    0.0042368537342860535, 0.0039130492513123182, 0.0035625542194440071, 
    0.0031891484111080401, 0.0027971543723906548, 0.002391330427772342, 
    0.0019767345559792431, 0.0015585565480647006, 0.0011419475182863224, 
    0.00073183807759139008, 0.00033274332897678731, -5.1400338990831637e-05, 
    -0.00041737582421592321, -0.00076276215413891425, -0.0010859683121473493, 
    -0.001386169567486259, -0.001663201257578047, -0.0019173820652421427, 
    -0.0021493022899378381, -0.0023596604432669145, -0.0025490125251875421, 
    -0.0027176809297886463, -0.0028656444833719827, -0.0029924758095629064, 
    -0.0030973344688316625, -0.0031789850041478765, -0.0032357933859790237, 
    -0.0032658339396183958, -0.0032669268087327698, -0.0032367539142236774, 
    -0.0031729299088795854, -0.0030731056239201612, -0.0029350362592712054, 
    -0.0027567070010494563, -0.0025364225332530459, -0.002272902629278446, 
    -0.0019653644694350237, -0.0016135527600629508, -0.0012177536150921673, 
    -0.00077880567827110024, -0.00029807187362106764, 0.00022252622343480594, 
    0.00078054020374990392, 0.0013729660504111349, 0.0019962036331594504, 
    0.0026460726807692901, 0.0033177979773828066, 0.0040060200399383546, 
    0.0047049202283712893, 0.005408260607934352, 0.0061095393003801094, 
    0.00680220683246569, 0.007479878578326769, 0.0081365748106921529, 
    0.0087669373191306427, 0.0093664289791067466, 0.0099314309689100579, 
    0.010459224492544156, 0.010947899937815321, 0.011396207047454809, 
    0.011803318429280013, 0.012168629991635422, 0.012491588432104114, 
    0.012771414345792946, 0.013007040174120117, 0.013196973527134802, 
    0.013339362715274283, 0.01343226621463202, 0.013474040192269025, 
    0.013463742680910867, 0.013401676694639359, 0.013289705396493585, 
    0.013131498105815948, 0.012932673004200429, 0.012700671479952954, 
    0.012444573878911519, 0.012174708831955617, 0.011902227718452911, 
    0.011638565027240548, 0.011394847721679317, 0.011181386159504191, 
    0.0110071885077329, 0.010879603569270532, 0.010804111902386306, 
    0.010784279574135783, 0.01082182176457828, 0.010916775476296013, 
    0.011067643740239675, 0.011271590871914931, 0.011524628479170075, 
    0.011821636087375907, 0.012156612432981191, 0.012522663975815198, 
    0.012912008596067172, 0.013315892008538711, 0.013724408754747746, 
    0.014126359603567154, 0.014509121105093599, 0.014858818579521649, 
    0.015160500007313713, 0.015398527110460728, 0.015557174694585242, 
    0.015621206090229789, 0.015576538275629154, 0.015410859804739361, 
    0.015114179999694242, 0.014679145101203005, 0.014101220435741949, 
    0.013378671923606773, 0.012512312204852036, 0.011505328197825704, 
    0.010363061691482024, 0.0090928999479050737, 0.0077045368265881006, 
    0.0062101798969258128, 0.0046246257215769278, 0.0029652839521319336, 
    0.0012518151643929119, -0.00049455083392868692, -0.002251721096295678, 
    -0.0039979038795619135, -0.0057125210690470909, -0.0073772626071957623, 
    -0.0089768106985787938, -0.010499576324871897, -0.011937957979143819, 
    -0.013288362298382273, -0.014551231775038859, -0.015730603676008707, 
    -0.016833509349990772, -0.017869558278777134, -0.018849986476296866, 
    -0.019786959563661659, -0.02069273417104257, -0.021578683608656144, 
    -0.022454271724384252, -0.023326133150851601, -0.024197452107101881, 
    -0.025067303592007224, -0.025930493229823368, -0.026778049336715029, 
    -0.027597665300692222, -0.028374957788319392, -0.029094689421877588, 
    -0.029741605244659679, -0.030301521218900809, -0.030762419802497807, 
    -0.031114228759622407, -0.03134962338218257, -0.031464115596667737,
  // Fqt-total(5, 0-1999)
    0.99999999999999956, 0.99655969307961756, 0.98633011727300113, 
    0.96958005611644704, 0.94674127297620703, 0.91838606452204785, 
    0.88519866209941045, 0.84794285385980928, 0.80742825711919231, 
    0.76447754421198399, 0.71989656458451379, 0.6744487903446873, 
    0.62883499431616385, 0.58367854449124712, 0.53951621202029698, 
    0.49679406595674869, 0.4558677480777043, 0.4170063125938207, 
    0.38039870694455513, 0.34616208883660415, 0.31435116575646094, 
    0.28496792510605484, 0.25797122230764724, 0.23328582961811942, 
    0.21081071317181097, 0.19042634947177978, 0.17200103984817391, 
    0.15539620619224326, 0.14047070325049549, 0.1270842348157821, 
    0.1150999655712423, 0.10438644316892157, 0.094818952015654726, 
    0.086280396709910501, 0.078661821100374174, 0.071862638405755574, 
    0.065790649782942939, 0.06036190608209796, 0.055500448749847449, 
    0.051137987407695124, 0.047213506685231048, 0.043672855316004261, 
    0.040468292181324694, 0.037558029336939677, 0.03490574261743095, 
    0.032480077188805842, 0.030254148247585402, 0.028205037941536417, 
    0.026313304210643582, 0.024562503030507766, 0.022938731026417442, 
    0.021430207377596499, 0.020026892408862559, 0.018720157859066736, 
    0.017502513197471568, 0.016367385468237589, 0.015308961168563128, 
    0.014322080549029418, 0.013402169053852863, 0.012545215462306313, 
    0.011747748069149152, 0.011006827091701088, 0.010320018044674429, 
    0.0096853447728727643, 0.0091012158745012658, 0.0085663286232597214, 
    0.0080795341872184692, 0.0076396972593208556, 0.0072455231590630052, 
    0.006895396864164397, 0.0065872395140496804, 0.0063183954239705315, 
    0.0060855642943635734, 0.0058847886414017296, 0.005711503670776984, 
    0.0055606334117660368, 0.0054267429335086992, 0.0053042240232357785, 
    0.0051875049973234477, 0.0050712701376409612, 0.0049506605528346227, 
    0.0048214583622990343, 0.0046802257243841695, 0.0045243953589370299, 
    0.0043523083394079462, 0.0041631985064574002, 0.0039571324355116549, 
    0.0037349154006168536, 0.0034979695738351969, 0.0032481954719866179, 
    0.0029878476727828451, 0.0027194008142893871, 0.0024454360436664056, 
    0.0021685366320427146, 0.0018911893597859696, 0.0016157009307567062, 
    0.001344131838366921, 0.0010782418986954282, 0.00081945204649422169, 
    0.00056882835056525462, 0.00032708108730968618, 9.4569494790851664e-05, 
    -0.00012867717803972687, -0.00034293028774780499, 
    -0.00054872357558102445, -0.00074680852674383156, 
    -0.00093809895146174994, -0.0011236064455597018, -0.0013043662561569847, 
    -0.0014813476349775209, -0.0016553552577594972, -0.0018269268887228631, 
    -0.0019962278233304873, -0.0021629660552203171, -0.0023263227554586219, 
    -0.0024849263912705647, -0.0026368588666099689, -0.0027797182779500345, 
    -0.0029107112032105559, -0.0030267800103774131, -0.003124753440173956, 
    -0.0032015050575807022, -0.0032541159688007459, -0.0032800193955460494, 
    -0.0032771350020671464, -0.003243972164687834, -0.0031796934841787747, 
    -0.0030841511126130771, -0.0029578823799672979, -0.0028020732231348552, 
    -0.0026185035335164319, -0.0024094691726149107, -0.0021777029765305375, 
    -0.0019262869074421628, -0.0016585633646768055, -0.0013780537210612118, 
    -0.001088368406818165, -0.00079313019368474963, -0.00049590670865238358, 
    -0.00020014387401757767, 9.087884539532462e-05, 0.00037409159299106934, 
    0.00064666015328973384, 0.00090600645611269904, 0.0011498202820400968, 
    0.0013760660895951709, 0.0015829881365075473, 0.0017691050200920164, 
    0.0019332061054297327, 0.0020743416846706617, 0.0021918119638485367, 
    0.0022851480019993333, 0.0023541141518199594, 0.0023987104969545336, 
    0.0024191999279895306, 0.0024161425291106373, 0.0023904387168845742, 
    0.0023433660133107804, 0.0022765891817165414, 0.0021921459918546045, 
    0.002092409493088932, 0.0019800242322250824, 0.0018578379839111201, 
    0.0017288245280728748, 0.0015960091965843148, 0.0014623913833703406, 
    0.0013308715119254946, 0.0012041737667363016, 0.0010847819265923972, 
    0.00097487416471706294, 0.00087627717684805428, 0.00079043810899023532, 
    0.00071840369415972314, 0.00066081374994094995, 0.00061790014892446976, 
    0.00058948281195363508, 0.00057498100571889618, 0.00057342285913315662, 
    0.00058347073245928625, 0.00060345812222138543, 0.0006314363357396676, 
    0.00066524511934301417, 0.0007025858811604309, 0.00074112833731872652, 
    0.00077861462669991826, 0.000812984053936478, 0.00084248605219852061, 
    0.00086577460428914209, 0.00088198523978793328, 0.00089076841709934465, 
    0.00089228830757313263, 0.00088717811808938557, 0.00087646914907829317, 
    0.00086148891615260884, 0.0008437540752966353, 0.00082486280324993943, 
    0.00080638780992115238, 0.00078979515075730403, 0.00077635826795030072, 
    0.00076709618936021532, 0.00076272692477339114, 0.00076363770072963085, 
    0.00076987550110268501, 0.00078115680856675215, 0.00079689054566446529, 
    0.00081621755728373353, 0.00083806858450509306, 0.0008612180650134681, 
    0.0008843513252299013, 0.00090612975415794116, 0.00092525103405225828, 
    0.00094050291851009422, 0.00095081642205484371, 0.00095530505094852843, 
    0.00095329989806734955, 0.00094437794671983983, 0.00092837926992752522, 
    0.00090541591188812807, 0.00087585901693805284, 0.00084031786005864663, 
    0.00079959672409482931, 0.00075463148704926406, 0.00070641949080815758, 
    0.00065593681992544631, 0.00060405055525948527, 0.00055143482969033418, 
    0.00049849701725705796, 0.0004453126411373457, 0.00039158931547632022, 
    0.00033665538983249088, 0.00027947838210600813, 0.00021872130567242672, 
    0.00015282031252780647, 8.0088327996089988e-05, -1.176974413487079e-06, 
    -9.2573488371104648e-05, -0.00019549292322537204, 
    -0.00031102515623685357, -0.00043989044429898841, 
    -0.00058238637043862037, -0.00073835523318452909, 
    -0.00090717813009419293, -0.0010877901441408877, -0.0012787177652796072, 
    -0.0014781408808903971, -0.0016839647857634886, -0.0018939105520926185, 
    -0.0021056009812363079, -0.0023166424822977428, -0.0025246962651561387, 
    -0.0027275350939118237, -0.0029230943064090208, -0.0031095061051673849, 
    -0.0032851334553086042, -0.0034485941659910539, -0.0035987783883348204, 
    -0.0037348552167501595, -0.0038562686932856853, -0.0039627245057265474, 
    -0.0040541660497722121, -0.0041307404445570361, -0.0041927706154381624, 
    -0.0042407212938991223, -0.0042751832119055149, -0.0042968546576486362, 
    -0.0043065283943688462, -0.0043050692799310513, -0.0042933804428202001, 
    -0.0042723560634622413, -0.0042428139022346973, -0.0042054324054786743, 
    -0.004160677052489771, -0.0041087463779269483, -0.0040495300996822052, 
    -0.0039825947037587482, -0.0039071892901319698, -0.0038222869128651652, 
    -0.0037266454715049503, -0.0036188979794616674, -0.0034976534076658784, 
    -0.0033616161394958502, -0.0032097048849679343, -0.0030411660206352761, 
    -0.0028556754935920052, -0.0026534221429022897, -0.0024351645671498129, 
    -0.002202260607607661, -0.0019566605857154738, -0.0017008794300908711, 
    -0.0014379318807053343, -0.0011712546852319877, -0.00090460467099963751, 
    -0.00064194214151145376, -0.00038730529649920871, 
    -0.00014468541125760789, 8.2091243752839985e-05, 0.00028947534471433192, 
    0.00047428018980103117, 0.00063374833044876433, 0.00076559626782063514, 
    0.00086803892863342668, 0.00093979412940375917, 0.00098007340028795006, 
    0.00098856329403505176, 0.00096539910836620038, 0.00091113223999324429, 
    0.00082669382778381001, 0.00071336075145228236, 0.00057272411376746359, 
    0.00040665084696164973, 0.00021725670612904132, 6.8580923212739305e-06, 
    -0.00022207960649242738, -0.00046700360690381205, 
    -0.00072534170840763605, -0.00099456163336322984, -0.0012722197034677619, 
    -0.0015559920607647059, -0.0018436844717909251, -0.0021332246736916441, 
    -0.0024226441619637907, -0.0027100588056708677, -0.002993650583733241, 
    -0.0032716680280656424, -0.0035424427220568967, -0.0038044072644171801, 
    -0.0040561326554066001, -0.004296339655340215, -0.0045239153710708883, 
    -0.0047378884898218532, -0.0049373890708342087, -0.0051215787397171217, 
    -0.0052895677237284281, -0.0054403391597588778, -0.0055726800607456377, 
    -0.0056851546474375961, -0.0057761112312108096, -0.0058437404230161786, 
    -0.0058861672676840263, -0.0059015730505046337, -0.0058883291202064631, 
    -0.005845127463444723, -0.0057710958468503559, -0.0056658886505648407, 
    -0.0055297509387296226, -0.0053635396626330401, -0.0051687292815589675, 
    -0.0049473696219236082, -0.0047020311530818707, -0.0044357148403049934, 
    -0.0041517545138629892, -0.0038536972297148341, -0.0035451861718517495, 
    -0.0032298344318536843, -0.0029111246663837539, -0.0025923157873865665, 
    -0.0022763752766834272, -0.0019659229369984425, -0.0016631843848724781, 
    -0.0013699577695056445, -0.0010875826026711744, -0.00081692239376317895, 
    -0.0005583606855512509, -0.00031181533506150053, -7.6771214095664104e-05, 
    0.00014766274475016601, 0.00036268759946619553, 0.00056973360514296005, 
    0.00077038042355743552, 0.00096627963160848904, 0.0011590908777779582, 
    0.0013504308947389701, 0.0015418384136697489, 0.0017347531458097071, 
    0.00193050768378085, 0.0021303336423499027, 0.002335362084086821, 
    0.0025466319349090336, 0.0027650757988243557, 0.0029914970041647593, 
    0.0032265285930654425, 0.0034705730430265366, 0.0037237380628485114, 
    0.0039857643508932651, 0.0042559645001013745, 0.0045331776880019247, 
    0.0048157577491298904, 0.0051015875383587719, 0.0053881348975466968, 
    0.0056725298892981932, 0.0059516692186851131, 0.006222325534819449, 
    0.006481266420287379, 0.006725370388461732, 0.0069517364733079562, 
    0.0071577874044119515, 0.0073413506549036799, 0.007500724939567543, 
    0.007634716645834809, 0.0077426491772202627, 0.0078243456338191655, 
    0.0078800822593364708, 0.0079105328371221091, 0.0079166930561560163, 
    0.0078998069497163027, 0.0078612925654434566, 0.0078026741686643333, 
    0.0077255249528168915, 0.0076314113254306168, 0.0075218588116077794, 
    0.0073983231786065922, 0.0072621794705438041, 0.0071147246306329818, 
    0.0069571969552700225, 0.0067908054354034117, 0.0066167771397339856, 
    0.0064363910670209622, 0.0062510124774842737, 0.0060620991004413901, 
    0.0058711901265807035, 0.0056798610361212688, 0.0054896630046470827, 
    0.005302040698726398, 0.0051182494777921011, 0.0049392727279021003, 
    0.0047657555139393338, 0.0045979564942227455, 0.0044357284696153665, 
    0.0042785185725255515, 0.0041253978777804484, 0.0039750953630597434, 
    0.0038260475330149798, 0.0036764451149879172, 0.0035242821090188878, 
    0.003367408917229447, 0.0032035977204340682, 0.0030306228709790126, 
    0.0028463698736722136, 0.0026489655981453857, 0.0024369204263149213, 
    0.0022092762556467512, 0.0019657299361249465, 0.0017067197502268275, 
    0.0014334550304185196, 0.0011478873806462784, 0.00085262206887316795, 
    0.00055077897296736675, 0.00024581709668567098, -5.8658424415996339e-05, 
    -0.00035908925188453069, -0.00065213256029039875, 
    -0.00093479822554071309, -0.0012045530353883979, -0.0014594014760152107, 
    -0.0016979467875728009, -0.0019194352384980067, -0.0021237727045104126, 
    -0.0023114993137102378, -0.0024837112380593929, -0.0026419368552149107, 
    -0.0027879689100419932, -0.0029236864247330521, -0.0030508559567221016, 
    -0.0031709639292269959, -0.0032850658021617864, -0.0033936698068155946, 
    -0.00349666387326908, -0.0035932858499876604, -0.0036821415960252911, 
    -0.0037612691971504308, -0.0038282518671318207, -0.0038803672577784262, 
    -0.0039147721539856501, -0.0039286982419568812, -0.0039196471942485574, 
    -0.0038855789367271509, -0.0038250659660275465, -0.0037374168314013678, 
    -0.003622754830393992, -0.0034820524051254603, -0.0033171160020616383, 
    -0.003130533867259038, -0.0029255913178336157, -0.0027061656732243395, 
    -0.0024766013607282924, -0.0022415903244859133, -0.0020060457182587399, 
    -0.0017749876272434319, -0.00155343558777289, -0.0013463018197508133, 
    -0.0011582939768620135, -0.00099381947175282144, -0.00085687612881411987, 
    -0.00075095829642920532, -0.00067895497140428411, 
    -0.00064305514726041319, -0.00064466571792434497, -0.0006843317565121609, 
    -0.00076167333887562064, -0.00087533841896033043, -0.0010229948545711206, 
    -0.0012013449778212736, -0.0014061968730363225, -0.0016325656303324912, 
    -0.0018748198646388271, -0.002126844167053311, -0.0023822219980375705, 
    -0.0026344136917967578, -0.0028769463381634508, -0.0031035930084120666, 
    -0.0033085511741048038, -0.0034866164768750092, -0.0036333410078331265, 
    -0.0037451761810348592, -0.0038195809422089883, -0.0038550958205409843, 
    -0.0038513620780222975, -0.0038090975723997617, -0.003730021213705892, 
    -0.0036167419391204872, -0.0034726244441819513, -0.0033016370214343604, 
    -0.0031082049045321114, -0.0028970723080559502, -0.0026731792262425524, 
    -0.0024415537971571818, -0.0022072196539805466, -0.0019751216612497197, 
    -0.0017500469049622812, -0.0015365544387396419, -0.0013388935092705997, 
    -0.0011609274736058893, -0.0010060522865351855, -0.00087712454140101285, 
    -0.00077638165470131099, -0.00070537612269980416, 
    -0.00066491090986144747, -0.00065500324218243722, 
    -0.00067486604941802283, -0.00072292070906965526, 
    -0.00079683935102926884, -0.0008936068916510229, -0.0010096132821992873, 
    -0.00114076151301885, -0.0012825909023800341, -0.0014304165178582985, 
    -0.0015794686667611336, -0.001725040905059627, -0.0018626286526793273, 
    -0.0019880590893055212, -0.002097598857612164, -0.002188034501863622, 
    -0.0022567225359534275, -0.0023016066288080186, -0.0023211982059934311, 
    -0.0023145304297078821, -0.0022810851998908113, -0.0022207216097874429, 
    -0.0021335949666744483, -0.0020200959809016676, -0.0018807990653644108, 
    -0.0017164297557712878, -0.0015278476953765325, -0.0013160364057452987, 
    -0.0010821051137868518, -0.00082729664278739345, -0.00055300247855381022, 
    -0.00026077839017758141, 4.7637015289930073e-05, 0.00037029757886255333, 
    0.00070503295638476898, 0.0010494310462144558, 0.0014008263389924112, 
    0.0017562984338023824, 0.0021126752929947808, 0.0024665453351589667, 
    0.0028142813135593075, 0.0031520686854679138, 0.0034759543098623036, 
    0.0037819004974336133, 0.004065861981798714, 0.0043238655321288441, 
    0.0045521044065892115, 0.0047470412857614427, 0.0049055080903788809, 
    0.0050248101497244674, 0.0051028251399210601, 0.0051380831853974143, 
    0.0051298426086657861, 0.0050781376149482685, 0.004983801585065898, 
    0.0048484729430311275, 0.0046745647955055182, 0.004465217237828144, 
    0.0042242145308784129, 0.0039558802552833155, 0.0036649469975599154, 
    0.0033564010912160809, 0.0030353184827002569, 0.0027066941967872626, 
    0.0023752904008374266, 0.0020454971643502798, 0.0017212323788189064, 
    0.0014058649064574204, 0.0011021890166799653, 0.00081242282059482986, 
    0.00053824398154965513, 0.00028084700872179941, 4.1019221126853896e-05, 
    -0.00018077736074641692, -0.00038432596001014384, 
    -0.00056957808570776429, -0.00073659022588016382, 
    -0.00088547047903083178, -0.0010163448284188018, -0.0011293351331125496, 
    -0.0012245556874483283, -0.0013021191614027948, -0.0013621593835834414, 
    -0.0014048600485466337, -0.0014304907041915904, -0.0014394263490516855, 
    -0.0014321769111146669, -0.0014093994151944391, -0.001371898583950281, 
    -0.0013206203467593836, -0.0012566444786650378, -0.0011811686011993366, 
    -0.001095492980282552, -0.0010010024275339748, -0.00089914729355001903, 
    -0.00079142511973465763, -0.00067936734301534297, -0.0005645305206554924, 
    -0.0004484788794171753, -0.00033278233084451129, -0.00021899822019086286, 
    -0.00010865589404133896, -3.2351652999925104e-06, 9.5865331338365048e-05, 
    0.00018736969729930841, 0.00027016945604067268, 0.00034338068602992249, 
    0.00040639660241818842, 0.00045894671430389919, 0.00050114686361315587, 
    0.0005335553727919025, 0.0005571983396064987, 0.00057358816887269359, 
    0.00058470523541824461, 0.00059295376518373236, 0.00060108541033918701, 
    0.00061209312914859793, 0.00062908728907145098, 0.00065515986580709376, 
    0.00069324060156821866, 0.00074596160015253212, 0.00081553261702395168, 
    0.00090363224031394694, 0.0010113200688845597, 0.0011389726404519853, 
    0.0012862487580065796, 0.0014520832255165241, 0.0016347155397948003, 
    0.0018317504964883225, 0.0020402537342668588, 0.002256882182833288, 
    0.0024780317004427584, 0.0027000005661782884, 0.0029191536980134425, 
    0.0031320665149739964, 0.0033356383103870435, 0.0035271726667369034, 
    0.0037044101138003121, 0.0038655244260773882, 0.0040090770022706765, 
    0.004133943767567155, 0.0042392242610263921, 0.0043241363339758263, 
    0.0043879172840539772, 0.0044297349647209735, 0.0044486241631463306, 
    0.0044434561947142501, 0.0044129565848772118, 0.0043557642338776514, 
    0.004270521069799681, 0.0041559913823243262, 0.0040111910010025512, 
    0.0038355259549007546, 0.0036289279354672589, 0.0033919812388718065, 
    0.0031260313223239341, 0.0028332464192061882, 0.0025166465255988578, 
    0.0021800729218191444, 0.0018281144280417037, 0.0014659903987616753, 
    0.0010993918622795213, 0.00073430038775328999, 0.00037677928222307964, 
    3.2775045300151898e-05, -0.00029207455461134597, -0.00059259124981440577, 
    -0.00086417515930948781, -0.0011028829330491175, -0.0013054746771204012, 
    -0.0014694242366916192, -0.0015929117897533933, -0.0016747978665846569, 
    -0.0017145979296309317, -0.0017124548247709132, -0.0016691054976812876, 
    -0.0015858639173181297, -0.0014645977428925452, -0.0013077053098294459, 
    -0.0011180861078654973, -0.00089909830753629046, -0.00065449410261253526, 
    -0.00038833392597315095, -0.00010488735404529319, 0.00019148755928198835, 
    0.00049646980600481121, 0.00080589980579898527, 0.001115894740103981, 
    0.0014229512325015551, 0.0017240187534454316, 0.0020165539096463898, 
    0.0022985443779652654, 0.0025685006848633674, 0.0028254226664872857, 
    0.0030687389021409983, 0.0032982319941039276, 0.0035139600111587883, 
    0.0037161769454917126, 0.0039052568047294733, 0.0040816277110167819, 
    0.0042457138924529682, 0.0043978769852660287, 0.0045383782361911951, 
    0.0046673382809263577, 0.0047847144477105672, 0.004890285725091076, 
    0.0049836497770385669, 0.0050642248945080058, 0.0051312494626070742, 
    0.0051837922193511297, 0.0052207586270516934, 0.0052409127437235007, 
    0.0052429190707944185, 0.0052253946674876654, 0.0051869837736022457, 
    0.005126439477858861, 0.0050427081616635262, 0.0049350142231071245, 
    0.0048029329545197699, 0.0046464481183402734, 0.004465993879662622, 
    0.0042624830963122438, 0.0040373244594389341, 0.003792417642198836, 
    0.0035301443973077204, 0.0032533290520380532, 0.0029651896457283103, 
    0.0026692680634258122, 0.0023693458636452084, 0.0020693474797279631, 
    0.0017732479424042407, 0.0014849841152369072, 0.0012083716199371426, 
    0.00094703339394485754, 0.00070434131560176438, 0.00048335314514513566, 
    0.00028676257293385675, 0.00011684619993198038, -2.4586114809143988e-05, 
    -0.00013623120877734234, -0.00021732844324967332, -0.0002676871081618888, 
    -0.0002877001776131327, -0.00027834890755129896, -0.00024120133643681577, 
    -0.00017838639872115591, -9.2565023120349242e-05, 1.3119520638282387e-05, 
    0.00013511530394975216, 0.00026955107154456973, 0.00041234483613781158, 
    0.00055932558540713179, 0.00070636283004618617, 0.00084949494729741196, 
    0.00098504730038563386, 0.0011097387068360657, 0.0012207717519339282, 
    0.0013159037784922646, 0.0013934985842527841, 0.0014525625733320959, 
    0.001492757719216908, 0.0015143990343580369, 0.0015184288138554609, 
    0.001506375464828675, 0.0014802912262534035, 0.0014426731330612018, 
    0.0013963645093743495, 0.0013444383159622259, 0.0012900701936581836, 
    0.0012364176752492535, 0.001186492223454288, 0.0011430562569746394, 
    0.0011085444115662036, 0.0010850151830917117, 0.0010741254881437539, 
    0.0010771299199374132, 0.0010948971711165357, 0.0011279353760424455, 
    0.001176411561666384, 0.0012401809379590993, 0.0013188108682692097, 
    0.0014116005625612338, 0.0015176075844282929, 0.0016356663029623352, 
    0.0017644149366149281, 0.0019023182879437542, 0.0020476837606406067, 
    0.0021986881834647602, 0.002353396955069231, 0.0025097874642115272, 
    0.0026657758080398013, 0.0028192496050492596, 0.0029681000701473332, 
    0.0031102603950868939, 0.003243744934488891, 0.0033666900436137262, 
    0.0034773965159153111, 0.0035743663696624762, 0.0036563416728625643, 
    0.0037223290593842886, 0.0037716242370507691, 0.0038038155338277761, 
    0.0038187831070200062, 0.0038166747567566594, 0.0037978896048815251, 
    0.0037630412080258591, 0.0037129267771856263, 0.0036484951308552098, 
    0.0035708133318348764, 0.0034810424337859028, 0.0033804027825300232, 
    0.0032701490606174759, 0.0031515418159656643, 0.0030258190297953241, 
    0.0028941668114880253, 0.0027576944730693599, 0.0026174066976326128, 
    0.0024741780028526973, 0.0023287332689097382, 0.0021816296344059341, 
    0.0020332463406266422, 0.001883795660420156, 0.0017333448213785723, 
    0.0015818619950333987, 0.0014292867694291453, 0.0012756108367356755, 
    0.0011209746544036199, 0.00096575425499826283, 0.00081064479746781586, 
    0.00065670392096030055, 0.00050536894052184494, 0.00035841971035934834, 
    0.00021789368271815687, 8.596162193572834e-05, -3.5222070019277657e-05, 
    -0.00014368353047330748, -0.00023777024476709735, 
    -0.00031626404927542111, -0.00037845126563211654, 
    -0.00042415531573687388, -0.0004537299037277009, -0.00046804213712387096, 
    -0.00046841575143064836, -0.00045657322352875881, 
    -0.00043455804735226933, -0.00040464850879337144, 
    -0.00036925638947351717, -0.0003308314046141219, -0.00029175751043320646, 
    -0.00025426613274038971, -0.00022036741789112417, 
    -0.00019179599606447987, -0.00016999614448588962, 
    -0.00015612318717622153, -0.00015106938383116465, -0.0001554986148028587, 
    -0.00016988802998581202, -0.0001945559494665241, -0.00022968661956440745, 
    -0.00027533830806317932, -0.00033143813002159612, 
    -0.00039777217696007665, -0.00047396341512413194, 
    -0.00055946555218715493, -0.00065355284360450717, 
    -0.00075532325529418913, -0.00086371149462923132, 
    -0.00097751195807019059, -0.001095402400931573, -0.0012159809855411658, 
    -0.0013378029487631522, -0.0014594222863502449, -0.0015794369404048077, 
    -0.0016965311607919692, -0.0018095157546662514, -0.0019173606921869049, 
    -0.0020192228266027795, -0.0021144585715598013, -0.0022026279570249211, 
    -0.0022834784375951279, -0.0023569196648025861, -0.0024229857629384879, 
    -0.0024817766232271706, -0.0025334161770325246, -0.0025780042923471331, 
    -0.0026155809774663615, -0.0026461192821239225, -0.0026695275448183672, 
    -0.0026856725962515005, -0.0026944100167473218, -0.0026956187496586857, 
    -0.0026892285076222373, -0.0026752422082160035, -0.0026537480437965207, 
    -0.0026249164298131236, -0.0025889808233833266, -0.0025462100795650209, 
    -0.0024968576855810844, -0.0024411066646251364, -0.0023790040719078366, 
    -0.0023104060908530647, -0.0022349411988742051, -0.0021520047178029082, 
    -0.0020608063613227049, -0.0019604490050762679, -0.0018500537849409006, 
    -0.0017289004572564441, -0.0015965579090837054, -0.0014529966248533741, 
    -0.0012986516114651086, -0.0011344618520814638, -0.00096186326445657987, 
    -0.00078275565577786181, -0.00059945045333212571, 
    -0.00041458873605857257, -0.00023104441448100848, 
    -5.1809368809794524e-05, 0.0001201168947963928, 0.00028184557138211363, 
    0.00043069119964703103, 0.00056425670299987572, 0.00068049046985767931, 
    0.00077772851794684242, 0.0008547309555691679, 0.00091070309620342989, 
    0.00094532266087562805, 0.00095875575553870749, 0.00095166425174574639, 
    0.0009251932122842177, 0.00088093395442480674, 0.00082087172219183003, 
    0.00074729862625343764, 0.00066272451606103956, 0.00056977289755959031, 
    0.00047107806535469306, 0.00036918724383195017, 0.00026647744029395531, 
    0.00016509501300062123, 6.6901157175222939e-05, -2.6545986091498005e-05, 
    -0.00011400197700187884, -0.00019451899832077747, 
    -0.00026743462773268732, -0.00033233561371552481, 
    -0.00038903621399940884, -0.00043755027320437116, 
    -0.00047807125427753273, -0.0005109446862510608, -0.00053664604596294135, 
    -0.00055575513747370972, -0.00056892840624506668, 
    -0.00057687884320039131, -0.00058036535604948797, 
    -0.00058018846364535869, -0.00057719767483983776, 
    -0.00057229635167743264, -0.00056644135991622735, 
    -0.00056062759052347372, -0.00055586236334338897, 
    -0.00055312355803921324, -0.00055331153980683618, -0.0005571955741098968, 
    -0.00056536224846167661, -0.00057816153131591151, 
    -0.00059567013339067412, -0.00061765485270454795, 
    -0.00064355235183216478, -0.00067246271170823561, 
    -0.00070315391124638194, -0.00073408419064171777, 
    -0.00076342865661444513, -0.00078913311976725581, 
    -0.00080896270175860423, -0.00082058276135311742, 
    -0.00082163843850330839, -0.00080984559978681918, 
    -0.00078307941306720176, -0.00073945794356886855, 
    -0.00067741939341888142, -0.00059579192163833913, 
    -0.00049385291368043136, -0.00037139050117993564, 
    -0.00022875852250366576, -6.6922448574442261e-05, 0.00011249481287410079, 
    0.00030720144317448469, 0.00051424195042174123, 0.00073004057064407664, 
    0.00095047860239824754, 0.0011710149500263479, 0.0013868319588025745, 
    0.0015930214671266614, 0.0017847847098973273, 0.0019576469631054291, 
    0.0021076708019782662, 0.0022316473734432908, 0.0023272549119705333, 
    0.0023931601191730222, 0.0024290628247610434, 0.0024356719200534604, 
    0.0024146152886119431, 0.002368303733869777, 0.0022997516057282818, 
    0.0022123755049810912, 0.002109793676982052, 0.0019956270552886337, 
    0.0018733282232595403, 0.0017460359885262411, 0.0016164715424133995, 
    0.0014868757914587437, 0.001358981246709999, 0.0012340355383685102, 
    0.0011128456442695287, 0.00099585587606894712, 0.00088322725656179567, 
    0.00077492169507825009, 0.00067076649795171756, 0.00057049732914968689, 
    0.00047377834271770356, 0.00038021281485373592, 0.00028934341786292223, 
    0.00020066143784412606, 0.00011363790118915283, 2.7760715192532975e-05, 
    -5.740682895502314e-05, -0.00014216914295624982, -0.00022664630795556589, 
    -0.00031074791798840144, -0.00039415597525669114, 
    -0.00047631921252427878, -0.00055645192573424286, -0.0006335350445809642, 
    -0.00070632584309338335, -0.00077337277158893622, -0.0008330310532841691, 
    -0.00088349296231616007, -0.0009228153665544269, -0.00094895523578115623, 
    -0.0009598170049796319, -0.00095329085806648481, -0.00092731300457432001, 
    -0.00087992546119754678, -0.00080934921965130941, 
    -0.00071406639213819905, -0.00059290323745080672, -0.0004451055947689021, 
    -0.00027041266962113912, -6.9099779530277768e-05, 0.00015799026365036299, 
    0.0004094436372951322, 0.00068329816537360114, 0.00097708790701963037, 
    0.0012879095253186326, 0.001612506054113371, 0.0019473724705353214, 
    0.002288855596646577, 0.002633257544954731, 0.0029769183166729403, 
    0.0033162771030310679, 0.0036479161926207507, 0.0039685929051324976, 
    0.004275273048186732, 0.0045651728135175365, 0.0048358183436975821, 
    0.0050851123197510947, 0.0053114040333900334, 0.0055135553420589557, 
    0.0056910013127647935, 0.0058437849749145921, 0.0059725815779346717, 
    0.0060786799012221872, 0.006163950569340328, 0.006230764370911618, 
    0.0062818955411504647, 0.0063203864360144909, 0.0063493944509126245, 
    0.0063720305588104032, 0.0063912036076035792, 0.0064094720202711843, 
    0.0064289306821521258, 0.0064511247864924275, 0.0064770087645260313, 
    0.0065069474059820534, 0.0065407549361006503, 0.0065777701014324303, 
    0.0066169539890082955, 0.0066570008052052659, 0.0066964372914027938, 
    0.0067337224302088192, 0.006767323471424321, 0.0067957666600475591, 
    0.0068176688945151944, 0.0068317576984897122, 0.0068368590754296658, 
    0.006831899551327715, 0.0068158835035293831, 0.0067878911070233224, 
    0.0067470762221113504, 0.0066926776820301747, 0.0066240436454621538, 
    0.0065406560280251861, 0.0064421537574878684, 0.0063283589560945508, 
    0.0061992729170150035, 0.0060550711878693542, 0.0058960763358431954, 
    0.0057227190997511234, 0.0055354925290887081, 0.0053349103081706366, 
    0.0051214658782448956, 0.0048956147880850941, 0.0046577643708599322, 
    0.0044082959930222378, 0.0041475938301557963, 0.0038760930451138109, 
    0.0035943357151046853, 0.0033030213619301865, 0.0030030558544362142, 
    0.0026955917731647087, 0.0023820590863128646, 0.0020641925735843591, 
    0.0017440444466184644, 0.001423984587687097, 0.0011066886182117942, 
    0.00079510162357732757, 0.00049238544815447427, 0.00020184443969547991, 
    -7.3156944253483525e-05, -0.00032930024128010558, 
    -0.00056341629009257189, -0.00077258183566708571, 
    -0.00095422968039165829, -0.0011062371028364828, -0.0012270167679032311, 
    -0.0013155915018564003, -0.0013716615496372879, -0.0013956426855209214, 
    -0.0013886863749638604, -0.001352666455000529, -0.0012901334269108597, 
    -0.0012042521748866681, -0.0010987137571696792, -0.00097763792492867657, 
    -0.00084547682937549955, -0.00070690250554074428, 
    -0.00056670964482129031, -0.00042971400450953439, 
    -0.00030064107126096917, -0.00018401761290664186, 
    -8.4049478230153321e-05, -4.4969964636899446e-06, 5.1449234184468782e-05, 
    8.130306329196194e-05, 8.3401957801210221e-05, 5.700314762547899e-05, 
    2.3600609320767723e-06, -7.9243009147898137e-05, -0.00018549179245941794, 
    -0.00031310120760831832, -0.00045790018262832779, 
    -0.00061495813258709937, -0.00077874957386420563, 
    -0.00094334610111660745, -0.0011026264865663655, -0.0012504998130866483, 
    -0.0013811417950449661, -0.001489215584961043, -0.0015700867451306306, 
    -0.0016200088722600503, -0.0016362822632607862, -0.0016173714447418729, 
    -0.0015629799686281089, -0.0014740722185770645, -0.0013528494019730787, 
    -0.0012026836113083049, -0.0010280053327766984, -0.00083416517007368104, 
    -0.00062726391178952103, -0.00041397101578008699, 
    -0.00020132129601011084, 3.5010305541050432e-06, 0.00019338024441515648, 
    0.00036148900469064012, 0.00050151093313906367, 0.0006078490054983207, 
    0.00067581977095973933, 0.00070179616818737806, 0.00068332862390031138, 
    0.0006192060363247844, 0.00050946395543308642, 0.00035534370648768952, 
    0.00015920652222277368, -7.5594590167530915e-05, -0.0003448743944789487, 
    -0.00064379052325969142, -0.00096702907462890549, -0.0013089871458932835, 
    -0.0016639395956032071, -0.0020261800300529023, -0.0023901314168392924, 
    -0.0027504220264096073, -0.0031019433314947858, -0.0034398875834398962, 
    -0.0037597760733943763, -0.0040575068677610711, -0.0043293975844665164, 
    -0.0045722355509654165, -0.0047833319582970078, -0.0049605632797051049, 
    -0.0051024034537670527, -0.0052079548076032368, -0.0052769632341420469, 
    -0.0053098225498867391, -0.0053075849459183434, -0.0052719476743531028, 
    -0.005205225911688479, -0.0051102910665214839, -0.0049904899425524014, 
    -0.0048495272058144481, -0.0046913385781667564, -0.0045199433700759241, 
    -0.0043393146465861097, -0.004153252820139364, -0.0039652829028929493, 
    -0.0037785703101112403, -0.00359586019694362, -0.0034194334507610035, 
    -0.0032510836367938777, -0.0030921187546697811, -0.0029433644957938482, 
    -0.0028051791958163749, -0.0026774801665671887, -0.0025597586287545845, 
    -0.0024510951280587384, -0.0023501795436377724, -0.0022553462051334498, 
    -0.0021646243584120175, -0.0020758058698128806, -0.0019865288004618283, 
    -0.0018943688928437568, -0.0017969338105318169, -0.001691957134149733, 
    -0.0015774017236748756, -0.0014515540524374663, -0.0013131328348781168, 
    -0.0011613773724121646, -0.00099612640205253532, -0.00081788232134892059, 
    -0.00062783950630924707, -0.00042788629241828917, 
    -0.00022057910090536058, -9.0737396875544404e-06, 0.00020297142337857209, 
    0.00041152406759770101, 0.00061233300613556803, 0.00080109607094389068, 
    0.0009736324052035749, 0.0011260465995711563, 0.0012548880691115006, 
    0.0013572924391923021, 0.0014311086109201987, 0.0014750067133062488, 
    0.0014885645174880216, 0.0014723199692039202, 0.0014277794240065847, 
    0.0013573826336200682, 0.0012644169924829001, 0.0011528874244901893, 
    0.001027343775232107, 0.0008926904295631495, 0.00075399221615859329, 
    0.00061627330856725397, 0.000484330419337269, 0.00036256752186325893, 
    0.00025486113398480247, 0.00016443504580484261, 9.3781906692770345e-05, 
    4.4591180653930204e-05, 1.7696983893737504e-05, 1.3030456843822729e-05, 
    2.9600210278072781e-05, 6.5462098613297735e-05, 0.00011775060002008919, 
    0.00018273570966379654, 0.00025595646200460076, 0.00033240432428200252, 
    0.00040674255211379287, 0.0004735580013849223, 0.00052762397271958973, 
    0.00056414822650546932, 0.00057899934752769799, 0.00056889006699740118, 
    0.00053150635315372182, 0.00046558887225857073, 0.00037095269828539573, 
    0.00024846057787104392, 9.9950024279717224e-05, -7.1862932778689084e-05, 
    -0.00026352221834123282, -0.00047099506011262466, 
    -0.00068986146938945238, -0.00091552154272563958, -0.0011434085792824244, 
    -0.0013691862127772135, -0.0015889338687306448, -0.0017992921171705988, 
    -0.0019975793666390145, -0.0021818480011237748, -0.00235091280416153, 
    -0.0025043250120416623, -0.0026423014081082305, -0.002765625569280217, 
    -0.0028755126407038365, -0.0029734536356629143, -0.0030610578814105616, 
    -0.0031398963856449267, -0.0032113523277331316, -0.0032765103154714604, 
    -0.0033360666579848718, -0.0033902861003363206, -0.0034389981061114464, 
    -0.0034816387288170401, -0.0035173373872884159, -0.0035450352895355832, 
    -0.0035636080309896503, -0.0035719880058944927, -0.0035692424131903602, 
    -0.0035546174541252291, -0.0035275232306271288, -0.003487486779367048, 
    -0.0034340595309826135, -0.0033667312479575121, -0.0032848630485317336, 
    -0.0031876716854807546, -0.0030742641367029482, -0.0029437372820034918, 
    -0.0027953398041305946, -0.0026286394808844025, -0.0024437298827629595, 
    -0.0022414043554829601, -0.0020232931066721275, -0.0017919530775000535, 
    -0.0015508517496453573, -0.0013042872944100553, -0.0010571930313481761, 
    -0.0008148940333914009, -0.00058279696657341387, -0.00036605918098839746, 
    -0.0001692719190073415, 3.8196261740423899e-06, 0.00015052697897798061, 
    0.00026934166500690136, 0.00035995982184318083, 0.00042322568929526973, 
    0.00046099064488853303, 0.00047591852567834117, 0.00047127197536487062, 
    0.00045067108438110029, 0.00041788164847177388, 0.00037660943997044877, 
    0.00033035036846759951, 0.00028227536096696277, 0.00023516711819773309, 
    0.00019138074806778624, 0.00015285101255100065, 0.00012111757989182045, 
    9.7352757056209916e-05, 8.2407451702472463e-05, 7.6846835099231631e-05, 
    8.0982184175098273e-05, 9.4905004403409766e-05, 0.00011850056111653127, 
    0.00015144875148523194, 0.00019320183252526793, 0.00024295307867795056, 
    0.00029959007011891553, 0.00036163186804385409, 0.00042719786305703641, 
    0.00049396265037871445, 0.00055916306660641201, 0.00061961920535502613, 
    0.00067178023221804327, 0.000711818805583034, 0.00073573600667090143, 
    0.0007395071137559654, 0.00071924544465569516, 0.000671389604157534, 
    0.00059289624528421274, 0.00048142502863670131, 0.0003354921838450342, 
    0.000154589654997253, -6.0740339739519047e-05, -0.00030889109977537372, 
    -0.00058723174408679686, -0.00089217926757603674, -0.001219334114149999, 
    -0.0015636202487713296, -0.0019194746566281791, -0.002281018392584315, 
    -0.0026422543682315287, -0.0029972418649218393, -0.003340256715777284, 
    -0.0036659340462329875, -0.0039693744305795099, -0.0042462538282261693, 
    -0.0044929064015208787, -0.0047064224766039395, -0.0048847433619846371, 
    -0.0050267346585014892, -0.0051322450826085629, -0.0052021255560412896, 
    -0.0052382267412556553, -0.0052433727775018143, -0.0052213107548665346, 
    -0.0051766302305120806, -0.0051146532738712931, -0.0050412737711950911, 
    -0.0049627641128553246, -0.0048855531976883283, -0.0048159861749721665, 
    -0.0047600823946640728, -0.0047232913030614996, -0.0047102939213021638, 
    -0.0047248178180058983, -0.0047695083988786259, -0.0048458300182998388, 
    -0.0049539991436162159, -0.0050929397982534107, -0.0052602610620906811, 
    -0.0054522957582941725, -0.0056641619389570892, -0.0058898979325817799, 
    -0.0061226627872934701, -0.0063550075760101252, -0.0065791701577062149, 
    -0.006787389153518235, -0.0069722037225150614, -0.0071266977383192941, 
    -0.0072447001631129118, -0.007320940638612914, -0.007351161225827442, 
    -0.0073322013169439286, -0.0072620298473514248, -0.0071397440323844137, 
    -0.0069655214877807521, -0.0067405304695679191, -0.0064668185236918096, 
    -0.0061471678006527718, -0.0057849726199879865, -0.0053841186852108544, 
    -0.0049488819196902957, -0.0044838310897856223, -0.0039937504268747039, 
    -0.0034835552725922436, -0.0029582366759007277, -0.0024228085766216227, 
    -0.0018822893246815678, -0.0013416903499995285, -0.00080601209902973834, 
    -0.00028021341375732617, 0.00023082555272038683, 0.00072238104302578467, 
    0.0011899657918781996, 0.0016294277323899153, 0.0020370483349273711, 
    0.0024096571498954042, 0.0027447507741980102, 0.0030405985294983616, 
    0.0032963533608744112, 0.0035121289780578394, 0.0036890393731953399, 
    0.0038292033358337278, 0.0039356896020841074, 0.0040124056180820371, 
    0.0040639539384508209, 0.0040954295992942247, 0.0041122246600725602, 
    0.0041198096063847951, 0.0041235533055796608, 0.0041285545226198679, 
    0.0041394943570874157, 0.0041605374686896398, 0.0041952346784726981, 
    0.004246465506691369, 0.0043164008300613441, 0.0044064739673786626, 
    0.004517392482927084, 0.0046491396860256383, 0.0048010387681919784, 
    0.0049717960074197416, 0.0051595784530154322, 0.005362100298110596, 
    0.0055766911141284211, 0.0058003799973056552, 0.006029950606888281, 
    0.0062619871801509255, 0.006492897198317118, 0.0067189430376090285, 
    0.0069362642453661685, 0.0071409090203032695, 0.007328880089782914, 
    0.0074962071994393057, 0.007639016742345732, 0.0077536252828110021, 
    0.0078366104739541129, 0.0078848954535710239, 0.0078958553035715449, 
    0.0078674233966823416, 0.0077982496028669501, 0.0076878732342761328, 
    0.0075368850425992749, 0.0073470410722643927, 0.0071213108365171208, 
    0.0068637984371679225, 0.0065796016411648556, 0.0062745878641249442, 
    0.0059551876322437294, 0.0056281849612861258, 0.0053005326376356042, 
    0.004979179068419182, 0.004670904451108647, 0.0043821590897943205, 
    0.0041188660708009871, 0.0038862603143100583, 0.0036886944572309109, 
    0.003529479984222904, 0.0034107611258004538, 0.0033334272932565349, 
    0.0032970993944577663, 0.0033001904712394916, 0.0033400069525760506, 
    0.0034129136171755898, 0.0035145412400143052, 0.0036399760402360121, 
    0.0037839644970734296, 0.0039410821059202607, 0.0041058957507111504, 
    0.0042730946915171264, 0.0044376123288563185, 0.0045947274207152585, 
    0.0047401398735822421, 0.0048700700180161266, 0.004981313618040677, 
    0.005071332545793404, 0.0051383072612221263, 0.005181182350644813, 
    0.005199655248464964, 0.0051941667044109021, 0.0051658081840960596, 
    0.0051162336390567636, 0.005047513994014213, 0.0049620189047258527, 
    0.0048622363435358966, 0.0047506541103849555, 0.0046296488803486049, 
    0.0045014412121729174, 0.0043681026908714508, 0.0042316013753601195, 
    0.0040938602397684112, 0.0039568292301452113, 0.003822538180888675, 
    0.0036931410307186985, 0.0035709259749821644, 0.0034583087120455681, 
    0.0033578097346767546, 0.0032720107872014647, 0.0032034579043732267, 
    0.00315454513560065, 0.0031273415589444971, 0.0031233774667472685, 
    0.003143392463901616, 0.003187106727067139, 0.0032529747535197792, 
    0.0033380407074432481, 0.0034378843253228637, 0.0035466657664644219, 
    0.0036572961175855923, 0.0037616828639784106, 0.0038510766552558727, 
    0.0039164488214102795, 0.0039489220996907952, 0.0039401965750476432, 
    0.0038829819586002853, 0.0037713597549074197, 0.0036011145734709117, 
    0.0033699927528392823, 0.0030778550853515661, 0.0027267449389714537, 
    0.0023208404273055336, 0.0018662636595933421, 0.0013708154323868705, 
    0.00084361025980842126, 0.00029468000477326887, -0.00026544012643445278, 
    -0.00082607453333216781, -0.0013767277516830432, -0.0019073323471642397, 
    -0.0024084318679193101, -0.0028713416950537688, -0.003288242907536325, 
    -0.0036522808093578918, -0.0039576334611763943, -0.0041995540513930984, 
    -0.0043744350969679331, -0.0044798193140570455, -0.0045144126141899426, 
    -0.0044780708450346271, -0.0043717755290139538, -0.0041975953513507499, 
    -0.0039586541445345048, -0.0036590555004099913, -0.0033037829166155503, 
    -0.0028985528386826871, -0.002449627744233315, -0.0019636353431863192, 
    -0.0014473843646786325, -0.00090771616354751595, -0.00035136233513707611, 
    0.00021519175939314008, 0.00078580945480082173, 0.0013547874937125596, 
    0.0019169325424326982, 0.002467610961360024, 0.0030028192513671791, 
    0.0035192864028999842, 0.0040145666428528385, 0.0044871753409734027, 
    0.0049366646785741191, 0.0053636586242154401, 0.0057698038809725462, 
    0.0061576258488456707, 0.0065303294686554474, 0.0068915108522165812, 
    0.0072448961923627046, 0.0075940681083159255, 0.0079422373455986777, 
    0.0082920922548493734, 0.0086456977635005535, 0.009004422160004447, 
    0.0093689035616474382, 0.0097390187242496328, 0.010113843362583908, 
    0.010491605029641362, 0.010869652309020135, 0.011244436290065662, 
    0.011611531260026408, 0.011965718089630128, 0.012301119178655057, 
    0.012611404877129032, 0.012890041441989889, 0.013130537745738817, 
    0.013326740147698428, 0.013473059301886877, 0.013564702484580004, 
    0.013597861512443254, 0.013569856629476728, 0.013479255775599493, 
    0.013325935167988091, 0.013111070633714183, 0.01283704917379574, 
    0.012507286516701454, 0.012126005318983278, 0.011697979849670609, 
    0.011228242820079762, 0.010721863727299753, 0.010183697182961761, 
    0.0096181695060758056, 0.0090290721104000268, 0.008419450593751843, 
    0.0077914805905307987, 0.0071464743987412638, 0.0064849355215168894, 
    0.0058066828595278392, 0.0051110876937575543, 0.0043973206860528158, 
    0.0036646615502377317, 0.0029127716792955189, 0.0021419607217924622, 
    0.001353347671947405, 0.0005489886479405037, -0.00026810641370570424, 
    -0.0010939610538978416, -0.0019236953948905484, -0.0027515864853125275, 
    -0.0035711828035775981, -0.0043754122991917985, -0.0051567681494741812, 
    -0.0059074883162879557, -0.0066198211293773089, -0.0072862636175844457, 
    -0.0078998277718304328, -0.0084543166508086274, -0.0089445301784259763, 
    -0.0093664220892494265, -0.0097172421540605448, -0.0099955288101456242, 
    -0.010201097695454298, -0.010334922274792336, -0.010399001992222654, 
    -0.010396151517762277, -0.010329822090253366, -0.010203889683578805, 
    -0.010022499334879146, -0.0097899114413185322, -0.0095103869823257112, 
    -0.0091881367405989792, -0.0088272898212425743, -0.0084318927319685447, 
    -0.0080059362700984418, -0.0075533896087038562, -0.0070782104174384845, 
    -0.0065843575942744932, -0.0060757670257789954, -0.0055563674779976532, 
    -0.0050300273466638255, -0.0045005752946753273, -0.0039717869710172941, 
    -0.003447392530245977, -0.0029310988143357872, -0.0024265728943629983, 
    -0.0019374176070636314, -0.0014671221194900311, -0.001018929875464068, 
    -0.00059569957615826453, -0.00019974724804194889, 0.00016731617207491677, 
    0.00050467335935365954, 0.00081232723164171964, 0.0010910280068439175, 
    0.0013420840462708031, 0.0015671158172536649, 0.0017677474172745581, 
    0.0019453001267848566, 0.0021005539720070666, 0.0022335588649550937, 
    0.0023435529972288252, 0.0024289862172333899, 0.0024876017202797107, 
    0.0025166414148792668, 0.0025130704881467713, 0.0024738197561751402, 
    0.0023960716115037305, 0.0022774839509661525, 0.0021163984558912616, 
    0.001912002430038985, 0.0016643992661916041, 0.001374653642879402, 
    0.0010447888060846184, 0.00067774852127905989, 0.0002773368526075296, 
    -0.00015184468668096943, -0.00060446644770411847, -0.0010745616435806206, 
    -0.001555630352102571, -0.0020408097733333802, -0.0025230802303984555, 
    -0.0029955328597746867, -0.00345163884189253, -0.0038855166199360898, 
    -0.0042921930631304589, -0.0046677848846916606, -0.0050095934738538682, 
    -0.00531613131737361, -0.0055870722785121727, -0.0058230897899894472, 
    -0.0060256857557959096, -0.0061969322217615931, -0.0063392279008791848, 
    -0.0064550205896402877, -0.0065465770772032946, -0.0066157685130258321, 
    -0.0066639438655328991, -0.0066918069947384919, -0.0066994152238693512, 
    -0.0066861883766466965, -0.006650919793588549, -0.0065918763153169739, 
    -0.0065068843156976686, -0.0063935207482367284, -0.0062493313895748154, 
    -0.0060721259609295541, -0.0058603549040430877, -0.0056134728902274859, 
    -0.0053322936147708541, -0.0050193236926984828, -0.0046789152847965263, 
    -0.0043173624525032371, -0.0039427805774788337, -0.0035648584597592703, 
    -0.0031944268230423931, -0.0028429262331589981, -0.0025217733901195167, 
    -0.0022417499868452677, -0.0020123964118949076, -0.0018415795612061097, 
    -0.0017351581318832137, -0.0016969553561978139, -0.0017289426392901356, 
    -0.001831679887774532, -0.0020048337802897899, -0.0022475842073269052, 
    -0.0025587598308712462, -0.0029366894293086855, -0.0033788465782876643, 
    -0.0038814655241916738, -0.0044392082513611784, -0.0050449913076527344, 
    -0.0056899648835129863, -0.0063636608860659768, -0.0070542929861558091, 
    -0.0077491346601849167, -0.0084349732518750192, -0.0090985491122270151, 
    -0.0097269743910750397, -0.010308124138716613, -0.010830982051343202, 
    -0.011286036896269695, -0.011665619400671238, -0.011964167689999177, 
    -0.012178450735161493, -0.012307591166061284, -0.012353033116689496, 
    -0.01231838452745878, -0.012209142080607086, -0.012032393720036302, 
    -0.011796503251519026, -0.011510712694076747, -0.011184770808279204, 
    -0.010828523934888607, -0.010451489216685898, -0.01006240877892153, 
    -0.0096688543220274318, -0.0092768822639611292, -0.0088908105839760245, 
    -0.0085131319649054005, -0.0081445456354438516, -0.0077842096523985755, 
    -0.0074299884436805994, -0.0070789282465898882, -0.0067275867425346074, 
    -0.0063724388152066333, -0.0060101492141827013, -0.0056377865275600483, 
    -0.0052529135768944642, -0.0048536274793981489, -0.0044385744613253779, 
    -0.0040069062583176574, -0.0035583567986242361, -0.0030932838166902823, 
    -0.0026128653299636352, -0.0021192327318843552, -0.0016156469350546772, 
    -0.0011066078883247006, -0.00059788726189262495, -9.6489515666724088e-05, 
    0.00038948811696359518, 0.00085114626284514051, 0.001279190334225739, 
    0.0016643602094078966, 0.0019979654911405536, 0.0022724373510946581, 
    0.00248175799279505, 0.0026218593039126592, 0.0026908842523632017, 
    0.0026892844114494445, 0.0026198022500318074, 0.0024872951685430745, 
    0.0022984638948567019, 0.0020614606293447874, 0.0017855020672745605, 
    0.001480385817257858, 0.0011560847744840914, 0.00082229592232091833, 
    0.00048801247811144108, 0.00016115030563907244, -0.00015178367995504296, 
    -0.00044576917666637559, -0.00071725088328889321, 
    -0.00096379634723959759, -0.0011835501842250135, -0.0013747259543120864, 
    -0.0015350220291563779, -0.0016612914205667165, -0.0017495047609974355, 
    -0.0017950021958101502, -0.0017929483709403548, -0.0017390021499708488, 
    -0.0016300197248520813, -0.0014647665941159194, -0.0012445190889231609, 
    -0.00097343370726167935, -0.00065869868733344167, 
    -0.00031030725026275156, 5.9361435004761382e-05, 0.00043640530108213146, 
    0.00080622476839440683, 0.0011545548029709238, 0.0014682893220893168, 
    0.0017362120057721373, 0.0019493677242212115, 0.0021013112745026205, 
    0.0021881717557030549, 0.00220854558611892, 0.002163517416163004, 
    0.0020564525803906429, 0.0018928638096328818, 0.0016800998745159323, 
    0.001426948386773509, 0.0011432485264226309, 0.00083927361462724447, 
    0.00052521009046272273, 0.00021062762659592525, -9.5869199958462033e-05, 
    -0.00038695835781252285, -0.00065676124182831341, 
    -0.00090077478638996868, -0.0011158549142889335, -0.0013001145618091498, 
    -0.0014528042243750589, -0.0015743054959689571, -0.0016661010507558686, 
    -0.0017308639195410631, -0.0017723867699062359, -0.0017950966295493041, 
    -0.0018035342077457692, -0.001801341827273054, -0.0017902646593236709, 
    -0.0017690614214329295, -0.0017331102481122967, -0.0016742359285412997, 
    -0.0015815452591275098, -0.001442583836146708, -0.0012451065788954591, 
    -0.00097890564719341861, -0.00063749980085793013, -0.0002197436623338006, 
    0.00026933848782224553, 0.00081815602366094842, 0.0014090211822730934, 
    0.0020190796673332911, 0.0026220574015404499, 0.0031904227387606855, 
    0.0036976444868440429, 0.0041210828578331265, 0.0044440767741846582, 
    0.0046574712213361819, 0.0047603428519039492, 0.0047594898669153429, 
    0.0046683636021177879, 0.0045056019251875409, 0.0042936858016237025, 
    0.0040576231610244288, 0.0038239053262480727, 0.0036192748555904366, 
    0.0034689863760790658, 0.0033952235185476941, 0.0034153857127582989, 
    0.0035403692176263811, 0.0037744070060487444, 0.0041144645135569877, 
    0.0045517818676621274, 0.0050715382716513858, 0.005655527467089176, 
    0.0062822444473098777,
  // Fqt-total(6, 0-1999)
    0.99999999999999956, 0.99525477896692105, 0.98118203492540246, 
    0.95825887377193464, 0.92724489406017752, 0.88913362356896086, 
    0.84509179666781231, 0.79639235211502957, 0.74434703577655836, 
    0.69024387926757058, 0.63529367096269818, 0.58058806550855091, 
    0.52707054370528916, 0.475520106274198, 0.42654649842420117, 
    0.38059511041952593, 0.33795926501999224, 0.29879758152042524, 
    0.26315418310620686, 0.23097993873844364, 0.20215320403185549, 
    0.17649903200194833, 0.15380616303829428, 0.13384144315577334, 
    0.11636161981261176, 0.10112259128284649, 0.087886366084905562, 
    0.076426022433305943, 0.066528999078692433, 0.057999053385039662, 
    0.05065718871976075, 0.044341816785349569, 0.038908395527856937, 
    0.034228699195329303, 0.030189869056588551, 0.026693332357427726, 
    0.02365366227294614, 0.020997429060249363, 0.018662061059469638, 
    0.016594755756398284, 0.014751418347413437, 0.013095663155129717, 
    0.011597836530745011, 0.010234095539049233, 0.0089855167888666081, 
    0.0078372446681394085, 0.0067776960976422196, 0.0057978161358054753, 
    0.0048904180068153518, 0.0040495994418185497, 0.0032702716880185292, 
    0.002547798935699769, 0.0018777492351860668, 0.0012557654567936236, 
    0.00067753298161334573, 0.00013882468427818558, -0.00036439010252255709, 
    -0.00083580984043616214, -0.0012786664768482897, -0.0016956013968936201, 
    -0.0020885896396976283, -0.0024589100911700792, -0.0028071685662905978, 
    -0.0031333618895626361, -0.0034369817024644377, -0.0037171194639840448, 
    -0.0039726039225416046, -0.00420212526683036, -0.0044044008307353175, 
    -0.0045783470308469465, -0.0047232648476469305, -0.0048390013292585595, 
    -0.0049260691605052601, -0.0049856826419445435, -0.0050197031242487722, 
    -0.0050305105226369842, -0.0050207954850895299, -0.0049933246595873478, 
    -0.0049506995099818226, -0.0048951447311024769, -0.0048283547970490058, 
    -0.0047514192387787717, -0.0046648268211152118, -0.0045685523015440467, 
    -0.0044622062809636575, -0.0043452294042130857, -0.0042171019605832987, 
    -0.0040775481725176584, -0.0039267138625991311, -0.0037653001167647481, 
    -0.0035946387890787913, -0.0034167133444436256, -0.0032341284543008272, 
    -0.0030500289611085541, -0.0028679869896152924, -0.0026918461630510235, 
    -0.0025255467158731009, -0.0023729304906691651, -0.002237556816457438, 
    -0.0021225266217815954, -0.0020303368134859372, -0.0019627828792912337, 
    -0.0019208902486672662, -0.0019048902757129215, -0.0019142261982539712, 
    -0.0019475786111095839, -0.0020029169326895107, -0.0020775514106679649, 
    -0.0021682000199133604, -0.0022710559712161003, -0.0023818655893619186, 
    -0.0024960198711858773, -0.0026086581892258019, -0.0027148115991756415, 
    -0.0028095578414238428, -0.002888223571580517, -0.0029465928503258211, 
    -0.0029811355967446348, -0.0029892074390475399, -0.0029692134378993653, 
    -0.002920706226236326, -0.0028444053296286711, -0.0027421383823877724, 
    -0.0026167054909163011, -0.002471675122358677, -0.0023111292426190025, 
    -0.0021393681072144136, -0.001960613194117322, -0.0017787324038041968, 
    -0.0015970191646417717, -0.0014180521074598385, -0.0012436455299469297, 
    -0.0010748832697414354, -0.00091221715053920946, -0.00075560256496488268, 
    -0.00060466408703733631, -0.00045884417887661022, 
    -0.00031753290084062766, -0.000180178802841827, -4.6355180602145834e-05, 
    8.4194226333806244e-05, 0.00021153800997553114, 0.00033555299025671943, 
    0.00045593348020485293, 0.0005722035211700203, 0.0006837361540122809, 
    0.00078978332400788396, 0.00088950402190597167, 0.00098200815135671008, 
    0.0010663971932040239, 0.0011418034619149165, 0.0012074145197854302, 
    0.0012624846556100883, 0.0013063252451014501, 0.001338297787047695, 
    0.0013577982321348104, 0.0013642709389503707, 0.0013572302541645573, 
    0.0013362957248121334, 0.0013012175617495027, 0.0012518988983820664, 
    0.0011883860984968628, 0.0011108561467767627, 0.0010195847071192783, 
    0.00091493350009123409, 0.00079734643140365108, 0.00066738045110067024, 
    0.00052573556770289603, 0.00037331560751164715, 0.00021126139169002251, 
    4.0993752942961017e-05, -0.00013576509746424987, -0.00031699244527922586, 
    -0.00050038206430710658, -0.0006834035837600342, -0.00086338953902874069, 
    -0.0010376462389358851, -0.0012035816672784103, -0.0013588329176321525, 
    -0.0015013710281615751, -0.0016296000138260125, -0.0017424081837691995, 
    -0.0018392084065980156, -0.0019199361361551591, -0.0019850340844102914, 
    -0.0020353978240950895, -0.0020723098442491533, -0.0020973620743531957, 
    -0.0021123670413312717, -0.0021192684585458342, -0.0021200615285353209, 
    -0.0021167165077440658, -0.002111101021632381, -0.0021049226267199008, 
    -0.0020996619249531038, -0.0020965268935761562, -0.0020964145065900408, 
    -0.0020998726638208334, -0.0021070853202886271, -0.0021178514395578758, 
    -0.0021315740408027503, -0.0021472572880879902, -0.0021635175920283042, 
    -0.0021786109785353175, -0.0021904849386545923, -0.0021968486389378821, 
    -0.0021952614778127915, -0.0021832404822436334, -0.0021583692629613713, 
    -0.0021184066630375166, -0.0020613828895964417, -0.0019856777219800785, 
    -0.0018900659518995761, -0.0017737470628375379, -0.0016363401412333657, 
    -0.0014778598924116996, -0.0012986779975719099, -0.0010994740518579132, 
    -0.00088119740766290366, -0.00064503476125725391, 
    -0.00039239549360171264, -0.00012492909987076462, 0.00015544599505827689, 
    0.00044649371157366323, 0.00074560079923970753, 0.0010497273148519612, 
    0.0013553659739198956, 0.0016585301133755393, 0.0019547648605935108, 
    0.0022392087935230636, 0.002506692581875056, 0.0027518800920437007, 
    0.0029694444427722866, 0.0031542726263635978, 0.0033016733696116054, 
    0.0034075893460207901, 0.0034687867120425319, 0.0034830231895294013, 
    0.0034491762086968519, 0.0033673294413565512, 0.0032388069573157912, 
    0.0030661540594557569, 0.0028530529316366363, 0.0026041853802360351, 
    0.0023250384408071167, 0.0020216743294947906, 0.0017004764402166882, 
    0.0013678877111853625, 0.0010301682828967079, 0.00069318374109588929, 
    0.0003622345298969389, 4.1936572031240504e-05, -0.00026385681065513669, 
    -0.00055209213019742219, -0.0008205260686107973, -0.0010677177767973423, 
    -0.0012930102433289892, -0.0014964998797901943, -0.001678992615493547, 
    -0.001841935874299209, -0.0019873420932842744, -0.0021176892294311927, 
    -0.0022358064277624326, -0.002344761578632865, -0.0024477307990732741, 
    -0.0025478540010483944, -0.0026480761754172871, -0.0027509670446502822, 
    -0.002858540153171807, -0.0029720779584937944, -0.0030920100111557036, 
    -0.0032178282409931064, -0.0033481006362385646, -0.0034805461558488991, 
    -0.003612198738811319, -0.0037396155231141509, -0.0038591355175591315, 
    -0.00396714677869599, -0.0040603538427001389, -0.0041360008958422328, 
    -0.0041920635365918528, -0.0042273638746607202, -0.0042416121810542294, 
    -0.0042353648012761272, -0.0042099074321500221, -0.0041670651632500005, 
    -0.0041089589133536074, -0.004037730154385656, -0.0039552692952371836, 
    -0.0038629647239009483, -0.0037615175083258201, -0.0036508522969219905, 
    -0.0035301311903875843, -0.0033978873052723985, -0.0032522630233525239, 
    -0.0030913219348952122, -0.0029134080143830197, -0.0027174932984158841, 
    -0.0025034987914822086, -0.0022725282010958069, -0.0020270021912181359, 
    -0.0017706784355311503, -0.0015085633270186978, -0.0012467181445954911, 
    -0.00099197168149706811, -0.00075158167590386551, -0.0005328649887782628, 
    -0.00034281883074660432, -0.00018776869260314676, 
    -7.3072904738666304e-05, -2.8867658267848077e-06, 1.9980825857798186e-05, 
    -5.8753860894611497e-06, -8.0495826526568088e-05, 
    -0.00020265841362166121, -0.00037003637026983315, 
    -0.00057937668928765109, -0.00082666264542357421, -0.0011072467814440723, 
    -0.0014159408088433734, -0.0017470583188287671, -0.0020944456010840973, 
    -0.0024515040737156111, -0.0028112543269147579, -0.003166433172666158, 
    -0.003509653906206364, -0.0038336023177302941, -0.0041312680083798242, 
    -0.0043961818351646127, -0.0046226418957902044, -0.0048059177177537295, 
    -0.0049424111106114643, -0.005029769744430368, -0.0050669521098365752, 
    -0.0050542381526940874, -0.0049931887874190856, -0.0048865551209864144, 
    -0.0047381453112816524, -0.0045526510344600724, -0.0043354404008387618, 
    -0.004092321708536165, -0.0038292909665532814, -0.003552277198679277, 
    -0.0032668996257989142, -0.0029782441912130407, -0.0026906872138116912, 
    -0.0024077673786005675, -0.0021321113631911958, -0.0018654375044663534, 
    -0.0016086307156474473, -0.0013618821757060483, -0.0011248834117041201, 
    -0.00089703969854973821, -0.00067768120695270375, 
    -0.00046624925328018411, -0.00026243777007113167, 
    -6.6279314016796635e-05, 0.00012184275809270474, 0.00030124836632278271, 
    0.0004710603314020733, 0.00063034376571416753, 0.00077826007343212336, 
    0.00091420985488103285, 0.0010379503169413596, 0.0011496749793800263, 
    0.0012500428053970468, 0.0013401492141026225, 0.0014214565533474841, 
    0.0014956781856418093, 0.0015646480196810171, 0.0016301851307153814, 
    0.0016939798604330277, 0.0017575038680285125, 0.0018219648254047345, 
    0.001888281657429437, 0.0019570974641189101, 0.0020287940939632712, 
    0.0021035196168256408, 0.0021812097447672278, 0.0022615955018720053, 
    0.0023442059938355649, 0.0024283530337491639, 0.0025131053543799805, 
    0.0025972617816379675, 0.0026793282209685207, 0.0027575044698192512, 
    0.0028296999605811361, 0.002893570097146741, 0.0029466007076143158, 
    0.0029862276093916016, 0.0030100013668114519, 0.0030157781438901209, 
    0.0030019364180623098, 0.0029675746208344444, 0.0029126852175230152, 
    0.002838281381576636, 0.002746463429833992, 0.0026404128170535112, 
    0.0025243038884238036, 0.0024031392400180817, 0.0022825026804188047, 
    0.0021682447702359316, 0.0020661320009655476, 0.0019814710561297591, 
    0.001918756140344277, 0.0018813534959225106, 0.0018712638312989834, 
    0.0018889791928094262, 0.0019334482790216987, 0.00200213985268374, 
    0.0020912205049825124, 0.0021957999978446646, 0.002310242329983172, 
    0.0024285096736856369, 0.002544521342698051, 0.0026525039702833659, 
    0.0027473128372386721, 0.002824708097320416, 0.0028815641952899245, 
    0.0029160061213450287, 0.0029274557729300744, 0.0029165844441208576, 
    0.0028851792522500874, 0.0028359244717994056, 0.0027721338757509496, 
    0.0026974636174847254, 0.0026156365660760209, 0.002530204029955361, 
    0.0024443580444156636, 0.0023608004064202821, 0.0022816623821706908, 
    0.0022084784970962694, 0.0021421999294385006, 0.0020832500029499016, 
    0.0020316123351398542, 0.0019869425171858066, 0.0019486949257790051, 
    0.0019162599747324389, 0.0018890899460674837, 0.0018668103562227529, 
    0.0018492934450550216, 0.0018366756877691011, 0.0018293271640488634, 
    0.0018277588144164564, 0.0018324950417754231, 0.0018439264047329052, 
    0.0018621580086400195, 0.0018868843670492442, 0.0019172933005459666, 
    0.0019520228824510316, 0.0019891560148138738, 0.0020262853102432322, 
    0.0020606190790852619, 0.0020891284280242475, 0.002108711995361614, 
    0.0021163495818250938, 0.0021092272513188923, 0.0020848268394845788, 
    0.0020409947779681465, 0.0019759911720126653, 0.0018885336074148792, 
    0.0017778302414028786, 0.0016436135981684656, 0.0014861571571927411, 
    0.0013062825347051066, 0.0011053546156464199, 0.00088526752616579531, 
    0.0006484224267524402, 0.00039770712034781171, 0.00013646633102289818, 
    -0.00013154003653356532, -0.00040219507070953365, 
    -0.00067110490789983198, -0.00093370551665363183, -0.0011853784814610663, 
    -0.0014215878127608733, -0.0016380140157720505, -0.0018306897537622303, 
    -0.0019961274957754661, -0.0021314204557806005, -0.0022343334056859209, 
    -0.0023033606889190064, -0.0023377579669780963, -0.002337550314718368, 
    -0.0023035099733420918, -0.0022371151325882785, -0.0021404865340579502, 
    -0.002016308682748465, -0.0018677367494585517, -0.0016982882926151353, 
    -0.0015117325360240682, -0.0013119730616071347, -0.0011029358343460417, 
    -0.00088846501137609501, -0.00067222277210565154, 
    -0.00045758871666686088, -0.00024757383803565434, 
    -4.4717692782763799e-05, 0.00014899556417596822, 0.00033220742302511759, 
    0.00050422342793039808, 0.00066500559782202808, 0.00081512584848565564, 
    0.00095567601350747945, 0.0010881379304889553, 0.0012142300888630174, 
    0.0013357227796012266, 0.0014542556891142858, 0.0015711642971869789, 
    0.001687333039138428, 0.0018030820120594779, 0.0019180970472939744, 
    0.0020314113429803467, 0.0021414197030843502, 0.0022459526580033964, 
    0.0023423801173453741, 0.0024277547475337288, 0.0024989838104320194, 
    0.0025530178966409784, 0.0025870511298541113, 0.0025987091648176776, 
    0.0025862222267282876, 0.0025485528276506519, 0.0024854899180452605, 
    0.0023976797486331019, 0.0022866050591719808, 0.0021545134935304715, 
    0.0020042921302349656, 0.0018393137314598167, 0.0016632528350401896, 
    0.0014799094921282535, 0.0012930327812122964, 0.0011061670678621138, 
    0.00092250728744259342, 0.00074478048565840152, 0.00057514309819945439, 
    0.00041511917658234898, 0.00026557367296246712, 0.00012672312842630144, 
    -1.8264485956392496e-06, -0.00012102396605924287, 
    -0.00023230251600035655, -0.00033751110261225607, 
    -0.00043884122494293996, -0.00053874017192574297, 
    -0.00063981445272521316, -0.00074472168830668189, -0.0008560456080094434, 
    -0.00097616073978782801, -0.0011070923774184655, -0.0012503757835441757, 
    -0.0014069180437121052, -0.0015768834678629626, -0.0017595943030539677, 
    -0.0019534737194358037, -0.0021560263087450453, -0.0023638628089564292, 
    -0.0025727682916939299, -0.0027778123244246054, -0.0029735026956238019, 
    -0.0031539821745541602, -0.0033132675935568716, -0.0034455171843676192, 
    -0.0035453119138912988, -0.0036079368634150295, -0.0036296396575280958, 
    -0.0036078504886789841, -0.003541343653638175, -0.0034303210548712673, 
    -0.0032764290272347986, -0.0030826884447104196, -0.0028533567473800329, 
    -0.0025937213572223335, -0.0023098504383665119, -0.0020083123547936089, 
    -0.0016958889589723028, -0.0013792960592242977, -0.001064936977841061, 
    -0.00075869309773481054, -0.00046576567145290742, 
    -0.00019056471148481017, 6.3354305761140667e-05, 0.00029331711048304597, 
    0.00049752082254095234, 0.00067501310824217588, 0.00082564458234701832, 
    0.00095001144041644209, 0.0010493880653865088, 0.0011256331910312362, 
    0.0011810882181150003, 0.0012184558648054053, 0.0012406680101936778, 
    0.0012507471197696367, 0.0012516761190199733, 0.0012462636319785158, 
    0.0012370276948666793, 0.0012260761268824891, 0.0012150069412838619, 
    0.0012048188271631646, 0.001195841970304101, 0.0011877172892382668, 
    0.0011794095549009958, 0.0011692904192562132, 0.0011552638940980943, 
    0.0011349475119417369, 0.0011058660824916722, 0.0010656444646587123, 
    0.0010121755809614078, 0.00094373464149207246, 0.00085905546651173263, 
    0.00075734509405221034, 0.00063826074258067889, 0.00050187612805684741, 
    0.00034863223830060769, 0.00017929956243815606, -5.0494235587312728e-06, 
    -0.00020305733916138233, -0.00041309322993572667, -0.0006332609732882335, 
    -0.00086140430934948339, -0.0010951137496332196, -0.001331727012651497, 
    -0.0015683390394704848, -0.0018018109941972369, -0.0020287979345666551, 
    -0.0022457979349371862, -0.0024492451811147192, -0.0026356347927580129, 
    -0.0028016943959028044, -0.0029445707365300922, -0.0030619991033773446, 
    -0.003152445379791805, -0.0032151761034491327, -0.0032502783521750739, 
    -0.0032586072198483667, -0.0032416923110435399, -0.0032015988185997049, 
    -0.0031407726715842899, -0.0030618719007050967, -0.0029675989790973372, 
    -0.0028605512743218996, -0.002743095179276886, -0.0026172762328625482, 
    -0.0024847717897484899, -0.002346885092458716, -0.0022045758747220065, 
    -0.002058514626528481, -0.0019091592574055104, -0.0017568444840135671, 
    -0.0016018632793534217, -0.0014445429447705722, -0.0012853137826450932, 
    -0.0011247608742576294, -0.0009636623484050457, -0.00080301767375605708, 
    -0.00064406919368571215, -0.00048830793930323925, 
    -0.00033747729925636088, -0.00019355714733926244, 
    -5.8740783443290707e-05, 6.4619390195554767e-05, 0.00017407391043417636, 
    0.00026716049942976904, 0.00034149912026922767, 0.00039489159762057631, 
    0.00042542891560703251, 0.00043160160377509024, 0.00041240496218877809, 
    0.00036743385234919683, 0.00029695885436386828, 0.00020197966039818931, 
    8.4243009625918158e-05, -5.3770199081769538e-05, -0.00020890157778786001, 
    -0.00037739578201533388, -0.00055502464499584123, 
    -0.00073724964419034369, -0.00091941504309823519, -0.0010969645732644992, 
    -0.0012656656389019489, -0.0014218378878756669, -0.0015625541341394544, 
    -0.0016858126605807295, -0.0017906410136356847, -0.0018771467300722261, 
    -0.0019464904395633878, -0.0020007947010408063, -0.002042999266178853, 
    -0.0020766523027490572, -0.0021056799997808185, -0.0021341296721450504, 
    -0.0021659056338799005, -0.0022045353729922626, -0.00225296830295544, 
    -0.0023134359789086932, -0.0023873711324204827, -0.0024754049589660967, 
    -0.002577403204419201, -0.0026925553083346513, -0.0028194743016835412, 
    -0.0029562852895283829, -0.0031007113054346822, -0.0032501328017062532, 
    -0.0034016349753026925, -0.0035520548540777554, -0.0036980301930939186, 
    -0.0038360658272166394, -0.0039626272683714169, -0.004074271139134362, 
    -0.0041678059466923045, -0.0042404805561174616, -0.0042901658692601763, 
    -0.0043155254628331864, -0.004316133321516597, -0.0042925221564891923, 
    -0.0042461587648252811, -0.0041793369964745067, -0.0040950012853098721, 
    -0.0039965278327671683, -0.0038874794392185926, -0.003771367864805713, 
    -0.003651436666101013, -0.0035304974325178085, -0.0034108180986875082, 
    -0.0032940809378624179, -0.0031814037985161856, -0.0030734141808106967, 
    -0.0029703602694403928, -0.0028722458960617728, -0.0027789706772054891, 
    -0.0026904628951326661, -0.0026067975583987605, -0.0025282940874335595, 
    -0.0024555807259270543, -0.0023896169371644582, -0.0023316580806700448, 
    -0.0022831690794313849, -0.0022456821244397737, -0.0022206179338049568, 
    -0.002209103417215327, -0.0022118012984431923, -0.0022287776541148564, 
    -0.0022594102622332068, -0.0023023497303172455, -0.0023555207286344118, 
    -0.0024161640917185101, -0.0024809164267323124, -0.0025459135420250064, 
    -0.0026069078172593616, -0.0026594128662536113, -0.0026988617072990525, 
    -0.002720784142307719, -0.0027210167358516476, -0.0026959100012528782, 
    -0.0026425504509465731, -0.0025589687189015646, -0.0024443253018991032, 
    -0.0022990562384625009, -0.0021249630319679046, -0.0019252261857977762, 
    -0.0017043401629142784, -0.0014679557401708211, -0.0012226413797042752, 
    -0.00097556858175815934, -0.00073413136001136464, 
    -0.00050554212801525681, -0.00029641855042917235, 
    -0.00011240646147939725, 4.2122652345330025e-05, 0.00016429468838534048, 
    0.00025282629523534864, 0.00030800802490455094, 0.00033157100783394249, 
    0.00032645571961537967, 0.00029651832239195001, 0.00024620384411687635, 
    0.00018021183673776328, 0.00010318791300842379, 1.945337936909349e-05, 
    -6.7204222658409751e-05, -0.00015368270422137106, 
    -0.00023764712544856905, -0.00031753803413965635, 
    -0.00039251679547196416, -0.00046235152167261299, 
    -0.00052725757367592756, -0.00058770987242603935, 
    -0.00064424095319675441, -0.00069725964947668878, 
    -0.00074687904329596337, -0.00079280860953772172, -0.0008342758676697249, 
    -0.00087001133147469282, -0.00089829560453859368, 
    -0.00091705168078190763, -0.00092399524570676282, 
    -0.00091681289821253129, -0.00089336968196386654, 
    -0.00085191962894304134, -0.00079130034157134769, 
    -0.00071110316638358295, -0.00061179133708229544, 
    -0.00049477387425281381, -0.00036240794063271617, 
    -0.00021795627229795355, -6.5475680588703334e-05, 9.0338035637432067e-05, 
    0.00024433101208784893, 0.00039110398675841506, 0.00052522174659069625, 
    0.0006414256501528989, 0.00073483446751395828, 0.0008011386621986611, 
    0.00083678790512625625, 0.00083916301218119266, 0.00080671990892155696, 
    0.00073910421967880962, 0.00063720358576069378, 0.00050313947498151202, 
    0.00034019463234591515, 0.00015267638057356824, -5.4279793625239819e-05, 
    -0.00027494490165060547, -0.00050326048005232705, 
    -0.00073310007821538164, -0.00095851852944635557, -0.0011739686110853386, 
    -0.0013744674003605072, -0.0015557128235845039, -0.001714148642511539, 
    -0.001846979380601306, -0.0019521462585802593, -0.0020282668183848043, 
    -0.0020745661150427448, -0.002090790618856446, -0.0020771343909112179, 
    -0.0020341669409079965, -0.0019627860628696134, -0.0018641770754657195, 
    -0.0017397890684127826, -0.0015913169833508393, -0.001420695566750208, 
    -0.001230090114335429, -0.0010218955647898977, -0.00079872934341038723, 
    -0.00056342796246251802, -0.00031903527215692, -6.880940198568798e-05, 
    0.00018377865053411331, 0.00043504193702290702, 0.00068106263518877936, 
    0.00091769768347879524, 0.0011406016394924948, 0.0013452819886828604, 
    0.0015272033639515538, 0.0016819362263897979, 0.0018053496214106158, 
    0.0018938217459372306, 0.0019444607595652296, 0.0019552896470306181, 
    0.001925400988062454, 0.0018550393861970736, 0.001745619175051859, 
    0.00159966468221704, 0.0014206878839185908, 0.0012129916577270164, 
    0.00098142896137105536, 0.00073113677361076449, 0.00046726076834849469, 
    0.00019470482305537331, -8.2063097079164481e-05, -0.00035913456180162794, 
    -0.0006332115368294991, -0.00090157540365537979, -0.00116201391366198, 
    -0.0014127349765438466, -0.0016522692016007528, -0.0018794125131150242, 
    -0.0020931846889805372, -0.0022928133168201941, -0.0024777286047090383, 
    -0.0026475569394223929, -0.0028021077996308644, -0.0029413399021420436, 
    -0.0030653124421869465, -0.0031741377832582257, -0.0032679201233010041, 
    -0.0033467020129241865, -0.0034104030562294775, -0.00345876557733177, 
    -0.0034913017126363679, -0.0035072501622083084, -0.0035055532958963216, 
    -0.0034848683003099643, -0.0034436161880966008, -0.0033800767968961165, 
    -0.003292515854981777, -0.0031793558219315849, -0.0030393531870712381, 
    -0.0028717767955432072, -0.0026765706523242346, -0.0024544722932995952, 
    -0.0022071019178637906, -0.0019369865032896594, -0.0016475477109326145, 
    -0.0013430431018599553, -0.0010284632329543646, -0.00070939823733323149, 
    -0.00039184795502213122, -8.2017000561475587e-05, 0.00021396217018641972, 
    0.00049031770457339246, 0.00074194130268286204, 0.00096466649013283263, 
    0.0011554748478395612, 0.0013126320068995165, 0.0014357393202422857, 
    0.0015257110133818617, 0.0015846973788401074, 0.0016159555635700915, 
    0.001623684872095528, 0.0016128374894244857, 0.0015889038758916528, 
    0.0015577053517397865, 0.0015251874712666955, 0.0014972275454142865, 
    0.0014794567779315396, 0.0014771055781318818, 0.0014948541162000241, 
    0.0015366943701354187, 0.0016057960916107954, 0.001704383566710183, 
    0.0018336187066259606, 0.0019934998799509057, 0.0021828025426124478, 
    0.0023990451943093371, 0.0026385403421640787, 0.0028964940053839011, 
    0.0031671823436441376, 0.0034441829966832295, 0.0037206443995921007, 
    0.0039895640434846171, 0.0042440494071381589, 0.0044775479495399798, 
    0.0046840376463749651, 0.0048581814935046135, 0.0049954576404752536, 
    0.0050922665042635986, 0.0051460336341703676, 0.0051552768406472448, 
    0.0051196567505318565, 0.005039988416679117, 0.0049181986195695748, 
    0.0047572328697967877, 0.0045609062707282193, 0.0043336952082683906, 
    0.0040805027018185952, 0.0038064017433159145, 0.0035163814660403763, 
    0.0032151228360405852, 0.002906811747513408, 0.002595012113853548, 
    0.0022825913174426881, 0.0019717138214137117, 0.0016638669988407462, 
    0.0013599510760161707, 0.0010603852137045808, 0.00076523704570002926, 
    0.00047436283425607035, 0.000187541368113155, -9.5393034400218147e-05, 
    -0.000374429027371896, -0.00064926237394764548, -0.00091919630179750165, 
    -0.0011830536043736519, -0.001439107602371297, -0.0016850506747929971, 
    -0.0019179966370974724, -0.0021345509563192003, -0.0023309338932358818, 
    -0.0025031781456964245, -0.0026473736718404675, -0.0027599648748115502, 
    -0.0028380467251184747, -0.0028796575641245022, -0.0028840456554872591, 
    -0.0028518634855102683, -0.0027853059404987081, -0.0026881422929196314, 
    -0.0025656517720731944, -0.0024244504643732485, -0.0022722017692478279, 
    -0.0021172351295066297, -0.001968072418216405, -0.0018328965117284178, 
    -0.0017189938849236435, -0.0016322328370027305, -0.0015765993027808849, 
    -0.0015538819167317647, -0.0015634984137389589, -0.0016025221101443456, 
    -0.0016658849260479294, -0.0017467641620577561, -0.001837100206881146, 
    -0.0019282177848001906, -0.0020114664343665795, -0.0020788292638966956, 
    -0.0021234431469639111, -0.0021399671161266695, -0.0021247915611907003, 
    -0.0020760946567220497, -0.0019937637372994276, -0.0018792532079497644, 
    -0.001735398825412772, -0.001566206935030382, -0.0013766297933659251, 
    -0.0011723185194612358, -0.00095935681747043495, -0.00074397552727740134, 
    -0.00053226341409935338, -0.00032989745474031404, 
    -0.00014191033425150972, 2.7503223773647931e-05, 0.00017511289636205682, 
    0.00029873362067045348, 0.00039725714786753298, 0.00047064166272521932, 
    0.00051986800324065204, 0.00054683671573272188, 0.00055423325632189991, 
    0.00054534346069237585, 0.00052383111832508638, 0.00049348619060697726, 
    0.00045797933734784645, 0.00042062637952483361, 0.00038420257758975884, 
    0.0003508071269708606, 0.00032181229929635836, 0.00029787591062823831, 
    0.0002790274101186799, 0.00026481178626215613, 0.000254469467578729, 
    0.00024713387135357232, 0.00024203260607450863, 0.00023865316178772422, 
    0.00023685941786793669, 0.00023693654703958896, 0.00023956001277113155, 
    0.0002456793933812623, 0.00025634667638425152, 0.00027252464734008042, 
    0.00029489634085019584, 0.00032370259968884279, 0.00035863823829694814, 
    0.00039878826746440161, 0.00044262576989733619, 0.00048804193179439456, 
    0.00053241908830638565, 0.00057273605089305443, 0.00060569498409073158, 
    0.00062787603452825968, 0.00063590097912401766, 0.00062661428339592766, 
    0.00059725503591029155, 0.00054562365476335483, 0.00047021269215097078, 
    0.00037031785306646144, 0.00024609432518698615, 9.8584779924288499e-05, 
    -7.0288081841417082e-05, -0.00025774768800285977, 
    -0.00046021417677540526, -0.00067337575052218686, 
    -0.00089228534929174715, -0.0011114937692136239, -0.0013252330247199809, 
    -0.0015276490745752928, -0.0017130803237295907, -0.0018763777111898304, 
    -0.0020132265819925977, -0.0021204493129785037, -0.0021962438083809126, 
    -0.0022403166236110396, -0.002253886390508917, -0.0022395654603613495, 
    -0.0022011048165587622, -0.0021430530970264557, -0.0020703550199751798, 
    -0.0019879285378042147, -0.0019002692260519033, -0.0018111147819261503, 
    -0.0017232066683065901, -0.0016381547064828819, -0.0015564160785467892, 
    -0.0014773684090975518, -0.0013994676133839827, -0.0013204592255764121, 
    -0.0012376321779754376, -0.0011480729347720152, -0.0010489272428399379, 
    -0.0009376137530678866, -0.00081200706470902851, -0.00067057921633238335, 
    -0.00051247907994546717, -0.00033755259724768324, 
    -0.00014630924668724871, 6.0173428795104466e-05, 0.00028038221646783408, 
    0.00051251840131217175, 0.00075465109341990892, 0.0010048546324739475, 
    0.0012613114468146157, 0.0015223799300627414, 0.0017866336269324247, 
    0.00205286266025548, 0.002320035162681804, 0.0025872484549716969, 
    0.0028536477397690272, 0.003118311831750268, 0.0033801423096665368, 
    0.0036377241401218687, 0.0038892169232256457, 0.0041322852446029068, 
    0.0043640734839598665, 0.0045812707406648881, 0.0047802232819339069, 
    0.0049571334926187035, 0.0051082705458508054, 0.005230213505045731, 
    0.0053200735685866411, 0.005375676104235433, 0.0053956886112992682, 
    0.0053796984249949243, 0.0053282144974152344, 0.0052426287009034985, 
    0.0051251442558394528, 0.0049786806847850733, 0.0048067679010227989, 
    0.0046134429398616431, 0.004403142280998135, 0.0041805841968985185, 
    0.0039506408813762611, 0.0037181976040979335, 0.0034879932928038862, 
    0.0032644586298278384, 0.0030515566050356596, 0.0028526436969446532, 
    0.0026703629039491316, 0.0025065850836853733, 0.0023623963372858187, 
    0.0022381515548380538, 0.0021335686696497625, 0.0020478856413169142, 
    0.0019800359883207731, 0.0019288589125585054, 0.0018932721109489168, 
    0.0018724241714967666, 0.001865775857151118, 0.0018731029512724154, 
    0.001894436678842371, 0.0019299216064145499, 0.0019796595374098704, 
    0.0020435250204327675, 0.0021210182292385727, 0.0022111517292371266, 
    0.0023124069572467063, 0.0024227531190428443, 0.002539739112641954, 
    0.0026606276423314515, 0.0027825659250416373, 0.0029027774457428112, 
    0.0030187264421178079, 0.0031282709117914221, 0.0032297631091828417, 
    0.0033221076214065559, 0.003404744025065526, 0.003477597156277947, 
    0.003540958642288458, 0.0035953254449334724, 0.0036412088339371545, 
    0.0036789186354721001, 0.0037083666927826674, 0.0037289101909992761, 
    0.0037392688792156179, 0.0037375199193559511, 0.0037212036077689764, 
    0.0036874894951063305, 0.0036334207942594421, 0.0035561744760395052, 
    0.0034533396568537027, 0.003323160232742409, 0.0031647218176577702, 
    0.0029780877659123734, 0.0027643444404451866, 0.0025255650913157341, 
    0.0022647177368259499, 0.0019854979726343985, 0.0016921324396146614, 
    0.0013891389743488341, 0.001081097713864831, 0.0007724170720397089, 
    0.00046711695528534064, 0.00016863928289952886, -0.0001203080624224956, 
    -0.00039785115274978007, -0.00066298848094364319, 
    -0.00091556309418271511, -0.0011561736517886004, -0.0013860283414073569, 
    -0.0016067634256011116, -0.0018202421033692369, -0.0020283377486882137, 
    -0.002232734849573384, -0.0024347343699367909, -0.0026350864401127314, 
    -0.0028338455281875963, -0.0030302509355462546, -0.0032226594884105469, 
    -0.0034085081141272907, -0.0035843556392052361, -0.0037459847083345494, 
    -0.0038885861948041479, -0.0040070120922226895, -0.0040960687830497895, 
    -0.0041508536683737083, -0.0041670718636046614, -0.0041413226562216597, 
    -0.0040713304734202004, -0.0039560800052363763, -0.0037958896234242625, 
    -0.0035924073805561163, -0.0033485412554415173, -0.0030683625544365364, 
    -0.0027569658907811039, -0.0024203164608030425, -0.0020650711840720574, 
    -0.0016984027223432871, -0.001327808510993661, -0.00096092099797264363, 
    -0.00060534444970764684, -0.00026847092100535687, 4.2678529251594861e-05, 
    0.00032163420688807314, 0.00056263766321226088, 0.00076081253781514228, 
    0.00091231829625199154, 0.0010144905847461676, 0.0010659493814290369, 
    0.0010666680616188387, 0.001018023890534843, 0.00092279248452007854, 
    0.00078510090836409407, 0.00061032257250086394, 0.00040489624972326585, 
    0.00017611028190088948, -6.8181942314950018e-05, -0.00031987072489433074, 
    -0.00057092533168320977, -0.00081373329827848185, -0.0010414164907784455, 
    -0.0012480993724889803, -0.0014291131597802158, -0.0015810765029724567, 
    -0.0017019095928061758, -0.0017907377018308651, -0.0018477326441973768, 
    -0.0018739228258843302, -0.0018709752757137669, -0.0018410063472305944, 
    -0.0017864015948375635, -0.0017096632863762924, -0.0016132750606660268, 
    -0.0014996067525321912, -0.0013708452569805936, -0.0012289669142414971, 
    -0.0010757632889968852, -0.00091290044834018726, -0.00074201376407391137, 
    -0.00056479543974645907, -0.00038306410418612361, 
    -0.00019879585970282372, -1.4120389602816084e-05, 0.00016873843180666728, 
    0.00034753634534548719, 0.00052012172703894957, 0.00068455083298449672, 
    0.00083920754834479071, 0.00098290368560017042, 0.0011149292212112242, 
    0.0012350652659540941, 0.0013435463488100893, 0.0014409620705286817, 
    0.0015281253174951211, 0.0016059141521296593, 0.0016751139112533865, 
    0.001736278365279701, 0.0017896332248295264, 0.0018349978132029391, 
    0.0018717734751654404, 0.0018989511420051683, 0.0019151430905962042, 
    0.0019186538570195705, 0.0019075558993020679, 0.0018798005657759201, 
    0.0018333481082625815, 0.0017663163121633394, 0.0016771271681276009, 
    0.0015646485474725992, 0.0014282875657930648, 0.0012680770751755709, 
    0.0010846998721875615, 0.00087951223140710815, 0.00065452052502900141, 
    0.0004123213938788378, 0.00015598284357190055, -0.00011112206753277715, 
    -0.00038551276117970837, -0.00066380593019093107, 
    -0.00094289559496697328, -0.0012200384151492029, -0.0014928866161327257, 
    -0.0017594364116589932, -0.002017949974842581, -0.0022668871276845574, 
    -0.0025048783852430079, -0.0027307227124118471, -0.0029434600634331981, 
    -0.0031424427574879778, -0.0033274604420505103, -0.003498867052218075, 
    -0.003657719774263879, -0.0038058697590368199, -0.0039459929588369479, 
    -0.0040815287279899861, -0.0042164987404346033, -0.0043552226246889895, 
    -0.0045019632367003905, -0.0046605232110419224, -0.0048338524524210507, 
    -0.0050237070424543218, -0.0052304072433189217, -0.005452720872055312, 
    -0.0056878889744624633, -0.0059317767780258891, -0.0061791319316617643, 
    -0.0064239360511031849, -0.0066597988044097946, -0.0068803760564825987, 
    -0.0070798015626499277, -0.0072530874852881318, -0.0073964836854642658, 
    -0.0075077537378741939, -0.0075863530702912386, -0.0076334746349739505, 
    -0.0076519595559664247, -0.0076460434234739442, -0.0076209699313403738, 
    -0.0075825035245628671, -0.0075363895952772755, -0.0074878242417520885, 
    -0.0074410135086972178, -0.0073988652625788277, -0.0073628507585068517, 
    -0.0073330212156443551, -0.007308190830643168, -0.0072862285543275904, 
    -0.0072644321378944445, -0.0072399227210283891, -0.0072100160663650659, 
    -0.0071725604229648391, -0.0071261660966211553, -0.0070703556766314709, 
    -0.0070055876061587844, -0.006933172967205462, -0.0068550843553592039, 
    -0.0067736657579204685, -0.0066912897806388223, -0.00660997616173603, 
    -0.0065310636202131466, -0.0064549669594534927, -0.0063811154153016218, 
    -0.006308056614559578, -0.0062336928905301972, -0.0061556037316843797, 
    -0.0060713734054431033, -0.0059788930189843921, -0.0058765865815415437, 
    -0.0057635795435685699, -0.0056397658038664479, -0.0055057907070334136, 
    -0.0053629447664217678, -0.005212980735774273, -0.0050578822870079978, 
    -0.0048995951113090883, -0.0047398098324515584, -0.0045797877903502853, 
    -0.0044202801948663335, -0.0042615551494716098, -0.0041035040761450521, 
    -0.0039458146930077482, -0.0037881515084295103, -0.0036303203284706411, 
    -0.0034723786016343699, -0.0033146723269495484, -0.0031578253201479758, 
    -0.0030026801565952352, -0.0028502191396558734, -0.0027014968238506204, 
    -0.0025575561974618376, -0.0024193687215645666, -0.002287767416688269, 
    -0.0021634112158153318, -0.0020467458160666613, -0.0019379963984597986, 
    -0.0018371598152689304, -0.0017440300411658131, -0.0016582012302457829, 
    -0.0015790923213494566, -0.0015059463364407476, -0.0014378195580112192, 
    -0.0013735610382426364, -0.0013117983645332908, -0.0012509274949161935, 
    -0.0011891311575593251, -0.0011244320230290208, -0.0010547846819942196, 
    -0.00097818412936658754, -0.0008928049306888749, -0.00079712402725433396, 
    -0.00069004234213544777, -0.00057098825281013928, 
    -0.00044000079565416393, -0.00029777447527215301, 
    -0.00014569971148659585, 1.415306895611175e-05, 0.00017906088725334733, 
    0.00034572032455174457, 0.00051034513311272174, 0.00066878486884055339, 
    0.00081665510569868267, 0.00094947214422021686, 0.0010627619410349112, 
    0.001152160150784618, 0.0012135015227190602, 0.0012428927887620108, 
    0.0012368089535643796, 0.001192201867503709, 0.0011067023813404694, 
    0.00097884758665961078, 0.00080836883404967759, 0.0005964598458292579, 
    0.00034600021302578495, 6.1661989919010294e-05, -0.00025011879817814908, 
    -0.00058131555504378231, -0.00092263579828311018, -0.0012639887225063132, 
    -0.0015950348318768343, -0.0019058108276443627, -0.0021873711602881365, 
    -0.0024323427122706913, -0.0026353580352698842, -0.0027932975784355045, 
    -0.0029052776449554028, -0.0029724600021161628, -0.0029976923452031362, 
    -0.0029850961520369373, -0.0029396384204878443, -0.0028667621648870109, 
    -0.0027720409553494947, -0.0026608762121324396, -0.0025381639007382205, 
    -0.0024079620602160375, -0.0022732012718112934, -0.0021355097510533123, 
    -0.0019952221376719819, -0.0018515440390011219, -0.0017028655480218458, 
    -0.0015471585448166957, -0.0013824274037473568, -0.0012071491593439584, 
    -0.0010206726760610824, -0.00082351983569706232, -0.00061757307831777257, 
    -0.00040610236930560306, -0.00019364708546713567, 1.4222063131733113e-05, 
    0.00021124272336754107, 0.00039085333426960698, 0.00054659580341758515, 
    0.00067253508839210704, 0.00076364175075101736, 0.00081614600446618091, 
    0.00082782930979003648, 0.00079823325784575926, 0.00072875813473667291, 
    0.00062264522675909773, 0.00048484922505185007, 0.00032178539496701238, 
    0.00014099421284942789, -4.925018422454935e-05, -0.00024036487529227751, 
    -0.00042386714277834673, -0.00059175998153522731, 
    -0.00073691075516806146, -0.00085335362178697244, 
    -0.00093653169037999893, -0.00098346420347053716, 
    -0.00099278321939300692, -0.00096468303584093843, -0.0009007668869700393, 
    -0.00080381773995837384, -0.00067753878538531613, -0.0005262794337320462, 
    -0.00035475986047531829, -0.00016781377754070036, 2.9841857459769689e-05, 
    0.00023382031912194367, 0.00044023881619712559, 0.00064589314774174194, 
    0.00084835113784079196, 0.0010460616869214319, 0.0012383629976909728, 
    0.0014254474490929814, 0.001608278997114065, 0.0017884290122300787, 
    0.0019678741130762819, 0.0021487603816915078, 0.0023331545525619875, 
    0.0025227899334810898, 0.0027188438584030204, 0.0029217452294945955, 
    0.0031310316802622981, 0.0033452557461599421, 0.003561944891485834, 
    0.0037776165985721716, 0.0039878620270740028, 0.0041874838472629955, 
    0.0043707161660375832, 0.0045314625942841445, 0.0046635500278956361, 
    0.004760938070806439, 0.0048178832615970646, 0.004829036475631536, 
    0.0047895256224253788, 0.0046950440238453343, 0.0045420438793983432, 
    0.0043279877693383267, 0.0040516484107223317, 0.0037134223614111658, 
    0.0033155065152416481, 0.0028619659891603441, 0.0023586327747037593, 
    0.0018129160699689837, 0.0012335511288059451, 0.00063033064771968997, 
    1.3836773459843042e-05, -0.00060486854149045116, -0.0012145610675946875, 
    -0.0018041909010936539, -0.0023632163374473466, -0.0028819162845989885, 
    -0.0033516572285416995, -0.0037651251769580726, -0.004116479426605737, 
    -0.0044014740573273857, -0.0046175295739120477, -0.0047637914893777248, 
    -0.0048411689052716492, -0.0048523248546279291, -0.0048016475852521757, 
    -0.004695130034194985, -0.0045402074934991401, -0.0043455108068244166, 
    -0.0041205622057561677, -0.0038754559927866666, -0.0036204666635823498, 
    -0.0033656884654975393, -0.0031206735891476209, -0.0028940964001706363, 
    -0.0026934804681503837, -0.0025249857295230652, -0.0023932401291316308, 
    -0.0023012534330977743, -0.0022503709895235631, -0.0022402834909898972, 
    -0.0022691136279363272, -0.0023335395985961392, -0.0024289830785653066, 
    -0.0025498091730796419, -0.0026895755828772396, -0.0028413252233069333, 
    -0.0029979179890018827, -0.0031523546676238455, -0.0032981241338083272, 
    -0.003429486194517252, -0.003541683622066358, -0.0036310797958214731, 
    -0.0036951561931432078, -0.0037324262261178342, -0.003742238294708787, 
    -0.0037245382245637238, -0.0036795883989980188, -0.0036077340082313397, 
    -0.0035092123579327406, -0.0033840566672295579, -0.0032320664398662454, 
    -0.0030528784539760718, -0.0028460986842141524, -0.0026114876600397707, 
    -0.0023491543354986029, -0.0020597555604798044, -0.0017446718808580999, 
    -0.0014061302998396325, -0.0010472758883336448, -0.00067213626075236072, 
    -0.00028546455334690999, 0.00010754199245115711, 0.00050163363940536158, 
    0.00089195541127866623, 0.0012744990478766659, 0.001646421480169353, 
    0.0020062595494735411, 0.0023538974877858228, 0.002690388707761642, 
    0.0030175835245526248, 0.0033377107411316216, 0.0036529478821002168, 
    0.0039650018084345998, 0.0042747838473524372, 0.0045821755601801401, 
    0.0048858700421265397, 0.0051833233862488802, 0.0054707540302894068, 
    0.0057432457547936158, 0.0059948870434157935, 0.0062189940140090884, 
    0.0064083776650023889, 0.0065557016099622263, 0.0066537851454180211, 
    0.0066959791424732844, 0.0066764965636653267, 0.0065906484892868256, 
    0.0064350810854495412, 0.0062079108112064281, 0.0059087915713829453, 
    0.005538977020185405, 0.0051012923870901684, 0.0046001319119429685, 
    0.004041425991009622, 0.0034325512016877596, 0.0027822101667394615, 
    0.0021001780360042745, 0.0013969689103019243, 0.00068342006082707408, 
    -2.970180113117632e-05, -0.00073211769068458159, -0.0014143438806290404, 
    -0.0020679064894505595, -0.0026854741753005932, -0.0032608739312435121, 
    -0.0037889953220374803, -0.0042656593821690124, -0.004687476170567197, 
    -0.0050516877027970263, -0.0053561043108521292, -0.0055990689788522202, 
    -0.0057795430911761611, -0.0058972241928100001, -0.0059526834221908173, 
    -0.0059475111686797654, -0.0058843535509284887, -0.0057668466899199709, 
    -0.0055994646550684693, -0.0053872521678403375, -0.0051355258962411327, 
    -0.0048496197539639151, -0.004534663389332695, -0.0041954609481795226, 
    -0.0038364297012015241, -0.0034615913508963757, -0.0030745665318255276, 
    -0.0026785317724472035, -0.0022761542690074989, -0.0018694486891943614, 
    -0.0014596471316719994, -0.0010470358409994777, -0.00063082614882709368, 
    -0.00020909920285590308, 0.00022118040005889169, 0.00066401819802730663, 
    0.0011241162125128919, 0.0016064879775181619, 0.0021159577601332414, 
    0.0026565779134109409, 0.0032310511686013924, 0.003840226956472802, 
    0.004482753000452761, 0.0051549014209046271, 0.0058506334124702785, 
    0.0065618078441257444, 0.0072785010298037313, 0.0079894455042632245, 
    0.0086825023810247169, 0.0093451693377007913, 0.0099651285364339062, 
    0.010530787235295921, 0.011031818341141147, 0.011459624188367171, 
    0.011807742861682869, 0.012072110719041008, 0.012251190463873834, 
    0.012345925439390228, 0.012359565376912634, 0.012297347330903187, 
    0.012166087194156128, 0.011973766529369122, 0.011729075887409846, 
    0.011441044547416812, 0.011118743404524328, 0.010771083195806285, 
    0.010406696591704959, 0.01003384140345142, 0.0096603414038571467, 
    0.0092935185927486997, 0.0089400948192536051, 0.0086060738525473544, 
    0.0082965936230998578, 0.0080157575447165497, 0.0077664439174676865, 
    0.0075501941307007684, 0.0073670620829020123, 0.007215608243450162, 
    0.0070929173124121281, 0.0069947017749417036, 0.0069154996008688203, 
    0.006848917135180814, 0.0067879033518185913, 0.0067250408124154204, 
    0.0066527836515230341, 0.0065636779199439964, 0.0064504770650855364, 
    0.0063062455023201762, 0.0061244493032832741, 0.0058990682919929684, 
    0.0056247175639188452, 0.0052968345276443373, 0.0049118476054103542, 
    0.0044673027077955021, 0.0039620607937633822, 0.0033963981976657363, 
    0.0027721504926529351, 0.002092871068699897, 0.0013639336061644905, 
    0.00059266596179385444, -0.00021160299839199895, -0.001037647510893424, 
    -0.0018726691044173198, -0.0027027706831166155, -0.0035136777264642969, 
    -0.0042915351811168151, -0.0050237026867782321, -0.0056994047124299136, 
    -0.006310222996456733, -0.0068502739599816606, -0.0073161389828412995, 
    -0.0077065410908659406, -0.008021879117051477, -0.0082636458857541801, 
    -0.0084338388435823645, -0.0085344812062657701, -0.0085672445528147227, 
    -0.0085332356280128762, -0.0084329373888817078, -0.0082663345267921153, 
    -0.0080331466640919877, -0.0077331961650234969, -0.0073668051727638377, 
    -0.0069352322003122056, -0.0064410828835917509, -0.0058886118700366141, 
    -0.00528395914292257, -0.0046351798793851833, -0.0039521550696142811, 
    -0.0032463098502782863, -0.0025302745350521136, -0.0018174353967774905, 
    -0.0011214958790179616, -0.00045596273514629868, 0.00016629154721258788, 
    0.00073347337194381288, 0.0012352392026167812, 0.001662963087303262, 
    0.002009897995832401, 0.0022712613687022429, 0.0024441546975183148, 
    0.0025274465322979865, 0.0025215418250998578, 0.0024281719602251947, 
    0.0022501654454019845, 0.0019912542191790864, 0.0016559312991150112, 
    0.0012493473289534693, 0.0007772864960165504, 0.0002462115685020553, 
    -0.0003366796312886283, -0.0009633460250137785, -0.0016248202747193993, 
    -0.0023110943149431042, -0.0030110694150389454, -0.0037125066531641824, 
    -0.0044020901613955931, -0.0050655762665919434, -0.0056880775848655819, 
    -0.0062544903002174799, -0.0067500339768712505, -0.007160910693145367, 
    -0.0074749258267447225, -0.0076821814570623686, -0.0077756648728523675, 
    -0.007751743863312577, -0.0076106017171238653, -0.0073564726069366149, 
    -0.0069978011200429466, -0.006547183624604198, -0.0060210818210330473, 
    -0.0054392746504763698, -0.0048239728152623023, -0.0041985712896085037, 
    -0.0035862782823096362, -0.0030086655496751658, -0.002484490046416482, 
    -0.0020289866935638474, -0.0016537721965194428, -0.0013671286734984345, 
    -0.0011743907077636777, -0.0010780939955039293, -0.0010776860839190232, 
    -0.0011690525985217325, -0.0013441607086126948, -0.0015911814666975648, 
    -0.0018951637936112271, -0.0022391564292225455, -0.0026055242828298261, 
    -0.0029771910408258151, -0.0033385774094684406, -0.0036761152395738688, 
    -0.0039784924807758715, -0.0042366011887430563, -0.0044435239732534305, 
    -0.0045944488957519224, -0.0046866786760875112, -0.0047195360942560664, 
    -0.0046942272268537741, -0.0046136008189087939, -0.0044818140347559409, 
    -0.0043040411136506989, -0.0040861675300643977, -0.0038346944983178961, 
    -0.003556606159329435, -0.0032593603674628967, -0.0029507426879236665, 
    -0.0026386796750954679, -0.0023308300072799192, -0.0020341328055185114, 
    -0.0017541966506247721, -0.0014947498256473739, -0.0012572648157335826, 
    -0.001040678524926351, -0.00084149173758484908, -0.00065407058417980401, 
    -0.00047115098530703734, -0.00028451088199050886, 
    -8.5676560809795844e-05, 0.00013342535141284471, 0.00037991390574791765, 
    0.00065956842164051495, 0.0009765774316212103, 0.0013334275780244283, 
    0.0017308357863728763, 0.0021676918733216262, 0.0026409270221462674, 
    0.0031454933612776355, 0.0036743905767765935, 0.0042188654019771508, 
    0.0047688187807689133, 0.0053132837090594312, 0.0058409329502495866, 
    0.0063405886687688817, 0.0068016412020745279, 0.0072145376599934497, 
    0.0075711548850201293, 0.0078652539611147373, 0.0080928050621331508, 
    0.0082522198754705553, 0.0083445028959721005, 0.0083732180148069942, 
    0.008344263275784471, 0.0082655510989509181, 0.0081465175525489014, 
    0.0079976324956716055, 0.0078299283811402876, 0.0076545889734321356, 
    0.0074826385837749457, 0.0073247852374340857, 0.0071913179839710184, 
    0.0070920109720540928, 0.0070359936583165713, 0.0070315039673562148, 
    0.0070856462134759341, 0.0072040856115050513, 0.0073908242611501656, 
    0.0076480000509379972, 0.0079758784531700471, 0.0083728808215511579, 
    0.0088357661769487075, 0.0093597676884680289, 0.0099388892829705665, 
    0.010566024211068397, 0.011233087476590003, 0.011931061170746007, 
    0.012650048789461068, 0.013379299356926971, 0.01410732143591217, 
    0.014822137701934524, 0.01551166542225345, 0.016164180952548127, 
    0.016768754878477388, 0.017315887531529846, 0.017798038174534167, 
    0.018209991016628343, 0.018549233061971912, 0.018816366117697866, 
    0.019015204252981772, 0.019152855658073776, 0.019239613833723739, 
    0.019288609224799153, 0.019315324459775983, 0.019337004036750587, 
    0.019371995705083703, 0.019438861420476451, 0.019555420094360808, 
    0.019737409413463886, 0.019997220181287762, 0.020342568859830643, 
    0.020775554648212156, 0.021291996665163928, 0.021881381109356914, 
    0.022527305126986814, 0.023208370537712249, 0.023899396852223725, 
    0.024572633826624824, 0.025199041513890859, 0.025749486259793512, 
    0.026195574675308957, 0.026510740948835189, 0.026671155876679276, 
    0.026656585725472949, 0.0264514290803664, 0.026045597183309888, 
    0.025435352432726498, 0.02462420508271539, 0.023623451436595343, 
    0.022452632076239851, 0.02113947695100523, 0.019719126633777902, 
    0.018233005568496614, 0.016726739027685424, 0.015247556414400225, 
    0.013841453035448826, 0.012550200151438349, 0.011408428203242246, 
    0.010441155196341825, 0.0096617160329938376, 0.0090704174463809416, 
    0.0086543278612443361, 0.0083874701238863796, 0.008232508496586884, 
    0.0081430815590580585, 0.0080669913759500965, 0.0079499740028854595, 
    0.0077398423938152367, 0.0073904722465231686, 0.0068661778457640259, 
    0.0061448042211492875, 0.0052207617678664813, 0.0041065296494993356, 
    0.0028323530075566568, 0.0014441470069617337, -5.1363982805202529e-07, 
    -0.0014377250969025428, -0.0028041599470061749, -0.0040430532585009806, 
    -0.0051085735915532785, -0.0059689214265544821, -0.0066058285999857332, 
    -0.007014247051489661, -0.0072002249855703622, -0.0071782365971705389, 
    -0.0069713701375117253,
  // Fqt-total(7, 0-1999)
    0.99999999999999956, 0.99388909793499147, 0.97581459531923176, 
    0.94652877848077477, 0.90721850598674914, 0.85941532857128466, 
    0.80488524799822769, 0.74551032402294981, 0.68317393706644858, 
    0.61965967322392779, 0.55657087891804147, 0.49527457381347939, 
    0.43687028229180452, 0.3821817492960432, 0.33176762687712047, 
    0.285946339562826, 0.24483006737799398, 0.2083632067160773, 
    0.17636139886247373, 0.14854828223574512, 0.12458798553624788, 
    0.1041123716818456, 0.08674271975144017, 0.072106076599414828, 
    0.059846874198045019, 0.049634523012996187, 0.041167774198654548, 
    0.034176616196248628, 0.028422371994221228, 0.02369660168292103, 
    0.019819251457524067, 0.016636384559235717, 0.014017739823380108, 
    0.011854215980410227, 0.010055390806292801, 0.0085471056112393206, 
    0.0072691657051733695, 0.0061732022826394128, 0.0052207270060710808, 
    0.0043814334592283061, 0.0036317290794939689, 0.00295350895162716, 
    0.0023331228334842196, 0.0017605059024657335, 0.0012284323832185333, 
    0.00073185016814792455, 0.00026729531417032481, -0.00016763487989921146, 
    -0.00057472949189144669, -0.00095554121270399761, -0.0013116537884334649, 
    -0.0016448397258691471, -0.0019571044747051739, -0.0022506283744741784, 
    -0.0025276258795873755, -0.002790174367515056, -0.0030400420179265723, 
    -0.0032785603230876068, -0.0035065813533217975, -0.0037245143392859088, 
    -0.0039324528351342425, -0.0041303475044927119, -0.0043182033942985049, 
    -0.004496233424714737, -0.0046649717113097554, -0.004825273195970951, 
    -0.0049782519575408673, -0.0051251207085965577, -0.005266996870467648, 
    -0.0054046966325759088, -0.0055385596429185398, -0.0056683284458535835, 
    -0.0057930986661184547, -0.0059113156808066501, -0.0060208153089788873, 
    -0.0061188817361879366, -0.0062023143163195413, -0.006267503093351035, 
    -0.0063105140275633116, -0.0063272074751140545, -0.006313383618257209, 
    -0.0062649877770439687, -0.0061783417814332865, -0.0060504181841735775, 
    -0.0058791208773191503, -0.0056635564400094283, -0.0054042592867070043, 
    -0.0051033703473651847, -0.0047647361215818066, -0.0043939119406402136, 
    -0.0039980805333802907, -0.0035858638022569262, -0.0031670532432766562, 
    -0.0027522671097984543, -0.0023525550006655476, -0.0019789648498089864, 
    -0.0016421038728728862, -0.0013517072124663487, -0.0011162475049381632, 
    -0.0009426038892824106, -0.00083580799289199826, -0.00079889628606316968, 
    -0.00083285693352401035, -0.00093667668551467649, -0.0011074687531448225, 
    -0.0013406565349847548, -0.0016301956530566089, -0.0019687963242973577, 
    -0.0023481364423281253, -0.0027590483595052169, -0.0031916881905975905, 
    -0.0036356861975783052, -0.0040802980501501301, -0.0045145918294141911, 
    -0.0049276511644251262, -0.0053088460821392588, -0.0056481361475358861, 
    -0.0059364221591163471, -0.0061658973353197468, -0.0063303915904141753, 
    -0.0064256466494790219, -0.0064494929039651521, -0.0064018991569344845, 
    -0.0062848699070467626, -0.0061021935511945159, -0.0058590956271823823, 
    -0.0055618166979624342, -0.0052172014522505672, -0.0048323442087808751, 
    -0.004414332026297034, -0.0039701030708832559, -0.003506417895688074, 
    -0.0030299018401694091, -0.0025471451346624537, -0.0020647976238211663, 
    -0.0015896555228868759, -0.0011287018836643584, -0.00068908086634383034, 
    -0.00027802174067683908, 9.7299434557271126e-05, 0.00042996046906490937, 
    0.00071351375861546465, 0.00094224687930633975, 0.0011114375557505624, 
    0.0012175902240053966, 0.0012586273474148658, 0.0012340255728255788, 
    0.0011448587085857455, 0.00099376934833205876, 0.00078486459047220902, 
    0.0005235464352139048, 0.00021630673561687653, -0.0001295073816716437, 
    -0.00050594804765572571, -0.00090471765681540738, -0.0013174252596140235, 
    -0.0017358164824683091, -0.0021519870086845493, -0.0025585577353867076, 
    -0.0029488280479449207, -0.0033169052579726781, -0.0036578231058809869, 
    -0.0039676271674450054, -0.0042434372906194383, -0.0044834385732138394, 
    -0.0046868226198668508, -0.0048536701179931535, -0.0049848089184143726, 
    -0.005081634289770506, -0.0051459242798084807, -0.0051796331950340092, 
    -0.0051847044293178305, -0.0051629237948354091, -0.005115829978962357, 
    -0.0050447166348797428, -0.0049507134958702683, -0.0048349327071031938, 
    -0.0046986546918937264, -0.0045435163094085856, -0.0043716575422640975, 
    -0.0041858040577103977, -0.0039892460403358832, -0.0037857237723091883, 
    -0.0035792089139621004, -0.0033736362794952192, -0.0031726035744718854, 
    -0.0029790993208858871, -0.0027952998716779314, -0.0026224596182437025, 
    -0.0024609074739767763, -0.0023101486631430055, -0.0021690468565622001, 
    -0.0020360499773657546, -0.0019094440594077332, -0.0017875734193857724, 
    -0.0016690243892812037, -0.0015527370724671124, -0.0014380396786086659, 
    -0.0013246150953750942, -0.0012124015456313037, -0.0011014673652447226, 
    -0.00099188238367804563, -0.0008836254337857511, -0.00077654360199337039, 
    -0.00067037285828869589, -0.00056482648212201141, 
    -0.00045970848194705298, -0.00035504502960862486, 
    -0.00025119347862645995, -0.00014889662172380957, 
    -4.9279446031279992e-05, 4.6233211923624336e-05, 0.00013605935811254128, 
    0.00021865343062892252, 0.0002927228731407867, 0.00035743943538861533, 
    0.00041261880033505941, 0.00045884478606303218, 0.00049751710098061596, 
    0.00053080535313996115, 0.00056153815987400465, 0.00059300378448255166, 
    0.00062871257608111198, 0.00067213687052751785, 0.00072644953115953833, 
    0.00079431168900360972, 0.00087771020660887213, 0.00097786637752617718, 
    0.0010952161134828034, 0.0012294454555931659, 0.0013795610850738393, 
    0.0015439705830916574, 0.0017205406336650239, 0.0019066243647290874, 
    0.0020990372525710854, 0.0022940010379285136, 0.0024870689222641134, 
    0.0026730586012953224, 0.0028460331816727805, 0.0029993660494722872, 
    0.0031259097626965358, 0.003218282699987327, 0.0032692601559964132, 
    0.0032722391451743787, 0.0032217257630022165, 0.0031137991479968496, 
    0.0029464876966296292, 0.0027200242216570626, 0.0024369465902121189, 
    0.0021020421926609004, 0.0017221570492048275, 0.0013058776441707493, 
    0.00086313031118844354, 0.00040471527107379686, -5.819735935661662e-05, 
    -0.00051458030532555504, -0.0009540356024616435, -0.0013672302259927281, 
    -0.0017462268587280416, -0.0020846932801462238, -0.0023779697660072812, 
    -0.0026230011620553832, -0.0028181561224342069, -0.0029629983974267505, 
    -0.0030580384722525408, -0.0031045229544529587, -0.0031042767808152258, 
    -0.0030595882552085759, -0.0029731571753330798, -0.0028480605590136916, 
    -0.0026877445470663243, -0.0024960155129853325, -0.0022770391092763105, 
    -0.0020353146639296793, -0.0017756397227540255, -0.001503037573858245, 
    -0.0012226594633403479, -0.00093965644105628674, -0.00065902421428613812, 
    -0.00038544570108788224, -0.00012313123248748796, 0.00012430742139773036, 
    0.00035396073396122595, 0.00056367062397177546, 0.00075203841039883342, 
    0.00091839421654716605, 0.0010627318297185306, 0.0011856321232691339, 
    0.0012881824022350676, 0.0013719054253156266, 0.0014387013442972866, 
    0.0014908067754251808, 0.0015307601686781454, 0.0015613666403527066, 
    0.0015856410564333745, 0.0016067269352718972, 0.0016277753856907562, 
    0.0016517893163146852, 0.0016814309629858445, 0.0017188225942859185, 
    0.0017653506490724127, 0.0018215019687935479, 0.0018867430574662396, 
    0.001959476775520665, 0.0020370650332926783, 0.0021159305909735351, 
    0.0021917124146655065, 0.0022594835643700009, 0.002314007151533193, 
    0.0023500227156301179, 0.002362553421561608, 0.002347217823966425, 
    0.0023005108837625219, 0.0022200377648508548, 0.0021046765504778419, 
    0.001954654285644676, 0.0017715409247681954, 0.0015581911673019197, 
    0.0013186305874455357, 0.0010579270983932386, 0.00078203624449012135, 
    0.00049761675840995505, 0.00021180791742659923, -6.803965905773321e-05, 
    -0.0003346602298779206, -0.00058118092946087658, -0.000801392286503308, 
    -0.00098996031546951468, -0.0011425622931467265, -0.0012559462627982514, 
    -0.0013279345561384814, -0.001357389131447231, -0.0013441672851473563, 
    -0.0012890601455463992, -0.0011937293013877524, -0.0010606248218447431, 
    -0.00089288119649671277, -0.00069420867213075652, 
    -0.00046877929158200502, -0.00022112735893444488, 4.3954113939781112e-05, 
    0.00032149762428482817, 0.00060644213294883088, 0.00089371845149898343, 
    0.0011783197621180561, 0.0014553494735176989, 0.0017200513805110155, 
    0.0019678185678736818, 0.0021942029712759929, 0.0023949612718436025, 
    0.0025661527199041952, 0.002704296377859238, 0.0028065971658387794, 
    0.0028711805639915376, 0.002897296080654861, 0.0028854421474421121, 
    0.0028373581404514676, 0.0027558991653153916, 0.0026447798572685364, 
    0.0025082538118236771, 0.0023507402136199347, 0.0021764849012916991, 
    0.001989264604040713, 0.0017921782077633523, 0.001587539969426708, 
    0.0013768806577302787, 0.001161038396194379, 0.00094034341067064718, 
    0.00071487159232187954, 0.00048474557033860091, 0.00025043912925338797, 
    1.3062456147494174e-05, -0.00022543586217046017, -0.00046215930784618926, 
    -0.00069327969860002168, -0.0009141583085490975, -0.0011195555512867382, 
    -0.0013038933828027712, -0.0014615489969412314, -0.0015871638443455192, 
    -0.0016759491721562727, -0.0017239919778192293, -0.0017285380450750051, 
    -0.0016882519817119051, -0.0016034130479298913, -0.0014760259843006873, 
    -0.0013098265574179755, -0.0011101608633805743, -0.00088376803337969424, 
    -0.00063846388566569858, -0.00038277467779063303, 
    -0.00012554694298421551, 0.00012444342435888873, 0.00035886542506325661, 
    0.00057017202356416329, 0.00075189445111209757, 0.00089888349109122081, 
    0.0010074961575064845, 0.0010757159066895586, 0.0011032100818078824, 
    0.0010913036912992388, 0.0010428982252704488, 0.00096230844095191001, 
    0.00085504337317181278, 0.00072752911620550765, 0.00058677866636199394, 
    0.00044004024528961105, 0.00029443700980520297, 0.00015662535770199896, 
    3.2514675816729199e-05, -7.2944447435813265e-05, -0.00015586763006435623, 
    -0.00021345646944467042, -0.00024391547217618117, 
    -0.00024631554197909842, -0.00022042601935101506, 
    -0.00016654558912117341, -8.5382315459423208e-05, 2.2018664290605991e-05, 
    0.00015429751873426086, 0.00030975106451032268, 0.00048627895451687118, 
    0.00068133233474749013, 0.00089187077628981716, 0.0011143565785691292, 
    0.0013447881700694262, 0.0015787808322777551, 0.0018116774356037432, 
    0.0020386895866074104, 0.0022550426401046061, 0.0024561392280492574, 
    0.0026377060484559251, 0.0027959453437428235, 0.0029276612014471643, 
    0.003030382386509942, 0.0031024572851960997, 0.0031431358652011885, 
    0.0031526173233497488, 0.003132071340038246, 0.0030836174664894507, 
    0.0030102622590921315, 0.0029157801655254889, 0.0028045475581894908, 
    0.0026813202859112856, 0.0025509875795244477, 0.0024183324273679835, 
    0.0022877902017734535, 0.0021632715743763399, 0.002048021126072348, 
    0.0019445343249268159, 0.0018545138671382652, 0.0017788584645070434, 
    0.00171769274306626, 0.0016704456385388756, 0.0016359473083517959, 
    0.0016125214102552347, 0.0015980451886320162, 0.0015899855924051427, 
    0.0015854354832070482, 0.0015811994040226581, 0.0015739364108697082, 
    0.0015603698134284418, 0.0015375353227485328, 0.0015030064958679683, 
    0.0014550658189889881, 0.00139280009860015, 0.0013161001084948394, 
    0.0012255879847559421, 0.0011224842393299985, 0.0010084623091766605, 
    0.00088549058313991532, 0.00075568932470190331, 0.00062120427382318167, 
    0.00048409522566958678, 0.00034625464402388261, 0.00020934628820243328, 
    7.4763410571701395e-05, -5.6380779121950027e-05, -0.00018324853006339983, 
    -0.00030524914156313334, -0.00042199681636272888, 
    -0.00053325721675411344, -0.00063888273531933245, 
    -0.00073875511102343069, -0.00083271566530789215, -0.0009205155214518536, 
    -0.001001760254547482, -0.0010758629598081829, -0.0011420014009275432, 
    -0.0011990826575624346, -0.0012457351337598936, -0.0012803317352886091, 
    -0.0013010681480312303, -0.0013060833239289279, -0.0012936185645271326, 
    -0.0012621766593302014, -0.001210675669230528, -0.0011385495896912073, 
    -0.0010458099860324484, -0.00093305245942747325, -0.00080142682142133345, 
    -0.00065255713102508261, -0.00048845809210527956, 
    -0.00031141228217841671, -0.00012386281584522691, 7.1700625957111754e-05, 
    0.00027282705035804424, 0.00047715516648369157, 0.00068243120153305462, 
    0.00088647707424086616, 0.0010871597219839636, 0.0012823612100688873, 
    0.0014699861430939227, 0.0016480190420776948, 0.0018146089040901288, 
    0.0019681864455130403, 0.0021075691834574568, 0.0022320474862439917, 
    0.0023414348465959434, 0.0024360632281315128, 0.002516727002348004, 
    0.0025845746923880827, 0.0026409778802331638, 0.0026873693273946828, 
    0.002725098105343879, 0.0027553195314331748, 0.0027789385084095778, 
    0.0027966132262423754, 0.0028088230841436649, 0.0028159906894212501, 
    0.0028186165057810081, 0.0028174091435672287, 0.0028133658299256598, 
    0.002807775334071463, 0.0028021434353354508, 0.0027980461943851193, 
    0.0027969296989251578, 0.0027998974106627213, 0.0028075072754705777, 
    0.0028196047620294854, 0.0028352245497773277, 0.0028525476711791925, 
    0.002868927632811749, 0.0028809737629472356, 0.0028846843314123925, 
    0.0028756206326054174, 0.0028491382126511625, 0.0028006582653451843, 
    0.0027260037760195904, 0.0026217513589227833, 0.0024856014458343964, 
    0.002316714403363809, 0.0021159520286299412, 0.0018860117312047989, 
    0.0016314057757878353, 0.0013582938808439423, 0.0010741745671843652, 
    0.00078748844659675625, 0.00050716993475413078, 0.00024216507149086954, 
    9.5304159319603331e-07, -0.00020890522559099874, -0.0003811683002882104, 
    -0.00051121630169394358, -0.00059624843005903945, 
    -0.00063534796562718539, -0.00062943061700495683, 
    -0.00058106040626210002, -0.00049417481831655417, 
    -0.00037373073832865338, -0.00022530966236516522, 
    -5.4714519238118293e-05, 0.00013240038613590403, 0.00033084132501126639, 
    0.00053609618291624108, 0.00074445875037847825, 0.00095305030206380137, 
    0.0011597593986946491, 0.0013631137464512437, 0.0015621140790429014, 
    0.0017560666115935604, 0.0019444362320301383, 0.0021267274114513865, 
    0.0023024191061955909, 0.0024709349715772667, 0.002631637488296373, 
    0.0027838402233983472, 0.0029268201891556873, 0.0030598264364929371, 
    0.0031820713799346825, 0.0032927169131482014, 0.0033908407116925265, 
    0.0034753964950236089, 0.0035451805481627064, 0.0035988017545282988, 
    0.0036346719199013408, 0.0036510285335918154, 0.0036459822819876848, 
    0.0036176201774297287, 0.0035641322560240095, 0.0034839789611807851, 
    0.0033760884729128501, 0.0032400478755130733, 0.0030762818333218513, 
    0.0028861943968694157, 0.0026722423442961979, 0.0024379568667632005, 
    0.0021878801366947047, 0.0019274430394248523, 0.0016627766645180429, 
    0.0014004652051573686, 0.0011472568367291418, 0.00090972914945084012, 
    0.00069394934065995317, 0.00050512798500694739, 0.00034732488425337721, 
    0.0002232160773399745, 0.00013396273403499154, 7.9205158280590035e-05, 
    5.7175127926841179e-05, 6.492542886128781e-05, 9.8629320124416376e-05, 
    0.00015394188983042879, 0.00022632756959727512, 0.00031134971138257577, 
    0.00040487466475449331, 0.00050317667224312784, 0.00060297967406415791, 
    0.00070143129640509966, 0.00079604886601050294, 0.00088464065413794749, 
    0.00096525153464344354, 0.0010361252377286891, 0.0010957329345937729, 
    0.0011428588918967082, 0.0011767395089059519, 0.0011972302040810631, 
    0.0012049568967840078, 0.0012014227412876753, 0.0011890321267053981, 
    0.0011710249840658398, 0.0011513270648466068, 0.0011343226473608729, 
    0.0011245739735562528, 0.0011265138291616981, 0.0011441262762108618, 
    0.001180644001637335, 0.0012382844501863288, 0.0013180405833889562, 
    0.0014195272694034276, 0.0015409209672308773, 0.0016789855200117368, 
    0.001829186920077847, 0.0019859111530439802, 0.0021427675167063672, 
    0.0022929543581651363, 0.0024296728740988934, 0.0025465425892933257, 
    0.0026380058285488312, 0.0026996621780970113, 0.0027285261086932937, 
    0.0027231633734945472, 0.0026837120083021229, 0.0026117807430537958, 
    0.0025102541984549326, 0.002383030552197074, 0.0022347178378035104, 
    0.0020703097530137132, 0.0018948810093258404, 0.0017133096628640955, 
    0.0015300481801977818, 0.0013489469175775855, 0.0011731564195735598, 
    0.0010050807387257459, 0.00084639806932669483, 0.00069810880471826914, 
    0.00056060329747668859, 0.00043372942288654587, 0.00031685640263996745, 
    0.00020893680265737563, 0.00010857958981680902, 1.4126125071192008e-05, 
    -7.6264290388407737e-05, -0.00016452791902078973, -0.0002526200823189391, 
    -0.00034243991982927795, -0.00043576760237272553, 
    -0.00053417741334155211, -0.00063892278906419711, 
    -0.00075077949906349434, -0.00086986103262717742, 
    -0.00099543082642359151, -0.0011257646159212873, -0.0012580970860241083, 
    -0.0013887026096740709, -0.0015130978451085803, -0.0016263483340694955, 
    -0.0017234289533903696, -0.0017996011645307864, -0.0018508076110746602, 
    -0.0018740337346410667, -0.0018676421095363356, -0.0018316328630084775, 
    -0.0017677824755143062, -0.001679654274289884, -0.0015724508001723591, 
    -0.0014527197545898638, -0.0013279315638064855, -0.0012059766261425064, 
    -0.001094623478495057, -0.001000997393944795, -0.00093112546816724801, 
    -0.00088959435985430982, -0.00087934062608176005, -0.0009015811629820656, 
    -0.0009558723518331366, -0.0010402796127386787, -0.001151622675264548, 
    -0.0012857637734375149, -0.0014379100337453821, -0.0016029026142400872, 
    -0.0017754791701756365, -0.001950497200185372, -0.0021231060398376176, 
    -0.00228889056593202, -0.0024439723423931507, -0.0025850757878900575, 
    -0.0027095789699025066, -0.0028155325772309713, -0.0029016564843131832, 
    -0.0029673236400860805, -0.0030125117715357505, -0.003037763153129053, 
    -0.0030441334488930938, -0.0030331553491698823, -0.0030068025473258971, 
    -0.0029674260734322017, -0.0029176802504123876, -0.0028603845880267151, 
    -0.0027983688564616541, -0.0027342978420830059, -0.0026705108429376473, 
    -0.0026088875692127354, -0.0025507671372316655, -0.0024969086995398218, 
    -0.0024474981953131031, -0.0024021806032959829, -0.0023600969602831224, 
    -0.0023199139452835379, -0.0022798331597722334, -0.0022375967598853427, 
    -0.0021905034328307685, -0.0021354640012599961, -0.0020691315614205434, 
    -0.00198812072065774, -0.0018893040233575204, -0.0017701562195612894, 
    -0.0016290717979259408, -0.0014656207713092831, -0.0012806972889141935, 
    -0.0010765381232886383, -0.00085661869371082692, -0.00062542591014779934, 
    -0.00038813767224477427, -0.00015023735088120151, 8.2896990449949812e-05, 
    0.00030636142477535145, 0.0005160184669616817, 0.00070866228438609138, 
    0.0008820592092919073, 0.0010348441486556616, 0.00116633420841324, 
    0.0012762825540512202, 0.0013646374024578753, 0.0014313306569717077, 
    0.0014761353325639626, 0.0014985894520924622, 0.0014979886225936993, 
    0.0014734379907500185, 0.0014239587891210972, 0.0013486207733263516, 
    0.001246703822774775, 0.0011178675264675044, 0.00096232013082178148, 
    0.00078096076825746083, 0.00057549121255118382, 0.0003484694597840882, 
    0.00010329733051334258, -0.00015586762767798412, -0.00042425947471461741, 
    -0.00069672459489646989, -0.00096796603875686177, -0.0012328184812477033, 
    -0.0014865165648708309, -0.0017249309394947476, -0.0019447541428675504, 
    -0.0021436271232529521, -0.0023201785428856999, -0.002473996533408955, 
    -0.0026055329941121891, -0.0027159665067296832, -0.002807037218035712, 
    -0.0028808777913801238, -0.0029398398269813979, -0.0029863377621031544, 
    -0.0030227212556096263, -0.0030511646741882312, -0.0030735755230689109, 
    -0.0030915323236317144, -0.0031062274296824247, -0.0031184310421295538, 
    -0.0031284546277994207, -0.0031361529677443128, -0.0031409392922552557, 
    -0.003141839392208785, -0.0031375793725118835, -0.0031267104869127024, 
    -0.0031077492954834684, -0.0030793261834725209, -0.0030403328712479095, 
    -0.0029900457630846439, -0.0029282252911671581, -0.0028551686595687394, 
    -0.002771732211827064, -0.0026793002420590815, -0.0025797141220231731, 
    -0.0024751665369323957, -0.0023680599073416277, -0.0022608420809356296, 
    -0.0021558276298630731, -0.0020549988986101183, -0.0019598116023934356, 
    -0.0018710006495679856, -0.0017884060882760618, -0.0017108485385347741, 
    -0.0016360766199555027, -0.0015607928725946722, -0.0014807882328301577, 
    -0.0013911779306986793, -0.0012867066764395392, -0.0011621201563670274, 
    -0.0010125475370481975, -0.00083389427243921253, -0.00062317048382916059, 
    -0.00037878416368874215, -0.00010073214291162112, 0.00020927199164045367, 
    0.00054777010465005235, 0.00090960593232362527, 0.0012880591574923246, 
    0.0016750612546485699, 0.002061496321414215, 0.0024375753988401163, 
    0.0027932703688971542, 0.0031187869337411592, 0.0034050347198438056, 
    0.0036440643309875007, 0.0038294506876854319, 0.0039565819955341176, 
    0.0040228670526001979, 0.0040278262572384371, 0.0039731008262947178, 
    0.0038623579653301963, 0.0037011214425101361, 0.0034965256547090859, 
    0.0032570212787186117, 0.0029920261830316043, 0.0027115103468098554, 
    0.0024255614931656395, 0.0021439124190873187, 0.0018754758706951661, 
    0.0016279253792262267, 0.0014073462457209552, 0.0012179962069893192, 
    0.001062196423222234, 0.00094034107577447808, 0.00085102644505269344, 
    0.00079128105159575958, 0.00075685042931871425, 0.00074254179468292059, 
    0.00074255612295922929, 0.00075082298974175378, 0.00076129595124782405, 
    0.00076820967695963402, 0.00076629003562592082, 0.0007509257822075335, 
    0.00071829864657930878, 0.00066547995084163033, 0.00059049256069051883, 
    0.00049233342092932348, 0.00037095011522708839, 0.00022718362035574228, 
    6.2662883279408698e-05, -0.00012033614515261843, -0.00031905596189617838, 
    -0.00053043170005941456, -0.00075125819638601811, 
    -0.00097833514198410448, -0.0012085802167032447, -0.0014390920965554363, 
    -0.0016671780720808687, -0.0018903365554533017, -0.0021062011040279792, 
    -0.00231246758910787, -0.0025068039073848801, -0.0026867787362362754, 
    -0.0028498212461891392, -0.0029932576129586253, -0.0031144055015883063, 
    -0.003210759983941585, -0.0032802462894249251, -0.003321491327496704, 
    -0.0033340887205795108, -0.0033188029793824645, -0.0032776703366367375, 
    -0.0032139668476420737, -0.0031320635875775049, -0.0030371551128888681, 
    -0.0029349047810657137, -0.0028310472343249246, -0.0027309715082713226, 
    -0.0026393337592277811, -0.0025597464976377469, -0.0024945671715102019, 
    -0.002444814374652059, -0.0024102306989116458, -0.0023894629620223981, 
    -0.0023803421383409803, -0.0023802163657476293, -0.0023862966785133432, 
    -0.0023959697097371904, -0.0024070314480426707, -0.0024178453508367378, 
    -0.0024273844394510254, -0.002435170024167134, -0.0024411319032950065, 
    -0.0024453972951964309, -0.0024480596319199797, -0.0024489456992983576, 
    -0.0024474265744223924, -0.0024422738255092617, -0.0024315958244076528, 
    -0.0024128333917255995, -0.0023828526765911832, -0.0023380972097892003, 
    -0.0022748040307164377, -0.0021892547048771153, -0.0020780488175748783, 
    -0.0019383610868497628, -0.0017682054389537522, -0.0015666622425510655, 
    -0.0013340820644580677, -0.001072245803335927, -0.00078444406795361477, 
    -0.00047545587849137595, -0.00015140419711509806, 0.00018055186744306726, 
    0.00051264175982630787, 0.00083701551918992779, 0.0011463150812002548, 
    0.0014342134688049382, 0.0016958517620367624, 0.0019281287044259703, 
    0.0021297978297380453, 0.0023013765036718208, 0.0024448871434761812, 
    0.0025634777235177928, 0.0026609724035844785, 0.0027414393532728906, 
    0.0028088032974821972, 0.0028665771385930437, 0.0029177044184973719, 
    0.0029645219045801425, 0.0030088232948522319, 0.0030520012368366583, 
    0.0030952057552192914, 0.0031395233112057825, 0.0031861016617442824, 
    0.0032362362686540942, 0.0032913807021462981, 0.0033530785327608101, 
    0.0034228459450410232, 0.0035020134002313385, 0.0035915609626205811, 
    0.0036919863067057771, 0.0038032293622469954, 0.0039246609414969429, 
    0.0040550993368360221, 0.0041928715261874494, 0.0043358681677116402, 
    0.0044816094193872308, 0.0046273327293748171, 0.0047700948364008062, 
    0.0049068930425015178, 0.0050348169064467953, 0.0051511625475452062, 
    0.0052535101000556403, 0.0053397488110558848, 0.0054080621495334012, 
    0.0054568865330593451, 0.0054848778147976425, 0.0054908936638946035, 
    0.0054739995122824797, 0.0054335077352283987, 0.00536900415382728, 
    0.0052803925499082718, 0.0051679211958087449, 0.0050321987008470981, 
    0.0048741946111559922, 0.004695221226065774, 0.004496892463763405, 
    0.0042810695038919336, 0.0040498143470275904, 0.00380537615657244, 
    0.0035502566501973442, 0.0032873259182956238, 0.0030199889246771308, 
    0.0027523283658166127, 0.0024891709547643945, 0.0022360362792298175, 
    0.0019989402103410187, 0.0017840577940691719, 0.0015972862981635553, 
    0.0014437540674304384, 0.0013273379687759972, 0.0012502422262221651, 
    0.0012127088949479073, 0.0012129090005878727, 0.0012470403998542201, 
    0.0013096380369127323, 0.0013940873574102466, 0.0014932618279797519, 
    0.001600245198531771, 0.001709009252475853, 0.001814989846338365, 
    0.0019154538295921189, 0.0020096284383815393, 0.0020985666303929675, 
    0.00218478933477832, 0.0022717547020597497, 0.0023632446416271872, 
    0.0024627530568338139, 0.0025729463138524601, 0.002695263199221695, 
    0.0028296811748980215, 0.0029746676778202742, 0.003127314122970687, 
    0.0032836180007849406, 0.0034388799006606712, 0.0035881406305135438, 
    0.0037266001484331022, 0.0038499731845625181, 0.003954743346719242, 
    0.0040383107100172037, 0.0040990565960716775, 0.0041363395461613897, 
    0.0041504332468959857, 0.0041424458677966512, 0.0041141710262439192, 
    0.0040679156398620167, 0.0040062792671304919, 0.0039319053066388804, 
    0.0038472611065611746, 0.0037544292326272934, 0.0036549567138220856, 
    0.0035497819125459552, 0.0034392171353351732, 0.0033230098316187461, 
    0.0032004811226940735, 0.00307069848282184, 0.0029326907842466268, 
    0.0027856616038388613, 0.0026292034919596211, 0.0024634697491541968, 
    0.0022893184469818507, 0.0021083871681502652, 0.0019230969410482187, 
    0.001736537798665873, 0.0015522483567490602, 0.0013738699767576934, 
    0.0012047175781131941, 0.0010473249098794178, 0.00090301942475089474, 
    0.00077160169431351447, 0.00065118537302636748, 0.00053824199212596294, 
    0.00042782517681340968, 0.00031397336487922254, 0.00019022452796609168, 
    5.0189702643414836e-05, -0.0001118770549123385, -0.00030056046465524485, 
    -0.00051887853264886746, -0.00076800864198599977, -0.0010471723536130348, 
    -0.0013536624963979712, -0.0016829812234105937, -0.0020290737471044817, 
    -0.0023845969714869999, -0.00274121352117792, -0.003089878114137802, 
    -0.0034211352067235723, -0.0037253970920165529, -0.0039932217384618897, 
    -0.0042155877053789191, -0.0043841812037783909, -0.0044916734251212159, 
    -0.004532004744504302, -0.0045006605604676966, -0.0043949225332657448, 
    -0.0042140999487062713, -0.0039597136464200903, -0.0036356183696081026, 
    -0.0032480472675458188, -0.0028055641049126198, -0.0023188675846411606, 
    -0.0018004675660205024, -0.0012642054657366329, -0.00072464960358635652, 
    -0.00019639309617601838, 0.00030668803051531771, 0.000772131693904695, 
    0.0011894890162449361, 0.0015507387020317607, 0.0018505064999457021, 
    0.0020860686348338022, 0.0022571619995060957, 0.0023656558202318394, 
    0.0024151488792600903, 0.0024105290629270887, 0.0023575657679336796, 
    0.0022625598700275387, 0.0021320698207690988, 0.0019727263232922842, 
    0.0017911348169582602, 0.0015938375116569478, 0.0013873085940494904, 
    0.0011779582716267868, 0.00097210879687302293, 0.00077594546636790111, 
    0.00059543142325878143, 0.00043620662342115185, 0.00030348526115725748, 
    0.00020194617607110235, 0.00013566402871520713, 0.00010806081617805273, 
    0.00012187492194373914, 0.00017914388665360458, 0.00028118445049711961, 
    0.0004285177158542447, 0.00062077848798264507, 0.00085656755977935766, 
    0.0011333021065964197, 0.0014470538366520977, 0.0017924387969879422, 
    0.0021625652342703644, 0.0025490819788530957, 0.0029423391232019985, 
    0.0033316652385180019, 0.0037057670988990968, 0.0040532165782911677, 
    0.0043630220032167882, 0.0046252293374314914, 0.0048315149992269662, 
    0.0049757111010970845, 0.0050542350305878957, 0.0050663609734878066, 
    0.0050143122460516347, 0.0049031575229910489, 0.0047405258011388313, 
    0.0045361378823773795, 0.0043012017350277749, 0.0040476987009135743, 
    0.0037876246125854167, 0.0035322263815232924, 0.0032913170831555469, 
    0.0030727144049469278, 0.0028818489179610611, 0.0027215763762511928, 
    0.002592188320515461, 0.0024916078938993307, 0.0024157448292223861, 
    0.0023589593405988272, 0.002314587005461736, 0.0022754734761658148, 
    0.0022344895173448472, 0.0021849531545156428, 0.0021209814265511859, 
    0.0020377263611024241, 0.0019315075657223, 0.001799871744040542, 
    0.0016415756443770848, 0.0014565265140544877, 0.0012456916436636887, 
    0.0010109906193100373, 0.00075516419116452584, 0.00048163959868667875, 
    0.00019437837349671548, -0.00010227296424174618, -0.00040373092937697386, 
    -0.00070534433542650472, -0.0010025265288865239, -0.0012909306343980359, 
    -0.0015665883951797627, -0.0018260859260868562, -0.0020667190428186356, 
    -0.0022866525160948172, -0.0024850451806236588, -0.0026621389121400476, 
    -0.002819278325210737, -0.002958854388461133, -0.0030841594521572092, 
    -0.0031991197397136747, -0.003307930392326353, -0.0034145772387920805, 
    -0.00352232130688814, -0.0036331897027647056, -0.0037475726912912198, 
    -0.0038639829978313052, -0.0039790350613295149, -0.0040876486532183823, 
    -0.0041834718712306391, -0.004259454640641723, -0.0043085225658088776, 
    -0.0043242620763881603, -0.0043015776629659712, -0.0042372019772931556, 
    -0.0041300762614756162, -0.0039815174560877053, -0.0037951940833565027, 
    -0.0035768914913728959, -0.003334098995173044, -0.0030754554844947108, 
    -0.0028101028156061201, -0.0025470087961271186, -0.00229430659403274, 
    -0.0020587322845673547, -0.0018451763620907368, -0.0016564219031731569, 
    -0.0014930701522617893, -0.001353662074711317, -0.0012349730567652966, 
    -0.001132464307234022, -0.0010408189352313845, -0.00095452735956711376, 
    -0.00086846277754800999, -0.00077840014621483879, 
    -0.00068143681646397726, -0.00057627491140212856, 
    -0.00046339263861200488, -0.00034501785958807263, -0.0002249724031368866, 
    -0.00010834581749035877, -1.0492470946294744e-06, 9.0709082788057661e-05, 
    0.00016095434863778007, 0.00020443985735481176, 0.0002170422977259241, 
    0.00019604473695498907, 0.00014025616318166648, 5.0010441491699241e-05, 
    -7.293902073218691e-05, -0.00022559585309955401, -0.00040392907508120723, 
    -0.00060311392673179597, -0.00081776634256483733, -0.0010421901455487112, 
    -0.0012705807517207179, -0.0014972106404661117, -0.0017165756285073299, 
    -0.0019235039455888182, -0.0021132544611271284, -0.0022816175175801295, 
    -0.0024250158793744621, -0.0025406454339160418, -0.0026266143580038134, 
    -0.0026820801804247076, -0.002707380720232435, -0.0027041026834128479, 
    -0.0026750818635266306, -0.0026242942284407677, -0.0025566402153661106, 
    -0.0024776254006583865, -0.0023929500331885895, -0.0023080862817818084, 
    -0.00222786030163838, -0.00215612880305326, -0.0020955778908932276, 
    -0.0020476595149879918, -0.0020126563835143408, -0.001989843297143325, 
    -0.0019776918412700447, -0.0019740680260399942, -0.0019764161944117314, 
    -0.0019819091884661698, -0.0019875772718730552, -0.001990460378364207, 
    -0.0019877797058379942, -0.0019771473069577781, -0.0019567936338551108, 
    -0.0019258034367364632, -0.0018843071174290387, -0.0018336232648987084, 
    -0.0017762696257955192, -0.0017158869314709869, -0.0016570081165903209, 
    -0.0016047039137220128, -0.0015640955763792444, -0.0015397797294870233, 
    -0.0015352491155598146, -0.0015523817779545695, -0.001591125726979174, 
    -0.0016493993718646762, -0.0017232294303040556, -0.0018070663986469208, 
    -0.0018942481476290863, -0.001977524248952073, -0.0020495882957797047, 
    -0.0021035196275638228, -0.0021331311946979118, -0.0021331640789019795, 
    -0.0020993668832510037, -0.0020284928670112651, -0.0019182715889773201, 
    -0.0017673905457624224, -0.0015755103876199832, -0.0013432823833864321, 
    -0.0010724193581180886, -0.00076575452712012695, -0.00042730368256064789, 
    -6.2291973824982178e-05, 0.00032288325370966113, 0.00072076865241933144, 
    0.0011230709928594972, 0.0015209480169965305, 0.0019053868757171481, 
    0.0022676250538096556, 0.0025995875251190515, 0.0028942911824490587, 
    0.0031461779676059043, 0.0033513442644752269, 0.0035076434758152648, 
    0.0036146571037584561, 0.0036735431937416278, 0.0036868005812056644, 
    0.0036579956318398342, 0.0035914697373484101, 0.0034920830655232318, 
    0.0033649946104403658, 0.0032155233416484652, 0.0030490440165364214, 
    0.0028709488420102574, 0.0026866318256478696, 0.0025014666947966451, 
    0.0023207662916639397, 0.0021496721452534564, 0.0019929907897931571, 
    0.001854966552505494, 0.0017390365680852013, 0.0016476195637029013, 
    0.0015819922618567207, 0.0015422734976898414, 0.0015275079740706093, 
    0.0015358107573924312, 0.0015645205643736761, 0.0016103359174941855, 
    0.0016694471315572984, 0.0017376611659393369, 0.0018105712811065631, 
    0.0018837441558025522, 0.0019529511336313274, 0.0020143824508150497, 
    0.0020648322328847874, 0.0021018216482975387, 0.0021236570815014958, 
    0.0021294193218539289, 0.0021188997246989276, 0.002092482703721847, 
    0.0020509965930606278, 0.0019955299598846733, 0.0019272554977738526, 
    0.0018472670332072404, 0.0017564444882752148, 0.0016554108161442676, 
    0.001544534899658029, 0.0014240283792104156, 0.0012940553926126591, 
    0.0011548977200694914, 0.0010071008383513373, 0.00085159918302463774, 
    0.00068981686950772298, 0.00052369021161829759, 0.00035565779877521877, 
    0.00018858902806450782, 2.567735511474387e-05, -0.00012968623079210315, 
    -0.0002740181510258019, -0.0004038682368479946, -0.00051591180566453181, 
    -0.00060703022913001178, -0.00067440050735346362, -0.0007155914379001633, 
    -0.00072866265105451698, -0.00071230136474195391, 
    -0.00066596654109853223, -0.00059007547221976212, 
    -0.00048617640719054902, -0.00035711637655021157, 
    -0.00020713216233661025, -4.1838169116749137e-05, 0.00013193578456996064, 
    0.00030645985835722452, 0.00047356501482720317, 0.00062522531809445538, 
    0.00075417567466006625, 0.0008545332009839274, 0.00092231542946692258, 
    0.00095582800327825238, 0.00095585210856983041, 0.00092561124049957263, 
    0.00087051970464670355, 0.00079771543976329138, 0.00071545345899682656, 
    0.00063236883526112905, 0.00055672022314774249, 0.0004956502718799215, 
    0.00045451849173732968, 0.00043637909242900307, 0.00044162422237853014, 
    0.00046782034514723005, 0.00050978952671608846, 0.00055990985681972848, 
    0.00060861751814768946, 0.00064510145827711832, 0.00065809994944974245, 
    0.00063675603841812473, 0.00057145487992502552, 0.00045459192738576173, 
    0.00028123367001396497, 4.9603142043018473e-05, -0.00023862985282105357, 
    -0.00057826697359483282, -0.00096074941561261355, -0.0013745876715599852, 
    -0.001806009028729373, -0.002239829494759529, -0.0026604509314896597, 
    -0.0030528682745752469, -0.0034035984199512377, -0.0037014103871311757, 
    -0.0039378707150710159, -0.0041076293817832923, -0.0042085109308200551, 
    -0.0042414169357078927, -0.0042100473863663484, -0.0041204822408198016, 
    -0.0039806594979571825, -0.0037997754335900142, -0.0035876767755771174, 
    -0.0033542939088752059, -0.0031091580813748035, -0.0028610418791390926, 
    -0.002617670071893524, -0.0023855488041042341, -0.0021698210334271054, 
    -0.0019741582899145856, -0.0018007085775895587, -0.0016500709826618742, 
    -0.0015213358111698574, -0.0014121565313490428, -0.0013188867935201693, 
    -0.0012367792268450047, -0.0011603160845052964, -0.0010836311052435164, 
    -0.0010010036247503433, -0.0009073192115339598, -0.00079847233635519602, 
    -0.00067161844451527628, -0.00052534236456605328, 
    -0.00035971703245004375, -0.00017629665440802069, 2.1933745656679392e-05, 
    0.00023069113093056217, 0.00044457430925428694, 0.00065731631197874592, 
    0.00086212339338468996, 0.0010520153519667284, 0.0012201871884214514, 
    0.0013603591145219284, 0.0014670940813390045, 0.0015361000478208767, 
    0.0015644802164836043, 0.0015509388331622035, 0.0014959118351764219, 
    0.0014016355100626365, 0.001272118017971014, 0.0011130053185176639, 
    0.00093134122969810377, 0.00073522134649083612, 0.00053337173837359375, 
    0.00033467646248746505, 0.00014770262438842653, -1.9750892499841327e-05, 
    -0.00016106623666452445, -0.00027113827277852783, 
    -0.00034660404835087661, -0.00038596113249795216, 
    -0.00038950276345686219, -0.00035912626326621176, 
    -0.00029798504162611967, -0.00021005510205137747, 
    -9.9668077880689943e-05, 2.8919690917857244e-05, 0.00017186452099672911, 
    0.00032595039082429158, 0.00048868676575802221, 0.00065826883746338937, 
    0.00083347341828437984, 0.0010134803563558818, 0.0011976440969980108, 
    0.0013852890948327101, 0.0015754996044475078, 0.0017669537980705367, 
    0.0019578145220409062, 0.002145705970491912, 0.0023277800382105105, 
    0.0025008804828109202, 0.0026617697924035395, 0.0028074329150693422, 
    0.0029353714124522867, 0.003043899934042406, 0.0031323607319762672, 
    0.0032012432790150228, 0.0032522124795617206, 0.0032879818094011847, 
    0.0033121117014525752, 0.0033287244134710095, 0.0033421481913609259, 
    0.003356543454279535, 0.0033754845335191934, 0.0034015398074885, 
    0.0034358236362774246, 0.0034776115799109333, 0.0035240915408094042, 
    0.0035703955194619566, 0.0036100018886939659, 0.0036355198538538178, 
    0.0036397154970709274, 0.0036165525089126844, 0.0035619898642399771, 
    0.003474391830748904, 0.003354512951349298, 0.0032052128350680874, 
    0.0030310663462901201, 0.0028379022725764265, 0.0026323950712246027, 
    0.0024217195722459669, 0.0022132067092264151, 0.0020140926792389501, 
    0.0018312591172180855, 0.0016710235675312297, 0.0015389409887307493, 
    0.001439597828890899, 0.0013764384483920379, 0.0013515839114704561, 
    0.0013656911560693096, 0.0014177978953478448, 0.0015052568737643243, 
    0.0016237105127476874, 0.0017671730809102925, 0.0019282062276336862, 
    0.0020981884480019168, 0.0022676924076414423, 0.0024269210820513517, 
    0.0025662050437007325, 0.0026764909470999325, 0.0027498412019725592, 
    0.0027798431125632054, 0.0027619151734506603, 0.0026934441393310707, 
    0.0025737629466004801, 0.0024039573640442305, 0.0021865412316427364, 
    0.0019250678529147184, 0.0016237288535178637, 0.0012869793673418489, 
    0.00091926633041676368, 0.0005248341072473493, 0.00010760049336557844, 
    -0.00032884437235612186, -0.00078117752445654469, -0.0012462296956961697, 
    -0.0017208168417621916, -0.0022015856206280267, -0.0026848554505859231, 
    -0.0031665577752761553, -0.0036422420834181456, -0.0041071683344367721, 
    -0.0045564836540831393, -0.0049854781818774382, -0.0053898550055931343, 
    -0.0057659591245574149, -0.0061109345174799505, -0.0064227285929680548, 
    -0.0066999613115138936, -0.0069416706738732094, -0.0071470155544807864, 
    -0.0073149794702064182, -0.007444152077887475, -0.0075326878002387326, 
    -0.0075784179526217762, -0.007579083589971421, -0.0075326020714175101, 
    -0.0074372658562891873, -0.0072919047206272455, -0.007096036570271835, 
    -0.0068500255418422473, -0.0065552077188994881, -0.0062139428762331217, 
    -0.0058295136177582392, -0.0054058826628012226, -0.0049473603167284616, 
    -0.00445822491462419, -0.0039425180930345669, -0.0034039617786263492, 
    -0.0028461228013195081, -0.0022727661539737754, -0.0016882942615598874, 
    -0.0010981139151651973, -0.00050882555059075167, 7.1844506993997944e-05, 
    0.00063541869212898412, 0.00117326912547208, 0.0016772975037650558, 
    0.0021405971665837526, 0.0025579585493317471, 0.0029261379806672567, 
    0.0032439126568275865, 0.0035119149659776556, 0.0037323078501617559, 
    0.0039083613043814861, 0.0040439658182320152, 0.0041431308464480801, 
    0.0042094981906144555, 0.0042459235098008521, 0.0042542175021666488, 
    0.0042349680545264688, 0.0041875384837865943, 0.0041102017774636481, 
    0.0040004256571321986, 0.0038552278376833586, 0.0036716914760629533, 
    0.0034474229446115586, 0.0031810323773181783, 0.0028725023591188795, 
    0.0025234836807390506, 0.0021374342815855345, 0.0017196839499004427, 
    0.0012773524916953796, 0.00081916024933176019, 0.00035511963924972459, 
    -0.00010391036151906574, -0.00054675290277199655, 
    -0.00096254860118922224, -0.0013414149020966103, -0.0016750929098978363, 
    -0.0019575035634593189, -0.002185143678167713, -0.0023572688186857655, 
    -0.0024758855453644243, -0.0025454778585723443, -0.0025725681714044071, 
    -0.002565149789791978, -0.0025320663056246605, -0.0024823765373737051, 
    -0.0024248562004070364, -0.0023675400105681163, -0.0023174571718741969, 
    -0.0022804465868136842, -0.0022611213592118331, -0.0022628861886324369, 
    -0.0022880052934719374, -0.0023377169275838523, -0.0024123680368526297, 
    -0.0025115467041060611, -0.0026342782527437832, -0.0027792296621565525, 
    -0.0029449343142244834, -0.0031300171862115415, -0.0033333391637578977, 
    -0.0035540665817586155, -0.0037916212963720912, -0.0040454793781788765, 
    -0.0043149308441301328, -0.0045988131245476085, -0.0048952496351714267, 
    -0.0052015012806014074, -0.0055138863675069589, -0.0058278684550134565, 
    -0.00613822977782825, -0.0064394092918594603, -0.0067258510755509341, 
    -0.006992357198509656, -0.0072343915309015941, -0.0074483229376426955, 
    -0.0076316126308875803, -0.0077829459235471098, -0.0079022942882437299, 
    -0.0079908759046139217, -0.0080510389232453065, -0.0080860541718628179, 
    -0.0080997829057597951, -0.0080963359831845959, -0.0080796447763074233, 
    -0.0080530569134011198, -0.0080189450756040833, -0.0079783513181544939, 
    -0.0079307665712487554, -0.0078739905553185593, -0.0078041772633532739, 
    -0.0077160283125576939, -0.0076032394317629712, -0.0074590030022512223, 
    -0.0072766902467036876, -0.0070505541135726726, -0.006776399085330502, 
    -0.006452167035683006, -0.0060783352698906236, -0.005658131111781782, 
    -0.0051974908847411301, -0.0047047978251232685, -0.0041904208144346571, 
    -0.0036660397448383185, -0.0031438683080194682, -0.0026358130754346979, 
    -0.0021526552791140932, -0.0017033885870575965, -0.001294814166949057, 
    -0.00093133765158139677, -0.00061512290137833651, 
    -0.00034642648832736655, -0.00012405291798502159, 5.4145476202231908e-05, 
    0.00019088102161445936, 0.00028914020174577814, 0.00035203587283096478, 
    0.00038279319133907949, 0.00038483853092402217, 0.00036195823988888817, 
    0.00031843943564557398, 0.00025926488994394025, 0.00019024753252836122, 
    0.00011810097527873961, 5.0407991545061058e-05, -4.5553933266398556e-06, 
    -3.8138063129541924e-05, -4.1789988791840414e-05, 
    -7.6669262762908383e-06, 7.0744084804954155e-05, 0.00019797943826361099, 
    0.00037606880892851902, 0.00060417678107516927, 0.00087843704865520891, 
    0.0011920709820054563, 0.0015356816554132429, 0.0018977729769594819, 
    0.0022653971419701862, 0.0026248656559918139, 0.0029625452363411207, 
    0.0032655606380255137, 0.0035225185293062079, 0.0037240672440049089, 
    0.003863345188336947, 0.0039362524219667934, 0.0039415383971747693, 
    0.0038807223478081344, 0.003757832914637293, 0.0035790664612087709, 
    0.0033523347441638579, 0.0030867880382330721, 0.0027923108601128769, 
    0.0024790284923865116, 0.0021568410302202964, 0.0018350033651481727, 
    0.0015218153897176472, 0.0012243557761946406, 0.00094842035834483487, 
    0.00069855899601293386, 0.00047823404059423952, 0.00029013784036878649, 
    0.00013646084665478494, 1.9239966496665303e-05, -5.9414389213063835e-05, 
    -9.7172458347776384e-05, -9.1547018263765401e-05, 
    -4.0039592048715277e-05, 5.9488962217234903e-05, 0.00020838545867265675, 
    0.00040668261736118009, 0.00065260609620145416, 0.00094225175264807241, 
    0.0012693920438999653, 0.0016254475388970745, 0.0019996528704748751, 
    0.0023793989715356631, 0.0027506352795690155, 0.0030984376438298309, 
    0.0034076312228779565, 0.0036635238164966681, 0.0038526830067999447, 
    0.0039637590521935219, 0.0039881679608437014, 0.0039206544741062967, 
    0.0037595722200993069, 0.0035070061429199949, 0.0031686235586366627, 
    0.0027533027493789781, 0.0022725329434940358, 0.0017397107328165039, 
    0.0011692042869131181, 0.00057542123764464149, -2.8113133374927703e-05, 
    -0.0006294894709942577, -0.0012189413184164187, -0.0017890401652707181, 
    -0.0023346500419256428, -0.0028526635958626614, -0.0033415584089218232, 
    -0.0038008753800950054, -0.0042306210265499154, -0.0046308025551846385, 
    -0.0050010983481255404, -0.0053409098205644909, -0.0056498520190206812, 
    -0.0059285535928202066, -0.0061792586721913746, -0.0064058691239955411, 
    -0.0066133091018748856, -0.0068065495676715654, -0.0069896944837301656, 
    -0.0071655201651266353, -0.0073353694103676682, -0.0074993309721761436, 
    -0.0076566114928237929, -0.0078058531927269843, -0.0079454846665738214, 
    -0.0080739197951701421, -0.008189739733550876, -0.0082918521181490016, 
    -0.0083795721580768937, -0.0084527300591798714, -0.0085117443434734649, 
    -0.0085577582354835462, -0.0085927865021478214, -0.0086199559343848476, 
    -0.0086436173520038299, -0.0086693065832415886, -0.0087034221964319182, 
    -0.0087525390195747777, -0.0088225142194716961, -0.0089174357180405103, 
    -0.0090387061682681343, -0.0091842726509163072, -0.0093484050763797486, 
    -0.0095219023134838921, -0.00969290080305041, -0.0098480676230793106, 
    -0.0099741188571027366, -0.010059364990759547, -0.010095010565711384, 
    -0.010076111598605886, -0.010001892680854616, -0.0098756312508040209, 
    -0.0097040803220255697, -0.0094966697405393635, -0.0092644829068157953, 
    -0.009019327054280598, -0.0087726472192047582, -0.0085345982465712938, 
    -0.0083130969300862639, -0.0081131455389004195, -0.0079364850505156074, 
    -0.0077815427211787615, -0.0076438419142314321, -0.007516531720749728, 
    -0.0073912078472666105, -0.0072587367840441005, -0.0071103419717183239, 
    -0.0069385118198808538, -0.0067380136227301905, -0.0065067512123524801, 
    -0.0062462938108541512, -0.0059621624173046908, -0.0056636756548102312, 
    -0.0053634974805136602, -0.0050768665132173247, -0.0048207056178537731, 
    -0.0046126633133907503, -0.0044701742706803648, -0.0044096327504545754, 
    -0.0044457048204935672, -0.0045906954453767898, -0.0048539250035409881, 
    -0.0052412668370442356, -0.0057546369063446222, -0.0063917116929607144, 
    -0.0071458993937140881, -0.0080064667902567249, -0.0089590345105808565, 
    -0.0099862044314859774, -0.011068315951626825, -0.012184105502822231, 
    -0.013311450088705486, -0.014427916563758638, -0.015511503365121112, 
    -0.016541534775666434, -0.017499551090529444, -0.018370358324628168, 
    -0.019142796853425958, -0.019810332392769511, -0.020371405870401111, 
    -0.020829332060652295, -0.021192051281892339, -0.021471389424816367, 
    -0.021682142915966453, -0.021840758430711336, -0.021963706639091342, 
    -0.022065818508958973, -0.022158687009094305, -0.022249299074808545, 
    -0.022339335570642386, -0.022425277869481574, -0.02249932972957926, 
    -0.022551184385884541, -0.02257020366337965, -0.022547517428718359, 
    -0.022477374112685928, -0.022357685476761601, -0.022189783335488759, 
    -0.021977683344814654, -0.021727271521098004, -0.021445657751277894, 
    -0.021140691159324328, -0.020820989765041861, -0.020496027027365853, 
    -0.020176574175790028, -0.019874942181051364, -0.019604810594936711, 
    -0.019380823313593733, -0.01921754317698068, -0.019127929436542356, 
    -0.019121742046552936, -0.019203613758667023, -0.019371595387868853, 
    -0.019615951592122052, -0.019918562100933696, -0.020253227370377019, 
    -0.020586341853426345, -0.020878474873367237, -0.021086163599248541, 
    -0.021164373867570592, -0.021068923889508623, -0.020759471527896797, 
    -0.020202238187019505, -0.019372937630884601, -0.018259384107297466, 
    -0.016863287170631555, -0.015200965504738562, -0.013302436409290894, 
    -0.011209356122257083, -0.0089716289120017317, -0.006643834440364883, 
    -0.0042815524027103539, -0.0019381022683262396, 0.00033859703140303289, 
    0.0025082575785243437, 0.004541148783776751, 0.0064192556390835964, 
    0.0081366972023290095, 0.0096978929552718092, 0.011113965418146729, 
    0.012397524784097983, 0.013557032362535682, 0.014592165058949925, 
    0.015490744593065828, 0.016228531451865362, 0.016771481236658066, 
    0.017080292631844039, 0.01711599749706522, 0.016845989722704197, 
    0.016248562094692571, 0.015315667928524349, 0.014053345473193883, 
    0.012480800137949881, 0.010627794831208797, 0.0085317911814862292, 
    0.0062349576320649292, 0.0037822716213524532, 0.0012194278559345077, 
    -0.0014084492383777817,
  // Fqt-total(8, 0-1999)
    0.99999999999999956, 0.99221724269879774, 0.96927513582182034, 
    0.9323516072116903, 0.88328471607289216, 0.82440567373461593, 
    0.75833905558482073, 0.68779590371324673, 0.61538343115702832, 
    0.54344966293847818, 0.4739739548679846, 0.40850655416137394, 
    0.34815376668422071, 0.29360056325617118, 0.24515991770950615, 
    0.20283786399234219, 0.16640432778106581, 0.13546200212147022, 
    0.10950795085763762, 0.087985109248613511, 0.07032264693339231, 
    0.055965652914081801, 0.044395376638239996, 0.035141624267646401, 
    0.027789018249531051, 0.02197863653101376, 0.017406395850705483, 
    0.013819286000848691, 0.011010324148548804, 0.00881287983700107, 
    0.0070948021797815055, 0.005752656874113163, 0.0047063149584996994, 
    0.0038940159714355269, 0.003268058364854907, 0.0027911862581186677, 
    0.0024337305805698082, 0.0021714681176079496, 0.0019841300026186147, 
    0.0018544452243814222, 0.0017675562483943192, 0.0017106873668716663, 
    0.0016729165602220209, 0.0016450121535915407, 0.0016192557084743185, 
    0.0015892729700051446, 0.0015498640152159079, 0.0014968541737353466, 
    0.0014269629738012184, 0.0013376939190873939, 0.0012272508242815675, 
    0.0010944978420731736, 0.00093894652819949214, 0.00076078471469476423, 
    0.00056093316856979756, 0.00034109925695796693, 0.00010382815369124125, 
    -0.00014749193838713129, -0.00040868475383385984, -0.000674887541814162, 
    -0.00094072476429783844, -0.0012005346319465063, -0.0014486488462871353, 
    -0.0016797142406049142, -0.0018890559427258778, -0.0020730362289305077, 
    -0.0022293780606063547, -0.0023573644159090752, -0.0024578756181787152, 
    -0.0025332460387884046, -0.0025869752596632658, -0.0026233530661163721, 
    -0.0026470556680953466, -0.0026627246196368856, -0.0026745637732033044, 
    -0.002685937780264591, -0.0026990136305415574, -0.0027144651154604976, 
    -0.0027313006237561048, -0.0027468486005906901, -0.0027569372827139609, 
    -0.0027562621652617975, -0.0027388976369121494, -0.0026988947169031361, 
    -0.0026308831908849395, -0.0025305827804540013, -0.0023951575052015579, 
    -0.0022233677177525531, -0.0020155308008640797, -0.0017733065260644605, 
    -0.0014994149238735611, -0.0011973462248766604, -0.00087112947257461562, 
    -0.00052520158747685209, -0.00016435327769417503, 0.00020626094549842962, 
    0.00058109072738118299, 0.00095417077534711904, 0.0013191318562299137, 
    0.0016692727153270689, 0.0019977036352031318, 0.0022975474951891328, 
    0.0025622029168589949, 0.0027856257243716338, 0.0029626276169114189, 
    0.003089151215942778, 0.003162533114224, 0.0031817325335024766, 
    0.0031475363954857325, 0.0030627013912940672, 0.0029320332813926645, 
    0.0027623512797700033, 0.0025623080691403125, 0.0023420571640051517, 
    0.0021127479536969403, 0.0018858969091866387, 0.0016726812683233786, 
    0.0014832433016473421, 0.0013260910781945337, 0.001207664036270249, 
    0.001132097163970234, 0.0011011857863632564, 0.0011145366407285268, 
    0.0011698391640729497, 0.0012632056596612532, 0.0013895138310802435, 
    0.0015427230338116275, 0.0017161374527389051, 0.0019026435867669491, 
    0.0020949379630529341, 0.0022857741923921885, 0.0024682328906605313, 
    0.0026359931126735368, 0.002783574850838006, 0.0029065152367745433, 
    0.0030014535001799993, 0.0030661091247757718, 0.0030991817712248274, 
    0.0031001808007849185, 0.0030692365225097897, 0.0030069387968811975, 
    0.0029142239901701191, 0.0027923615505234443, 0.0026430305563515419, 
    0.002468484503035581, 0.0022717465809627187, 0.0020568131378132233, 
    0.0018287811053298744, 0.0015938632627840181, 0.0013592450240516093, 
    0.001132750275814479, 0.0009223499109134066, 0.00073553534137598797, 
    0.00057863887942569971, 0.00045619892251529641, 0.00037046276318418718, 
    0.00032111921105626602, 0.00030531988876070411, 0.00031800769409226482, 
    0.00035249777456845317, 0.00040122292029931762, 0.00045652724646718339, 
    0.00051136468867278107, 0.0005598358352595196, 0.00059752688540447687, 
    0.00062164297490222497, 0.00063100299974049999, 0.00062592490753148196, 
    0.00060805715142532146, 0.00058016857019334571, 0.00054590701084454888, 
    0.00050952338615120553, 0.000475551567194463, 0.00044846847935726172, 
    0.00043234974037060662, 0.00043054259185536551, 0.0004453855653388149, 
    0.00047798694766301432, 0.00052809759519509703, 0.00059408311640991385, 
    0.00067300079131923105, 0.00076079237590007446, 0.00085256711752475808, 
    0.00094296730077418514, 0.001026583077003046, 0.0010983852619747797, 
    0.0011541422773031073, 0.0011907991271589357, 0.0012067797033336503, 
    0.0012021970979434785, 0.0011789257708788041, 0.0011405335446394898, 
    0.0010920417694609916, 0.0010395271232356493, 0.00098959429222168467, 
    0.00094877080987664528, 0.00092291356840763837, 0.00091669631962901438, 
    0.00093325271210267899, 0.00097400578343885655, 0.0010387091234000431, 
    0.0011256743918564296, 0.0012321230473727788, 0.0013546091032199882, 
    0.0014894336653766805, 0.0016329849327308792, 0.0017819660755594787, 
    0.0019334925937558051, 0.0020850760694195464, 0.0022345405322267264, 
    0.0023799039396134596, 0.0025192852269133505, 0.0026508663890657579, 
    0.0027729208565016499, 0.0028838983771344055, 0.0029825462733807941, 
    0.0030680466102290258, 0.003140120178664513, 0.0031990892879713187, 
    0.0032458579489094523, 0.0032818212005503071, 0.0033086787254682911, 
    0.0033281963162318305, 0.0033419255493827736, 0.0033509469468946682, 
    0.0033556541034146948, 0.003355650188658404, 0.0033497488312246122, 
    0.0033360972793894349, 0.0033123932625601692, 0.0032761573105821655, 
    0.0032250242735277169, 0.0031570003619500703, 0.0030706741802129368, 
    0.0029653625733165713, 0.0028411863075161483, 0.0026990992891387754, 
    0.0025408751607693862, 0.002369063916107317, 0.0021869266487393453, 
    0.0019983442636976267, 0.0018076902915190643, 0.0016196496425565801, 
    0.0014389898925814173, 0.0012702714290662809, 0.00111752386186319, 
    0.00098392697360804118, 0.00087151499093705126, 0.00078095661980279608, 
    0.00071143812718489521, 0.0006606831609467773, 0.00062509934388638231, 
    0.000600067623027601, 0.00058032139180937017, 0.00056037737718372623, 
    0.00053494594773628766, 0.00049928180661743362, 0.00044940636094125438, 
    0.00038222302995383667, 0.00029552283704481101, 0.0001879376620999866, 
    5.8880484100119385e-05, -9.1494784387803992e-05, -0.00026227246553003816, 
    -0.00045172284500368123, -0.00065720675661113336, 
    -0.00087509434421992349, -0.0011007295680274913, -0.0013284775635309829, 
    -0.0015518973118730127, -0.0017640426412497661, -0.0019578687074103696, 
    -0.0021267285865033216, -0.002264891043221055, -0.002368030795305261, 
    -0.0024336338799389491, -0.0024612625331575325, -0.0024526592077521174, 
    -0.0024116415444780468, -0.0023438065860921235, -0.0022560474627483528, 
    -0.0021559414107606019, -0.0020510615514058935, -0.0019483158774920304, 
    -0.0018533807902310648, -0.001770313586540934, -0.0017013572532209652, 
    -0.0016469678979005769, -0.0016060113422707307, -0.0015760900509642372, 
    -0.0015539313213216548, -0.0015357763909376295, -0.0015177245896284665, 
    -0.0014959993194254653, -0.0014671339844783973, -0.0014280798798207216, 
    -0.0013762601340027703, -0.0013095873475086179, -0.0012264840481340951, 
    -0.00112590111057304, -0.0010073705858993764, -0.00087108653049643538, 
    -0.00071800686255033843, -0.00054996603182671773, 
    -0.00036976762055085838, -0.00018124365062306875, 1.0764584089754337e-05, 
    0.00020050199597441528, 0.00038151027436423516, 0.00054693600515405918, 
    0.00068993249684215041, 0.00080411017204334596, 0.00088398658074664654, 
    0.0009253613104477648, 0.00092556020154314922, 0.00088351114610354519, 
    0.00079965597550967697, 0.00067572454647910388, 0.00051444904750982175, 
    0.00031928129837902926, 9.4187433730680276e-05, -0.00015645472503143364, 
    -0.00042787127048162546, -0.00071485686689258272, -0.001011722994159484, 
    -0.0013122918316726307, -0.0016099177095623026, -0.0018975548071490734, 
    -0.0021678587242337779, -0.0024133326760651165, -0.0026265466453127273, 
    -0.0028004468985005251, -0.0029287658017345579, -0.0030065094451701396, 
    -0.0030304619325145716, -0.0029996386140829418, -0.002915606075157509, 
    -0.0027825956990482179, -0.0026073713086949878, -0.002398845367053544, 
    -0.0021674604062825406, -0.0019244151159727649, -0.0016808127738463317, 
    -0.0014468646866742441, -0.0012312180787239261, -0.0010405105616308323, 
    -0.00087915697176899434, -0.00074938225243609562, 
    -0.00065142236606294734, -0.00058386887964569046, 
    -0.00054406009436288628, -0.00052848671976638288, 
    -0.00053315398707896606, -0.00055387412820368941, 
    -0.00058646903607266086, -0.00062689125397801502, 
    -0.00067127133978263007, -0.00071592882813907208, 
    -0.00075737592361225972, -0.00079232871120620951, 
    -0.00081776011100078815, -0.00083097312255216204, -0.0008297065590494268, 
    -0.00081223772897034985, -0.00077751033230236285, 
    -0.00072524871039922171, -0.00065607429939662499, -0.0005716097158627965, 
    -0.00047452588046575239, -0.00036851855701770092, 
    -0.00025816756545405224, -0.00014867395525571857, 
    -4.5472339617945299e-05, 4.6229750390518461e-05, 0.00012194337603175506, 
    0.00017835400035021249, 0.00021366850333051177, 0.00022782839715583989, 
    0.00022254319067426185, 0.0002011471668064749, 0.00016830035654895941, 
    0.00012957007091215516, 9.0938101995865817e-05, 5.8291168172039901e-05, 
    3.6942065733158201e-05, 3.1247693173520347e-05, 4.4325985415987334e-05, 
    7.7912919468448532e-05, 0.00013233053816951977, 0.00020657673193091346, 
    0.00029848770845609663, 0.00040495281863218866, 0.00052212279626451621, 
    0.00064559460506573741, 0.00077054338182536489, 0.00089181957306907849, 
    0.0010040328826064482, 0.0011016522545860164, 0.0011791375813871795, 
    0.0012311149918265193, 0.0012525816684089168, 0.0012391236713095142, 
    0.0011871312655386801, 0.0010939824127675667, 0.00095818740397693284, 
    0.00077947563544036543, 0.0005588338187041403, 0.00029849310831209241, 
    1.8606682285627547e-06, -0.00032656112851705042, -0.00068127617856052344, 
    -0.001055909026942475, -0.0014433105533410823, -0.0018356909456860779, 
    -0.0022247678089818406, -0.0026019648052438412, -0.0029586461909046815, 
    -0.0032863977225774249, -0.0035773425108415616, -0.0038244997202887855, 
    -0.0040221455104874999, -0.0041661617699905789, -0.0042543151231400093, 
    -0.0042864198800832715, -0.0042643621204234783, -0.0041919691564934374, 
    -0.0040747716459445631, -0.0039196716984766303, -0.0037345646752090732, 
    -0.0035279441242605661, -0.0033085092977364703, -0.0030848018363617523, 
    -0.0028648822706828121, -0.0026560200942660544, -0.0024644057821287986, 
    -0.002294862104767374, -0.0021505796797686378, -0.0020329179913258833, 
    -0.0019413250721975128, -0.0018734165728227297, -0.0018252306277992696, 
    -0.0017916467877054838, -0.0017668971324293942, -0.0017451107274156338, 
    -0.0017208294686432456, -0.0016894454006831212, -0.0016475322646923778, 
    -0.0015930698984240347, -0.0015255495026231193, -0.0014459579932705449, 
    -0.0013566602063569838, -0.0012611895945071282, -0.0011639628661160751, 
    -0.0010699741210185914, -0.00098447842719028033, -0.00091268723648315405, 
    -0.00085949369417715317, -0.00082923433882650167, -0.0008254980031043496, 
    -0.00085099025418336005, -0.00090742996597436675, 
    -0.00099547223015736285, -0.0011146225068429506, -0.001263163221276788, 
    -0.001438084751929147, -0.0016350612633391466, -0.0018484973499781443, 
    -0.0020716561135491808, -0.0022968928475188841, -0.0025159698474691485, 
    -0.0027204580224275397, -0.0029021915496750868, -0.0030537632092122752, 
    -0.0031690106367044599, -0.0032434497556710334, -0.0032746181253164638, 
    -0.0032622660725162797, -0.0032083649978357147, -0.003116908488310496, 
    -0.0029935166078753498, -0.0028448683990927475, -0.0026780396662673088, 
    -0.0024998252654896817, -0.0023161320073284766, -0.002131536182406398, 
    -0.0019490441511263701, -0.0017700709946579141, -0.0015946282077753244, 
    -0.0014216800485552634, -0.0012495753086679631, -0.0010765347789837268, 
    -0.0009010720220525996, -0.00072232923307916021, -0.00054024143312773627, 
    -0.00035553556999873796, -0.00016955637213429318, 1.6026628771679422e-05, 
    0.00019952883978669906, 0.00037952080424956348, 0.00055495559879642758, 
    0.00072514429614459024, 0.00088959539974515535, 0.0010477442879363627, 
    0.0011986842450881232, 0.0013409496117031943, 0.0014724384974698804, 
    0.0015904740133450418, 0.0016920064287218991, 0.0017739047749950464, 
    0.0018332985817436044, 0.0018679405654441533, 0.0018765540272006513, 
    0.0018591295062664269, 0.0018171417643079615, 0.0017536197557125092, 
    0.0016730372326134407, 0.0015810075801716951, 0.0014837935701626297, 
    0.0013877024683392955, 0.0012984354132441545, 0.0012204929607396464, 
    0.0011566911691741539, 0.0011078798568214991, 0.0010728778905417118, 
    0.0010486398526340891, 0.0010306394983645086, 0.0010134168455976234, 
    0.00099122717588695682, 0.00095871600953726689, 0.00091155250664770853, 
    0.00084694478129652994, 0.00076400119427107453, 0.00066388477679203185, 
    0.00054974755986998745, 0.00042643039624702835, 0.0002999832997603978, 
    0.00017703149508380102, 6.4091217331295735e-05, -3.3088568486063724e-05, 
    -0.00011005836076920014, -0.0001640032862492114, -0.0001938637625727378, 
    -0.00020025421189555316, -0.00018523873939621418, 
    -0.00015201958269601601, -0.00010459857174028268, 
    -4.7455093665499448e-05, 1.4720622639917018e-05, 7.7253877139113621e-05, 
    0.00013563860985680364, 0.00018566991682734995, 0.00022355944013712661, 
    0.00024608800359920697, 0.00025079405265188907, 0.00023622428507864962, 
    0.00020218439427549517, 0.00014996225836468995, 8.2461587104318512e-05, 
    4.2037985201763777e-06, -7.8842368170696324e-05, -0.00015958758935596937, 
    -0.00023030684137090608, -0.00028323569798473322, 
    -0.00031124411138609194, -0.00030852177807341936, 
    -0.00027120903398228331, -0.00019790004422119581, 
    -8.9951617631567167e-05, 4.8444062250276066e-05, 0.00021045409316652701, 
    0.00038706324781662366, 0.0005677629011404282, 0.00074141620846785827, 
    0.00089718560913415023, 0.0010254660252042025, 0.0011186689129742309, 
    0.0011718131243122578, 0.001182825753476305, 0.0011525633392781484, 
    0.0010845459443361407, 0.00098448225015127303, 0.00085963545925728366, 
    0.00071811851072495279, 0.0005682011472812915, 0.00041767978273469635, 
    0.00027335753775502622, 0.00014067018109078451, 2.3485607050055934e-05, 
    -7.5931053753899676e-05, -0.00015679968406248534, 
    -0.00021956853340336673, -0.00026557541350764045, 
    -0.00029665717343062059, -0.00031476607007691542, 
    -0.00032163637033737392, -0.0003185487219192313, -0.00030620833716286537, 
    -0.00028475527924085291, -0.00025388154286729931, 
    -0.00021305505273453657, -0.00016175811012233586, 
    -9.9730861363945444e-05, -2.7172944458490778e-05, 5.5117544126753103e-05, 
    0.00014566434973323732, 0.00024227232160517606, 0.00034202890188338126, 
    0.00044132540098260916, 0.00053591524413535124, 0.00062099547754874485, 
    0.00069136350303554818, 0.00074163475021033582, 0.00076653279048326001, 
    0.00076126017788737436, 0.00072192585299425281, 0.0006459802712012033, 
    0.00053260421769898731, 0.00038299417436291847, 0.0002004766248041376, 
    -9.5898736795339122e-06, -0.00024011340954995016, 
    -0.00048274868877818555, -0.00072848681050815579, -0.0009682859075914016, 
    -0.0011936687094932872, -0.0013972384585426122, -0.0015730589542036998, 
    -0.001716913111283322, -0.0018264269880894925, -0.0019010697006992907, 
    -0.0019420436314945841, -0.0019520629822021734, -0.0019350273307982718, 
    -0.0018956281381795055, -0.0018388999112609135, -0.0017697580897105883, 
    -0.0016925681147933515, -0.0016107673624800388, -0.0015266076280906454, 
    -0.0014410407188228259, -0.001353797358410191, -0.0012636374596210038, 
    -0.0011687691240262214, -0.0010673256794222483, -0.00095786495074633735, 
    -0.00083976639312316828, -0.00071350891288554348, 
    -0.00058077377565121484, -0.0004444069806074338, -0.00030824265769560541, 
    -0.00017681848349972564, -5.5015104636547983e-05, 5.2352606096679833e-05, 
    0.00014096776492508343, 0.00020744248998605573, 0.00024969706345193853, 
    0.00026726558175041779, 0.00026146622869103862, 0.00023543867168140638, 
    0.00019399631391854406, 0.00014331862616808876, 9.0499600358284274e-05, 
    4.2965558024199046e-05, 7.8558105567620298e-06, -8.6034934494017504e-06, 
    -1.6392906362279855e-06, 3.1656693316130835e-05, 9.2099010795527504e-05, 
    0.00017837331562323497, 0.00028720913920768484, 0.00041370261838268805, 
    0.00055177340497797095, 0.00069467444923495983, 0.00083550668886109313, 
    0.00096770250752989439, 0.0010854321134070456, 0.0011839241473911603, 
    0.0012596873547047508, 0.0013106335428731122, 0.0013361153945140574, 
    0.0013368910204489362, 0.0013150141645117787, 0.0012736380515353939, 
    0.0012167429257614651, 0.0011487701913590242, 0.001074221065389412, 
    0.00099726090999811552, 0.00092138201111217465, 0.0008491771143854087, 
    0.0007822285615243041, 0.00072108623008099832, 0.00066534669142058597, 
    0.00061376791868968442, 0.00056442454789569637, 0.00051488138532214595, 
    0.00046235199145659467, 0.00040385356135024957, 0.00033636772120151291, 
    0.00025701789232156149, 0.00016326744617423556, 5.3148200878967974e-05, 
    -7.4495379703672513e-05, -0.00021976021928842148, -0.0003814956973262088, 
    -0.00055718302852530998, -0.00074296295332318928, 
    -0.00093382249518951022, -0.0011239537973054905, -0.0013072671348793872, 
    -0.0014779993654633202, -0.0016313262029948932, -0.0017638898247547615, 
    -0.0018741215531137181, -0.0019623121067188507, -0.0020303886357791465, 
    -0.0020814391819337927, -0.0021190706496139536, -0.0021467091968522881, 
    -0.002166955798543807, -0.0021810888632476772, -0.0021887985976991441, 
    -0.0021881600825867068, -0.0021758417890461951, -0.0021475287283604229, 
    -0.0020984783221400876, -0.0020241545154080286, -0.0019208568495718734, 
    -0.0017863038428402747, -0.0016200918968089038, -0.0014240220992373144, 
    -0.0012022202927213042, -0.00096107287848435535, -0.00070890278308267018, 
    -0.00045543706174952856, -0.00021107459445968713, 1.3955596340866159e-05, 
    0.00021044746445142372, 0.00037098622431441385, 0.0004905497354620172, 
    0.00056686319465916522, 0.00060052185248116749, 0.00059487898910860239, 
    0.00055573125543782894, 0.00049085599364883184, 0.0004094440989568821, 
    0.00032148003823781322, 0.00023710868668735578, 0.00016604383048683137, 
    0.00011705274668387593, 9.7557714736833413e-05, 0.00011338252755541299, 
    0.00016864321239630752, 0.00026576498974896371, 0.0004055734034740904, 
    0.00058742078959760568, 0.00080930841737917388, 0.0010679747240865847, 
    0.0013589625750500482, 0.0016766461523859254, 0.0020142550674216823, 
    0.0023639119776495219, 0.0027167330842696219, 0.0030630132819949966, 
    0.0033925221661161424, 0.0036949134517028663, 0.0039602152777642053, 
    0.0041793691409899442, 0.0043447430064149735, 0.0044505842587788365, 
    0.004493328373840322, 0.0044717584129455572, 0.0043869985534339476, 
    0.0042423619679210645, 0.0040430846004874061, 0.0037959973544849524, 
    0.0035091695677824169, 0.0031915463902771101, 0.0028526030041745769, 
    0.0025020156266567575, 0.002149332751511474, 0.0018036726102087376, 
    0.0014734214645382273, 0.001165964931577981, 0.00088747169384252914, 
    0.00064275870900428367, 0.00043524930145796272, 0.00026703839689915047, 
    0.00013903715036113313, 5.1172240159931747e-05, 2.5728062033592893e-06, 
    -8.2747594606131475e-06, 1.6540017562920601e-05, 7.4330191351262717e-05, 
    0.00016174217225646775, 0.00027463416631030824, 0.00040795535103578068, 
    0.00055566719225849919, 0.00071072364775015963, 0.00086515873835023803, 
    0.0010102904102522253, 0.0011370406175852329, 0.0012363625762266848, 
    0.001299759551864969, 0.0013198265851630886, 0.0012907788858435923, 
    0.001208920449741691, 0.0010730061290191821, 0.00088447054284675349, 
    0.00064749768920841801, 0.00036891535003519445, 5.791628130975316e-05, 
    -0.00027441276592635942, -0.00061571080084418188, 
    -0.00095308271497468618, -0.001273887818034935, -0.0015665072313225132, 
    -0.0018210193516079881, -0.002029702550137613, -0.0021873508453280083, 
    -0.0022913659338404751, -0.0023416452841011847, -0.0023402999934425536, 
    -0.0022912534254567584, -0.0021997744262824536, -0.0020719953189052209, 
    -0.0019144667746354485, -0.0017337817903327493, -0.001536277307771033, 
    -0.0013278138469492069, -0.0011136431889799932, -0.00089833513101821786, 
    -0.00068576708036329544, -0.00047915471558127422, 
    -0.00028113166325422612, -9.3860447250328785e-05, 8.0825556846630478e-05, 
    0.00024127654029921003, 0.00038588597613303674, 0.00051297659138169107, 
    0.00062075342126976672, 0.00070732766131803679, 0.00077083131866937586, 
    0.00080959879049266104, 0.00082241485279761295, 0.00080875716263364907, 
    0.00076901280974406424, 0.00070461705533957661, 0.00061809045443266897, 
    0.00051295855629756584, 0.00039356980903681749, 0.00026482335721797115, 
    0.00013184049643016787, -3.9757836268134163e-07, -0.00012742149936895901, 
    -0.00024562845521554339, -0.00035259308681557172, 
    -0.00044729367468539742, -0.00053020943276387348, 
    -0.00060325019415914173, -0.00066950040299630002, 
    -0.00073279965519437327, -0.0007972052593199101, -0.00086643583005525352, 
    -0.00094336721181298834, -0.0010296616364709672, -0.0011255794493931701, 
    -0.0012299716312697202, -0.0013404495575454944, -0.0014536761553208025, 
    -0.0015657394544445755, -0.0016725523495780914, -0.0017702578186258005, 
    -0.001855570299463814, -0.0019260323505410784, -0.0019801408042117385, 
    -0.0020173252761950303, -0.0020378077445981821, -0.002042364442699578, 
    -0.0020320637744514827, -0.0020080163494641174, -0.0019711715137070806, 
    -0.0019222168565881965, -0.0018615624571376658, -0.0017894148373270938, 
    -0.001705929791873865, -0.0016113718997522897, -0.0015062658624489078, 
    -0.0013914776391184621, -0.0012681984168995597, -0.0011378528360338378, 
    -0.0010019164758145063, -0.00086169292051280634, -0.00071808203892822576, 
    -0.00057138990188976366, -0.00042120206028519879, 
    -0.00026636653445666754, -0.00010508893620814093, 6.4856525269997613e-05, 
    0.0002457926336447886, 0.00043972946662500765, 0.00064788427326329268, 
    0.00087022265040347731, 0.0011050503104263064, 0.001348742747567751, 
    0.0015956742104347593, 0.0018383570126807504, 0.0020678155211954203, 
    0.0022741571965920306, 0.0024472505051985269, 0.0025774733533719739, 
    0.0026564163113603299, 0.0026775064513569861, 0.0026365151476501667, 
    0.0025319371220403849, 0.0023652249668324561, 0.0021408556752747793, 
    0.0018662095887920528, 0.0015512404724816573, 0.0012079554677895965, 
    0.00084974092193916973, 0.00049059783805609561, 0.0001443616761083465, 
    -0.00017601097108209588, -0.00045904954818133176, 
    -0.00069523670511497575, -0.00087733090447069469, -0.001000546139390735, 
    -0.0010626218296080582, -0.0010637788479202607, -0.0010065993104446465, 
    -0.000895837988780692, -0.00073816333579698897, -0.00054186471148971955, 
    -0.00031649684817706308, -7.2498019589221978e-05, 0.00017920067907259879, 
    0.00042755453250131276, 0.00066175725469800619, 0.00087155891544414999, 
    0.0010475864046125371, 0.0011816709064715895, 0.0012672018239614732, 
    0.0012994850468357388, 0.0012760749027690768, 0.0011970024968526974, 
    0.0010648551654364416, 0.00088465833794731138, 0.00066355955353983895, 
    0.00041032161745089781, 0.00013466885056808721, -0.00015343932367870873, 
    -0.00044451356927566616, -0.00073016581174658191, -0.001003587847774983, 
    -0.0012598420760172604, -0.0014959720901439641, -0.0017109407806163376, 
    -0.0019054326248959654, -0.0020815463317346884, -0.002242421205943155, 
    -0.0023918066013508201, -0.0025336083499326776, -0.0026714542281017113, 
    -0.0028082872699321214, -0.0029460324136621192, -0.0030853629094038794, 
    -0.0032255899118806587, -0.0033646906784716639, -0.003499474166079214, 
    -0.0036258820758235232, -0.0037393938278455496, -0.0038354854451761464, 
    -0.0039101013628382976, -0.0039600636427215294, -0.0039833688776312708, 
    -0.003979331415010918, -0.0039485474158340019, -0.0038926944859546814, 
    -0.0038142107593219093, -0.0037159291107639945, -0.0036007431095213599, 
    -0.0034713575876055064, -0.0033301880800827776, -0.003179395713653286, 
    -0.0030210343498086969, -0.002857264362401414, -0.0026905727426401742, 
    -0.0025239387070130582, -0.0023609036342515273, -0.0022055345754557702, 
    -0.0020622838154557735, -0.0019357678419894774, -0.0018304754439371288, 
    -0.0017504266267421402, -0.0016987900729313527, -0.0016774821248065844, 
    -0.0016867798546336239, -0.0017250375946883615, -0.0017885344479402084, 
    -0.0018715239992983205, -0.001966508597711573, -0.002064717613721981, 
    -0.0021567669688606649, -0.0022334168354502921, -0.002286350934466011, 
    -0.0023088695913620742, -0.0022964554511935055, -0.0022471211073501057, 
    -0.0021615297495145196, -0.0020428910327341702, -0.0018966577001289732, 
    -0.001730081009899341, -0.001551662905459556, -0.0013705390949428969, 
    -0.0011958212203240094, -0.0010359255360190189, -0.00089795378333373506, 
    -0.00078716585967806977, -0.00070658924145473401, 
    -0.00065681697519964365, -0.00063598569238281139, 
    -0.00063994914677961137, -0.00066263900218633761, 
    -0.00069658279559876488, -0.00073356817412874428, -0.0007653970708465977, 
    -0.0007846495639549266, -0.00078540467560932073, -0.00076378901845085192, 
    -0.00071832317893734789, -0.00064996839459518347, 
    -0.00056187139662772256, -0.00045885270290505056, 
    -0.00034667800818652606, -0.00023125101614154806, 
    -0.00011784779080637706, -1.0509794219409146e-05, 8.8297337570369605e-05, 
    0.00017771324169611855, 0.00025822201565620253, 0.00033116861477856693, 
    0.00039817638187289797, 0.00046058532593655044, 0.00051904070409951428, 
    0.00057328871140563886, 0.00062220991999601338, 0.00066404279794922373, 
    0.00069675245521975526, 0.00071842879825984799, 0.0007276448172739827, 
    0.0007237372019949169, 0.00070696236120083562, 0.00067855611773113189, 
    0.00064069216546420614, 0.0005963618537638154, 0.00054918275865183542, 
    0.00050314991009328539, 0.0004623558827570876, 0.00043071543481333445, 
    0.00041172367041145439, 0.0004082678794627153, 0.00042252242153687327, 
    0.00045588658539805226, 0.00050893709088841701, 0.00058138913379822627, 
    0.00067203917392341065, 0.00077871655984213244, 0.00089826363507770532, 
    0.0010265717384236807, 0.0011586768590147118, 0.0012889312683268053, 
    0.0014112533140966748, 0.0015194373413691805, 0.0016075317995203999, 
    0.0016702433547443954, 0.0017033542305054221, 0.0017040780134320601, 
    0.0016713133887703731, 0.0016057378097816927, 0.0015097246261017298, 
    0.0013870668674601156, 0.0012425652076849516, 0.001081540997427166, 
    0.00090937564042551787, 0.00073112324362643638, 0.00055129284283418102, 
    0.00037377513183476708, 0.00020192692099105602, 3.8745564673012175e-05, 
    -0.00011291028287482411, -0.00025014130229969673, -0.0003699144212439393, 
    -0.00046910340533127854, -0.00054464638160714104, 
    -0.00059380989336166323, -0.00061452795923930411, 
    -0.00060576820232511209, -0.00056788523846214517, 
    -0.00050291430053289894, -0.00041471641898587348, 
    -0.00030893573109912653, -0.0001927143320570089, -7.4159866493158033e-05, 
    3.8371536247023913e-05, 0.00013709689792319263, 0.00021562882303721883, 
    0.00026966964756857916, 0.00029748733202287863, 0.0003000990185545371, 
    0.00028115100410838024, 0.00024651069954023663, 0.00020362674801258107, 
    0.00016072574458509927, 0.0001259529520922019, 0.00010653289768368128, 
    0.00010803424869829788, 0.00013381298513817145, 0.00018467960899643085, 
    0.00025885033315381999, 0.00035215047751882366, 0.00045850834311617945, 
    0.00057063203934375477, 0.00068084126286161405, 0.00078188760381836975, 
    0.00086769516877505332, 0.00093391418064347337, 0.00097825399918209286, 
    0.0010005970148584389, 0.0010029073262940778, 0.00098899673412802618, 
    0.00096417062451514498, 0.00093477628623009454, 0.0009076542152560848, 
    0.00088950318201248574, 0.00088617697504809979, 0.00090198258318968942, 
    0.00093904990527634766, 0.00099687236642193272, 0.0010721115990375174, 
    0.0011587016523246937, 0.0012482682529239369, 0.0013308229635139739, 
    0.0013956579958595706, 0.0014323324898694193, 0.0014316343718471182, 
    0.0013864391323433222, 0.0012923568149774271, 0.0011481355089342491, 
    0.00095579646647156913, 0.00072048483787766652, 0.00045007169763457638, 
    0.00015455586237224578, -0.00015466523614889103, -0.00046556364017068767, 
    -0.00076622910741282299, -0.0010455192036595529, -0.0012935878557787635, 
    -0.0015022327527963915, -0.0016651094112571545, -0.0017777701823552137, 
    -0.0018375916375718043, -0.0018436081247680883, -0.0017963090016817093, 
    -0.0016974613004610178, -0.0015499757650012497, -0.0013578429472362534, 
    -0.0011261452124881439, -0.00086109182723151725, -0.00057002735521506805, 
    -0.00026135571306722452, 5.567007145955707e-05, 0.00037129942256305151, 
    0.00067577013554816071, 0.00095988126177848614, 0.0012155801533360407, 
    0.0014364977482590141, 0.0016183634122265852, 0.0017592696720042658, 
    0.0018597553224405045, 0.0019227007599510993, 0.0019530716977671457, 
    0.0019575057084455869, 0.0019438052538745562, 0.0019203683470850022, 
    0.0018955906191116031, 0.0018772933272221753, 0.0018722375960078088, 
    0.0018857639876532495, 0.0019215665537426021, 0.0019816349205061395, 
    0.0020663256877502165, 0.0021745395251681621, 0.0023039403849433324, 
    0.0024511850694576209, 0.0026121608569531314, 0.0027822250850012315, 
    0.0029564467068955414, 0.0031298833322637122, 0.0032978515695220598, 
    0.0034561951288722796, 0.0036015077274189292, 0.003731294779612127, 
    0.0038440400402646934, 0.0039392035140436623, 0.0040171095157627984, 
    0.0040787926268339523, 0.0041257976515841821, 0.0041599717679562977, 
    0.0041832874136905418, 0.0041976738186201342, 0.0042049061369119171, 
    0.0042065067489501021, 0.0042036552506389928, 0.0041970921300546853, 
    0.0041870007282990718, 0.0041728797247736317, 0.0041534506976048519, 
    0.004126646624848648, 0.0040897224006959318, 0.0040394899666256322, 
    0.0039726446230497411, 0.0038861473969937312, 0.0037775614074456935, 
    0.0036453083072426171, 0.0034888312119570192, 0.0033086227774387356, 
    0.0031061717914695761, 0.002883857929723403, 0.0026448183232912104, 
    0.0023928077145817695, 0.0021320468175185978, 0.0018670343958215384, 
    0.0016023194247838026, 0.0013422060455409298, 0.0010904307918719071, 
    0.00084984138395679425, 0.00062214888346586751, 0.00040779650964817152, 
    0.00020599791290920851, 1.4944535180388097e-05, -0.00016779826608081204, 
    -0.00034479623086318482, -0.00051819447801886693, 
    -0.00068919009003237989, -0.00085762613060222598, -0.0010217635375362223, 
    -0.0011782568312921765, -0.0013223510245691248, -0.0014482754033008688, 
    -0.0015498109137943349, -0.0016209751372473244, -0.001656701629525365, 
    -0.0016534371215132107, -0.0016095424391349609, -0.0015254750602973438, 
    -0.001403682760698318, -0.0012482427864873628, -0.001064344542580813, 
    -0.00085765413378912736, -0.00063372490978921088, 
    -0.00039755936141786961, -0.0001533683528064443, 9.5418674626217886e-05, 
    0.0003459561184839173, 0.00059565406686319623, 0.00084185725880323156, 
    0.0010815893134426247, 0.0013114451679502013, 0.0015276612483429276, 
    0.0017263411058643418, 0.0019038489938272638, 0.0020572674553921162, 
    0.0021848846932289181, 0.0022865990745641949, 0.0023641694319660347, 
    0.002421278500236935, 0.0024633956100132467, 0.0024974934937565703, 
    0.0025316781046506214, 0.002574769508289203, 0.002635854948576349, 
    0.0027238466887719343, 0.002846995369028881, 0.0030123807904203844, 
    0.0032253703034584749, 0.0034890725020077767, 0.0038038357838921103, 
    0.0041668877713896563, 0.0045721372230129956, 0.0050102153927904843, 
    0.005468742944647588, 0.0059328156996929044, 0.0063856528884758913, 
    0.006809343494057791, 0.0071856625271769234, 0.0074968776243727938, 
    0.0077265463289878039, 0.007860260146294042, 0.007886324193649737, 
    0.007796353562983872, 0.0075857646445718499, 0.0072541245684981433, 
    0.0068053512547261216, 0.0062477183714389449, 0.0055936371973736637, 
    0.004859227575233196, 0.0040636359595360074, 0.0032281253912812891, 
    0.0023749736665767238, 0.0015262792140699497, 0.0007028215057869573, 
    -7.6939332979640419e-05, -0.00079759740008481168, -0.0014472816189058438, 
    -0.0020178505624176822, -0.0025048319318075811, -0.0029071484349568705, 
    -0.0032266262916110611, -0.0034674259966929232, -0.0036353946583393354, 
    -0.0037374715919960967, -0.0037811934968889475, -0.0037743063285267404, 
    -0.0037244641811445991, -0.0036389996740168909, -0.0035247496558960261, 
    -0.0033879164935755818, -0.003233973806885811, -0.0030675972537001872, 
    -0.0028926202022475692, -0.0027120149291611985, -0.0025278881881310375, 
    -0.0023414596308328709, -0.0021530553195760298, -0.0019620725418456109, 
    -0.0017670030465692082, -0.0015654908090351996, -0.0013545315216123091, 
    -0.0011307506054375055, -0.00089079394434302117, -0.0006318052237106541, 
    -0.00035192127230606885, -5.0713436503869109e-05, 0.00027047139007254067, 
    0.00060834858247764184, 0.000957748976826819, 0.0013118716289707828, 
    0.0016627220679934344, 0.0020016736413508347, 0.0023201251596822086, 
    0.002610150735161671, 0.0028651002042245862, 0.0030800933336274433, 
    0.0032523473770263156, 0.0033812696155234804, 0.0034683446311307427, 
    0.003516750195098727, 0.0035307807820063376, 0.0035151299729499728, 
    0.0034741153985533299, 0.003411017729938349, 0.0033276165354911261, 
    0.0032240915579171713, 0.0030992931348616868, 0.0029513213838665425, 
    0.0027782786498675928, 0.0025790447303485394, 0.0023538671801721102, 
    0.0021046946649965785, 0.0018351855163893369, 0.0015503873834959035, 
    0.0012561430072689722, 0.00095831355318128238, 0.0006619704734347453, 
    0.00037065533014711218, 8.5958471583207576e-05, -0.00019250916217259539, 
    -0.00046669889469823204, -0.00073928298319795118, -0.0010125954141204784, 
    -0.0012875477378411024, -0.001562734788717214, -0.0018338870327666563, 
    -0.0020937272773592932, -0.0023322308393095219, -0.0025372972706105661, 
    -0.0026957689594672286, -0.0027947028170829859, -0.0028227587410558351, 
    -0.0027715028938730653, -0.0026364308725894941, -0.0024175611497909118, 
    -0.0021194825222711775, -0.0017509070495722418, -0.0013237993699898479, 
    -0.00085228537438978734, -0.00035150617129787602, 0.00016339603943417433, 
    0.00067808015086930312, 0.0011795338602841828, 0.0016563860398575529, 
    0.0020990653797764236, 0.0024999069376673484, 0.0028532631898867235, 
    0.0031556091207029101, 0.0034056711322674564, 0.0036044596201832597, 
    0.0037551893358923581, 0.003863006362138256, 0.0039345268497011296, 
    0.0039772140940996323, 0.0039986519608301539, 0.0040058111673858064, 
    0.0040043852018618997, 0.0039982685121038924, 0.0039892318745216532, 
    0.0039768113139897589, 0.0039584129063127867, 0.0039295830579986315, 
    0.0038844310088575677, 0.0038161003417812363, 0.0037173004368602747, 
    0.0035808230450287428, 0.0034000739306094107, 0.0031696057838124787, 
    0.0028855952118704126, 0.0025462725927739194, 0.0021521970946870722, 
    0.0017063632246270596, 0.0012141412769327588, 0.00068306416946401773, 
    0.00012251102000670271, -0.00045666087722431869, -0.0010425010311988219, 
    -0.0016223319158798395, -0.0021831206097704123, -0.002711842072127736, 
    -0.0031958625992986435, -0.0036233805553226128, -0.0039838909796824779, 
    -0.004268673705101267, -0.0044712529032466019, -0.0045878090704268119, 
    -0.0046174714013318208, -0.0045624365002618567, -0.0044279042584578288, 
    -0.0042217697444924505, -0.0039540931252157567, -0.0036363906180050458, 
    -0.0032808324189380418, -0.0028994737960101082, -0.002503647117823183, 
    -0.0021035671864047729, -0.0017081956292157535, -0.0013252885575882835, 
    -0.00096154908778878071, -0.00062275168780713856, 
    -0.00031380301914419787, -3.8719494918042197e-05, 0.0001994398288674336, 
    0.0003986100614270834, 0.00055771334267450557, 0.00067661425184197585, 
    0.00075609639517704727, 0.00079791549477898846, 0.00080488294351881129, 
    0.00078099514076927085, 0.00073146813837456483, 0.0006626372995117497, 
    0.00058167745453831926, 0.00049615357138194809, 0.00041347220820930398, 
    0.00034036441404985577, 0.00028244124336099154, 0.00024390378704998005, 
    0.00022739663525687942, 0.0002340048324372452, 0.00026341531133364661, 
    0.0003141826340131659, 0.0003840917654848343, 0.00047049027734962135, 
    0.00057059990660402588, 0.00068170973334488185, 0.00080128600565389728, 
    0.00092700676203482236, 0.0010567604092099753, 0.0011886382403768056, 
    0.0013209372337303071, 0.0014521813725747309, 0.0015811521393781947, 
    0.0017069221211816876, 0.0018288633461929571, 0.0019466686394009147, 
    0.002060351975245618, 0.0021701913109646326, 0.00227662908298158, 
    0.0023800622751462574, 0.0024806194310433112, 0.0025778930699982064, 
    0.0026707761779352097, 0.0027574313923772091, 0.0028354278013202126, 
    0.0029019674519290212, 0.0029541712103648941, 0.002989379693360804, 
    0.003005408028574815, 0.0030007273007387936, 0.0029745861707178656, 
    0.0029270287846427301, 0.0028588484810835048, 0.0027714262657077132, 
    0.0026665328015767036, 0.0025460952163062862, 0.0024119940930356788, 
    0.0022659304535144059, 0.0021093730330227489, 0.0019436009632716174, 
    0.0017697986687633491, 0.0015891876409302741, 0.001403150184075443, 
    0.0012133664984500063, 0.0010219198762884288, 0.00083139201876282899, 
    0.00064494200636864218, 0.0004663180695578171, 0.00029983470604647689, 
    0.00015023274580823432, 2.2446985003710095e-05, -7.8716033823454098e-05, 
    -0.00014893915321476664, -0.00018481364580518801, 
    -0.00018421224872268297, -0.00014664344017010166, 
    -7.3544180355008312e-05, 3.1499485494167794e-05, 0.00016263419788700812, 
    0.00031170049072244319, 0.00046837121826619015, 0.00062048910172151804, 
    0.00075466892562119623, 0.00085715743562642219, 0.00091494446738642535, 
    0.00091700208170061512, 0.00085557509455352931, 0.00072733481820890455, 
    0.00053422740205390695, 0.00028387442626974703, -1.0616198700588033e-05, 
    -0.000331488688355614, -0.00065774810599632727, -0.00096695918071388904, 
    -0.0012371615895516192, -0.0014486353910315381, -0.0015854028720524176, 
    -0.0016363615901759817, -0.0015960307368254763, -0.0014649221247451691, 
    -0.0012495529053303646, -0.00096208757929887442, -0.00061963775522884423, 
    -0.00024319348503673368, 0.00014382989038057477, 0.0005173325264806346, 
    0.0008544808317160899, 0.0011356071521820197, 0.0013459044994250356, 
    0.0014766702803011447, 0.0015259267961558226, 0.0014984282341555914, 
    0.0014049886224299891, 0.0012612678642605602, 0.0010861307193004831, 
    0.00089971837278924965, 0.00072150601061882994, 0.00056851416759734128, 
    0.00045391019846152041, 0.00038608839345420507, 0.00036837231018640787, 
    0.00039919946441335427, 0.00047279794737324952, 0.00058017923789238646, 
    0.00071027168107625101, 0.00085111929876955652, 0.00099095672838021972, 
    0.0011191704455351973, 0.0012270416258274219, 0.0013083376720268857, 
    0.0013596942925694162, 0.0013807953598119857, 0.0013742934904287863, 
    0.0013454420779759366, 0.001301533822703759, 0.0012511981878367668, 
    0.0012036850678575977, 0.0011681867807632051, 0.0011532563925560121, 
    0.0011662803600997237, 0.001213066015451939, 0.0012974879997244418, 
    0.0014212198374584429, 0.0015835547395289852, 0.0017813359832841782, 
    0.0020090361015966405, 0.0022589702874362149, 0.002521728516379617, 
    0.0027867684206211189, 0.0030431752954258504, 0.0032805104055895606, 
    0.0034896217896730444, 0.0036633509601863507, 0.0037970284503555116, 
    0.0038886859661076503, 0.0039389888452192479, 0.0039508717880648555, 
    0.0039289706935444948, 0.0038789966716290809, 0.0038071017479195139, 
    0.003719353310509444, 0.00362132481952752, 0.0035177875850802422, 
    0.0034126062907188434, 0.0033087841313041407, 0.0032087195128438417, 
    0.0031145467075083294, 0.003028468480922396, 0.0029529295065138278, 
    0.0028905418425762019, 0.0028437641599536852, 0.0028143626368137336, 
    0.0028028451333973934, 0.0028079594926360613, 0.0028264999285239705, 
    0.0028534496972117324, 0.0028824395893966726, 0.0029064630774834487, 
    0.0029186342674430562, 0.0029128443289893969, 0.0028842786818643975, 
    0.0028297111867765646, 0.002747617965501901, 0.0026381603657107482, 
    0.0025030895592548265, 0.0023455990935755573, 0.0021700918020436753, 
    0.001981947574787089, 0.0017871585487476912, 0.0015919390209862428, 
    0.0014023199079462292, 0.0012238087957249322, 0.0010611855837156558, 
    0.0009185123424584195, 0.00079931806852822306, 0.00070691383398630285, 
    0.00064475366221386195, 0.00061666597022981356, 0.000626932264535586, 
    0.00068010227734104436, 0.00078059187861183972, 0.00093213809687679153, 
    0.0011371051538050466, 0.0013958314737196086, 0.0017060569746952063, 
    0.0020625912671103299, 0.0024572448311255754, 0.0028790739899809533, 
    0.003314899932346343, 0.0037499836549677139, 0.0041688737430186978, 
    0.0045562826732208368, 0.0048979313339594316, 0.0051813814607557639, 
    0.0053967200253598599, 0.0055371482391569759, 0.0055994292277575389, 
    0.0055841667946766003, 0.0054959250892468812, 0.0053430920298665899, 
    0.0051375156618458607, 0.0048938223023237649, 0.0046285357595370162, 
    0.0043590345416112683, 0.0041024648844942609, 0.0038747203407003016, 
    0.0036896128331957256, 0.0035582525032115645, 0.0034886348527753187, 
    0.0034854125267161891, 0.0035498402764905248, 0.003679803271076467, 
    0.0038700035622169591, 0.0041122432382555965, 0.0043958237152279976, 
    0.0047080676761414317, 0.0050349347245318855, 0.0053617087948421753, 
    0.0056737695322372382, 0.0059573874543886896, 0.0062004983416665913, 
    0.0063933396083486827, 0.0065289625632094341, 0.0066034689572017167, 
    0.0066160599343951538, 0.0065688304968071487, 0.006466370562204597, 
    0.0063152067644219254, 0.0061231333713873291, 0.0058985101675003947, 
    0.0056496372371610034, 0.0053842162755280854, 0.0051089738302475237, 
    0.0048295083984048288, 0.004550314340046803, 0.0042749715308943595, 
    0.004006479220690572, 0.0037476494104093719, 0.0035014773156026536, 
    0.0032714437123359829, 0.0030616689081573831, 0.0028768784187027841, 
    0.002722165418536648, 0.0026025253545190535, 0.002522232341704823, 
    0.0024840643373900814, 0.0024886206428492725, 0.002533770450575532, 
    0.0026143638938663787, 0.0027223935973160209, 0.002847446226980084, 
    0.0029775403394405242, 0.0031000858798465908, 0.0032029639848665009, 
    0.003275392234312789, 0.0033085782791209828, 0.0032959865611338875, 
    0.003233267742642897, 0.0031178288916019685, 0.0029482478702863892, 
    0.0027236948872622858, 0.0024435088976567966, 0.0021071198073481174, 
    0.0017143520805493933, 0.001266027497151333, 0.00076475171868268231, 
    0.00021560660671703853, -0.0003733309393590413, -0.00099095980211214908, 
    -0.0016234957904327847, -0.0022553532178671795, -0.0028703007019893669, 
    -0.0034529138852967987, -0.0039899752035922496, -0.0044716779340064289, 
    -0.0048923258512756944, -0.005250469495904006, -0.0055483907672810202, 
    -0.0057911325780996593, -0.0059852093152869554, -0.0061372636533509571, 
    -0.0062529314604184228, -0.0063360167016113349, -0.00638806446582698, 
    -0.0064084145449064206, -0.0063945940707388583, -0.0063430952033301565, 
    -0.0062503383980816807, -0.0061136733156646524, -0.0059322925265392554, 
    -0.0057077449089761702, -0.0054440821707173138, -0.0051475132867408804, 
    -0.0048256881526082974, -0.004486786302874874, -0.0041385590596876654, 
    -0.0037875511468106774, -0.0034385033503068875, -0.003094131634345001, 
    -0.0027551625506055302, -0.0024206445175332389, -0.0020885173968652115, 
    -0.0017562399523778712, -0.0014215575484012196, -0.0010830815860704808, 
    -0.00074085713778542493, -0.00039661609970084006, 
    -5.3829324477431295e-05, 0.00028248734107207683, 0.00060616453464057603, 
    0.00091046925268395917, 0.0011887923005601863, 0.0014353094813616962, 
    0.00164558530050027, 0.0018170164257005552, 0.0019491437777408955, 
    0.0020437125640471523, 0.0021045860697536142, 0.0021375734443649709, 
    0.0021500657673751387, 0.0021506433618199063, 0.0021485975543923692, 
    0.0021532835204242152, 0.002173406461660267, 0.0022162113621316368, 
    0.0022867340778956672, 0.0023869863798547195, 0.0025154629864407689, 
    0.0026668258220287522, 0.0028320212057003809, 0.0029987272638850333, 
    0.0031521986910534473, 0.0032764807283769087, 0.0033557557519004202, 
    0.0033758498455712404, 0.0033256916558165547, 0.0031986795353296099, 
    0.0029937026581037351, 0.0027157224364203845, 0.0023757359278261713, 
    0.001990018625979386, 0.0015787058818884309, 0.0011638226515037827, 
    0.00076709305370055263, 0.00040767294964259366, 0.00010023812728017357, 
    -0.00014635191648764369, -0.00032966860853204596, 
    -0.00045353420843879472, -0.00052712020975540603, 
    -0.00056334302471735208, -0.00057686707126114933, 
    -0.00058188047875688375, -0.00058983130597223201, 
    -0.00060761421940631736, -0.00063644451274556455, 
    -0.00067175164672301786, -0.0007040270573904139, -0.00072025995208706544, 
    -0.0007055476910465899, -0.0006446528725998484, -0.00052341388161702778, 
    -0.00033007379932137977, -5.6348001913304574e-05, 0.00030173131820110388, 
    0.00074342356139975795, 0.0012632213238629229, 0.0018511709059075498, 
    0.0024935301559849011, 0.0031736334391062808, 0.0038728750159037467, 
    0.0045716745662063973, 0.0052502625040712382, 0.0058893355627102247, 
    0.0064705696882714639, 0.0069772599593989158, 0.0073949693480249504, 
    0.0077123084223605365, 0.0079215928746267216, 0.0080192944317841429, 
    0.0080060502376373219, 0.0078862437809088838, 0.0076672396364364853, 
    0.0073584936294027658, 0.0069704863225840156, 0.006513885915548732, 
    0.0059988660333590476, 0.0054347534022476073, 0.0048298456126467902, 
    0.0041915512938369868, 0.0035265516303143092, 0.0028410218049404875, 
    0.0021407766432471002, 0.0014314454115589787, 0.00071870328663530328, 
    8.6196795479700495e-06, -0.00069196894185373633, -0.0013752498400158156, 
    -0.0020324824486464672, -0.0026543245843057462, -0.0032313409912030295, 
    -0.0037544893234609735, -0.0042154784493388976, -0.0046068989189167967, 
    -0.0049220233732518636, -0.0051544323929300336, -0.0052974555819574245, 
    -0.0053436291014130836, -0.0052845393760154293, -0.0051111918796176272, 
    -0.0048148835440347398, -0.0043885625575183964, -0.0038283696459952489, 
    -0.0031350676575349944, -0.0023151650187278822, -0.0013814130499384756, 
    -0.00035269328681518765, 0.00074667204792604463, 0.0018883069754426361, 
    0.0030416005649402493, 0.0041757669926101477, 0.0052619659722017084, 
    0.0062752753524919214, 0.0071962526378592656, 0.0080118129959306384, 
    0.0087153783237562555, 0.0093061163863984303, 0.0097876049051572878, 
    0.010165967455385404, 0.010448076034499433, 0.010640084367050049, 
    0.01074648323103539, 0.010769823838350429, 0.010710696619625665, 
    0.010567816496467694, 0.01033790164336657, 0.010015309440330552, 
    0.0095918500254085701, 0.0090569622895018392, 0.0083986483071701191, 
    0.007604858148295428, 0.0066655874052395812, 0.0055749497690043169, 
    0.0043334407175046521, 0.0029498236504045599, 0.0014424135982526614, 
    -0.00016050656797181033, -0.0018215416584072149, -0.003496380751817687, 
    -0.0051370770384632286, -0.0066961457601291746, -0.0081305401554407266, 
    -0.0094049640417148764, -0.010493615913283849, -0.011380249706590588, 
    -0.012056740562311184, -0.012520942963857805, -0.012775020529234689, 
    -0.012824781898257587, -0.012680150339354511, -0.012355896720009828, 
    -0.011872145773574904, -0.011254127499064983, -0.01053116109605543, 
    -0.0097351505305839324, -0.0088990618352364874, -0.0080551228580481096, 
    -0.0072333677014318693, -0.0064602247977054647, -0.0057575795388936637, 
    -0.0051419491749799392, -0.0046239623301302189, -0.0042081349850813903, 
    -0.0038928582387191177, -0.0036706590629910297, -0.0035286439193331258, 
    -0.0034491924723501093, -0.0034110834824511542, -0.0033908483023886793, 
    -0.0033644687631744349, -0.0033093117540687312, -0.0032061252549983889, 
    -0.0030411817838694923, -0.0028086246064099132, -0.0025122829651182494, 
    -0.0021668200438349329, -0.0017972931097567665, -0.0014368750185715518, 
    -0.0011224566053359161, -0.00088872770122701869, -0.0007618944387056181, 
    -0.0007542153274949536, -0.00086131564890173809, -0.0010630951482872688, 
    -0.0013279217150700779, -0.0016192953351488527, -0.0019033990119816471, 
    -0.0021565329907752531, -0.0023706002582639897, -0.0025569478553566344, 
    -0.0027471975782948467, -0.0029920664900301157, -0.0033561646796666407, 
    -0.0039101878855535678, -0.0047196012115384009, -0.0058322096762083589, 
    -0.0072668224510637827, -0.0090056044612758287, -0.010993261460563529, 
    -0.013143048325747851, -0.015347665776179364, -0.017494726458162701, 
    -0.019482967727729245, -0.021234274289279913, -0.02270198758747052, 
    -0.023872107706858176, -0.024760313480756101, -0.025407019930365198, 
    -0.025870921294734346, -0.02622422284214751, -0.026546896104964388, 
    -0.026920198305524227, -0.027418957668548929,
  // Fqt-total(9, 0-1999)
    0.99999999999999944, 0.99040669518327629, 0.96222899527673156, 
    0.9172037856185381, 0.85800909162886374, 0.78797875978805598, 
    0.71077020720158313, 0.6300339434217187, 0.54912725863559297, 
    0.47090151033659094, 0.39757641191033699, 0.33069941550246268, 
    0.27117664609268077, 0.21935508208070251, 0.17513377948327211, 
    0.13808420526646181, 0.10756423624070506, 0.082816008813984404, 
    0.06304295880015573, 0.047465630802037695, 0.035358375336397831, 
    0.026070527557531295, 0.019035891433008264, 0.013774009254379212, 
    0.0098860980655303115, 0.0070477949349174989, 0.0050002620516538861, 
    0.0035407213246603517, 0.0025130970770581179, 0.0017992320213657011, 
    0.0013109075333337242, 0.00098285097920191027, 0.00076681957624367741, 
    0.00062679921882881275, 0.00053534029836511206, 0.00047097808297374017, 
    0.00041664580226226014, 0.00035888581248630109, 0.00028763329891732202, 
    0.00019628877378126256, 8.1839337152882585e-05, -5.5173644294252988e-05, 
    -0.00021093802697515825, -0.00037894032694886027, 
    -0.00055078613921411912, -0.00071721407349090464, 
    -0.00086918545960859084, -0.00099896481299784805, -0.0011010402074068104, 
    -0.0011727813011858071, -0.0012147140643407194, -0.0012303505734018393, 
    -0.0012255999764592201, -0.0012078222637342876, -0.0011846758003169959, 
    -0.0011629279891270134, -0.0011474122378268407, -0.0011402950531128038, 
    -0.0011407478471402853, -0.0011450727412478461, -0.001147258708941363, 
    -0.0011398972305660868, -0.0011153354079484908, -0.001066923444721736, 
    -0.00099020764001228677, -0.00088388844762149748, 
    -0.00075041716988572937, -0.00059608532691517743, 
    -0.00043054492997925256, -0.00026576432078077384, 
    -0.00011457148785049725, 1.0994189717051742e-05, 0.00010121622910487564, 
    0.00014987980266169197, 0.00015489607669577651, 0.00011835165461213341, 
    4.6008021593951905e-05, -5.3618307883765893e-05, -0.00017041157475866666, 
    -0.00029387298253892189, -0.00041422319851361448, 
    -0.00052326704063675709, -0.00061493557242091421, 
    -0.00068548687970619289, -0.00073337724939174912, 
    -0.00075889566432045703, -0.00076361741901130457, 
    -0.00074982807167090848, -0.00072000559681680335, 
    -0.00067645252952573361, -0.00062116841980579273, 
    -0.00055592687196103299, -0.00048252782098513817, 
    -0.00040312169258116157, -0.00032048468299175474, 
    -0.00023815836371674545, -0.00016039719481285495, 
    -9.1919101591361895e-05, -3.7494084734936709e-05, 
    -1.4403285622883875e-06, 1.2896772816100193e-05, 3.5915970489071108e-06, 
    -2.9539506681894445e-05, -8.4795971523341665e-05, -0.000158632623067797, 
    -0.0002458787767711558, -0.00034009776097916248, -0.00043404425422304758, 
    -0.0005201631380214283, -0.00059107448935994279, -0.00063999341723882741, 
    -0.00066106658870106877, -0.00064960993716188541, 
    -0.00060226844861130976, -0.00051712977540205036, 
    -0.00039379036243402559, -0.00023340283592583293, 
    -3.8674175478770027e-05, 0.00018619669994786263, 0.00043565006934356886, 
    0.00070297589293555969, 0.00098058626505182996, 0.0012603354458573894, 
    0.0015338772361706771, 0.0017930303826919425, 0.0020301548393651466, 
    0.0022385395398136529, 0.0024127701020697145, 0.0025490856906807201, 
    0.0026457027649737642, 0.0027030537318808905, 0.0027238880159017528, 
    0.0027131634442155712, 0.0026776916585877384, 0.0026255271815292147, 
    0.0025651730700579751, 0.0025047120905538041, 0.0024509911312271364, 
    0.0024089742975157229, 0.0023813828280603048, 0.0023686387776061203, 
    0.00236912260244383, 0.0023796689706339111, 0.0023961975694490514, 
    0.002414384734130783, 0.0024302265365806243, 0.0024404627910266838, 
    0.0024427787975856066, 0.002435812044997428, 0.0024189999658386801, 
    0.0023923142845385, 0.0023559853370855848, 0.00231022692982923, 
    0.0022550380619816941, 0.002190059565030409, 0.0021145009138000648, 
    0.0020271389746378387, 0.0019264056621323717, 0.0018105806277614672, 
    0.0016780686302522352, 0.0015277227019975697, 0.0013591271521722454, 
    0.001172753079139196, 0.00096995395956809432, 0.00075281929728112978, 
    0.00052398045222100723, 0.00028646606843304323, 4.3686531777662501e-05, 
    -0.00020045979170330372, -0.00044142672728683647, 
    -0.00067388678143476971, -0.00089170378130344868, -0.0010880409475564467, 
    -0.0012556144460456802, -0.0013870866142281914, -0.0014755470734789246, 
    -0.0015150450790471089, -0.0015011285475392746, -0.0014313159030767144, 
    -0.0013054665181121419, -0.0011260181419089558, -0.00089802997651380141, 
    -0.00062904779045440482, -0.00032875888378432503, 
    -8.4442590925211591e-06, 0.00031972503173276342, 0.00064352127314285499, 
    0.0009515363040647146, 0.0012340333913999297, 0.0014836612480503685, 
    0.0016959328084309394, 0.001869381364877559, 0.0020053548784859797, 
    0.0021074648662973154, 0.0021807848627738149, 0.0022309101049605064, 
    0.0022630515313289525, 0.0022812823581580001, 0.0022880667599229423, 
    0.0022841106805837146, 0.0022685698319410692, 0.0022395583042108327, 
    0.0021948735893247331, 0.0021328094426928275, 0.0020529130600167398, 
    0.0019565531785346534, 0.0018472163143181208, 0.001730468078285559, 
    0.0016135999136145432, 0.0015050205146944632, 0.0014134541586976175, 
    0.0013470882078050863, 0.0013127499735988513, 0.0013152133706093173, 
    0.0013567207151404591, 0.0014367519275918601, 0.0015520618424473308, 
    0.0016969520994865922, 0.0018637354898103258, 0.0020433174242952454, 
    0.0022258220779455074, 0.0024011887903908394, 0.0025596966719244165, 
    0.0026923963764715914, 0.0027914667742666736, 0.0028505215653320663, 
    0.0028649160340263988, 0.0028320738135825161, 0.0027518213955965531, 
    0.0026267119193093195, 0.0024622433597587187, 0.0022668980538563914, 
    0.002051921067315702, 0.0018308029042492162, 0.0016184409615336878, 
    0.0014300685934837312, 0.0012800411704715318, 0.0011806134963871866, 
    0.0011408717594469789, 0.0011659274394995524, 0.0012564813674954124, 
    0.0014087750922915014, 0.0016149117895165889, 0.0018634805386817828, 
    0.0021403924400361786, 0.0024298106952474136, 0.0027151017572251985, 
    0.002979720274575728, 0.003207992376196068, 0.0033857916765986824, 
    0.0035011105028047019, 0.0035445662193780937, 0.003509839631495397, 
    0.0033940647564659611, 0.0031981106260001737, 0.0029267006649893873, 
    0.002588276454348626, 0.0021945448075571497, 0.0017597107525262003, 
    0.0012994310269398722, 0.00082961535457360455, 0.00036520167169024412, 
    -8.0932817329913782e-05, -0.00049881080969191912, 
    -0.00088184000562703806, -0.0012268723841056457, -0.0015338460441634847, 
    -0.0018050544158355528, -0.0020441894958277878, -0.0022553050053368173, 
    -0.0024418934003678431, -0.0026062227732822079, -0.0027490083117316893, 
    -0.0028694399792946489, -0.0029655100957970376, -0.0030345650324850107, 
    -0.0030739544257766226, -0.0030816714289892857, -0.0030568729163645801, 
    -0.0030002225497915182, -0.0029140051395837897, -0.0028020141881962518, 
    -0.0026692541187669427, -0.0025215045252465484, -0.0023648206241564159, 
    -0.0022050562396829939, -0.0020474647889040577, -0.0018964320899772626, 
    -0.0017553376901023885, -0.0016265583383200466, -0.0015115534660339459, 
    -0.0014109919054062284, -0.0013249041857134579, -0.0012528114099997613, 
    -0.001193858663298023, -0.0011469546468157721, -0.0011109274001732858, 
    -0.0010847035937870978, -0.0010674809798045285, -0.0010588904136186216, 
    -0.0010591035919146514, -0.001068877233721567, -0.0010895215962790671, 
    -0.0011227851593417462, -0.0011706801315571752, -0.001235234312156499, 
    -0.0013181869005926303, -0.0014206538896370563, -0.0015427855467910489, 
    -0.0016834443729476687, -0.0018399654270407873, -0.0020080325326964684, 
    -0.0021816976096228251, -0.0023535726229314013, -0.0025151835112381194, 
    -0.0026574891627087257, -0.0027715020153258013, -0.0028489666146007311, 
    -0.0028829660459920446, -0.0028683719451060522, -0.0028020606240325274, 
    -0.0026828925545496073, -0.0025115079058829937, -0.0022900536615568122, 
    -0.0020219440536808886, -0.0017117151881416654, -0.0013649543637418687, 
    -0.0009882660607293365, -0.00058919671712230517, -0.000176080618286286, 
    0.00024220383334355657, 0.00065651729495838672, 0.0010577875773623156, 
    0.0014373348873563069, 0.001787206096646222, 0.0021005161603617618, 
    0.0023717832140895366, 0.002597210385556669, 0.0027748796834477286, 
    0.0029048015944992483, 0.0029888095714461775, 0.0030302952400289018, 
    0.003033821661112135, 0.0030046581626382183, 0.0029483052593409637, 
    0.0028700793765932564, 0.0027748063233138101, 0.0026666759527343899, 
    0.0025492537955924864, 0.0024256586861598414, 0.002298833327439027, 
    0.0021718400852942452, 0.0020480872563233337, 0.0019314331001853411, 
    0.0018261235943710381, 0.0017365705629512221, 0.0016669676823498453, 
    0.0016207865315258684, 0.0016002162306780539, 0.0016056347773308768, 
    0.0016351960238901097, 0.0016846132344041887, 0.001747214446767797, 
    0.0018142647853151281, 0.0018755787315527484, 0.0019203390630419888, 
    0.0019380325444399566, 0.0019193737006955936, 0.0018570875652987235, 
    0.0017464398266935661, 0.0015854780035421383, 0.0013749569651804188, 
    0.0011180389980731079, 0.0008198162186860478, 0.00048675676660664814, 
    0.00012615357395032634, -0.0002543815825196197, -0.00064732527314134204, 
    -0.0010455149425014439, -0.0014422679291694034, -0.0018313420605755907, 
    -0.0022067662674867821, -0.0025625802583341432, -0.002892571012645596, 
    -0.0031900665481862591, -0.0034478621432837298, -0.003658331454500978, 
    -0.0038137631179871235, -0.0039069038753090377, -0.0039316917097580893, 
    -0.0038840872019255969, -0.0037629016261173385, -0.0035704467597405028, 
    -0.0033128523731434322, -0.0029999449031202171, -0.0026446678257621876, 
    -0.0022621277941539271, -0.0018684074982986049, -0.0014793214923242877, 
    -0.0011092780104647831, -0.00077038728467128999, -0.00047191722613219731, 
    -0.00022011996027803372, -1.8396803167509772e-05, 0.00013230548517763964, 
    0.00023300711384299056, 0.00028624979938205949, 0.00029580721435085508, 
    0.00026656737319485972, 0.00020457759164363738, 0.00011712778378116526, 
    1.276990155220733e-05, -9.883753519543665e-05, -0.00020732295231896597, 
    -0.00030221919334664696, -0.00037375359183227372, 
    -0.00041371853923074381, -0.00041629722803459434, 
    -0.00037871095517539119, -0.00030156683105642145, 
    -0.00018884552025761082, -4.7489063948148987e-05, 0.0001133150108445762, 
    0.00028307580742889049, 0.00045098596848897575, 0.00060686157527928665, 
    0.00074188213169547551, 0.00084910609157116739, 0.00092371835846465598, 
    0.00096300679138563137, 0.00096615031931696202, 0.00093385415467128101, 
    0.00086794200662074867, 0.00077099181556338425, 0.00064609814013603668, 
    0.0004968098787710908, 0.00032725039696651609, 0.00014236457918294311, 
    -5.1816606575037716e-05, -0.00024802676667127604, 
    -0.00043782933748916404, -0.00061195866824304858, 
    -0.00076092204407300591, -0.00087578495677193469, 
    -0.00094903147566980164, -0.00097536733657678618, 
    -0.00095234202257694662, -0.00088069655770533096, 
    -0.00076435456639623533, -0.00061003438756868664, 
    -0.00042649960036914865, -0.00022355491366536829, 
    -1.0955740288354647e-05, 0.00020257208876999511, 0.00041003176332982718, 
    0.00060652047312369554, 0.00078929690744076303, 0.00095758144902133779, 
    0.0011121469883879098, 0.001254738387042092, 0.0013873987608661617, 
    0.0015118130531058848, 0.0016287833301590127, 0.0017379329757162938, 
    0.0018376809592031951, 0.0019254642574455245, 0.0019981563902704657, 
    0.0020525978079383232, 0.002086147015662647, 0.0020971793268404603, 
    0.0020854826187790302, 0.0020524865029774822, 0.0020013100040805185, 
    0.0019365970259824501, 0.001864154164647998, 0.0017904369854660235, 
    0.001721925978956754, 0.001664501154739264, 0.0016228753233217478, 
    0.0016001994996166439, 0.0015978682804342554, 0.0016155810939948573, 
    0.0016516143712238967, 0.0017032515074806194, 0.0017672981171101307, 
    0.0018405434136508202, 0.001920113983166646, 0.0020036374922179738, 
    0.0020891857010630938, 0.0021750465462989726, 0.0022593654189663982, 
    0.0023397855924542433, 0.0024131884690678502, 0.002475627122564997, 
    0.002522469430011845, 0.0025487309399041319, 0.0025494883749306954, 
    0.0025202903717292113, 0.0024574763961476404, 0.0023583614974188455, 
    0.0022212965977017572, 0.0020456421109794148, 0.0018316952385457053, 
    0.001580628858862647, 0.0012944716255515259, 0.00097615937558060285, 
    0.00062962753439710351, 0.00025989374483015965, -0.00012691572337033492, 
    -0.00052362897976363876, -0.00092221856573329423, -0.001314114232860864, 
    -0.0016905847934943535, -0.0020431708328282568, -0.0023640873632783193, 
    -0.0026465760287677858, -0.0028851871082662454, -0.0030759923771623053, 
    -0.0032167497252554335, -0.0033070039161410833, -0.0033481194652539925, 
    -0.0033431985795441001, -0.003296898162330968, -0.0032151159879711851, 
    -0.003104614889047131, -0.0029726176730562374, -0.0028264389509257948, 
    -0.0026731737105158567, -0.0025194433504912243, -0.0023711876000599682, 
    -0.0022334888372646279, -0.0021104271776598727, -0.0020049783373935191, 
    -0.0019189602337839138, -0.0018530485930288486, -0.0018068402505183323, 
    -0.0017790039402417637, -0.0017674941006982916, -0.0017698125723988498, 
    -0.0017832374557217034, -0.0018049991464771896, -0.0018323580081813999, 
    -0.0018625888089753521, -0.0018929165793094807, -0.0019204328192872701, 
    -0.0019420547559076842, -0.001954556334119372, -0.0019547198576766499, 
    -0.0019395792933726069, -0.0019067161882773082, -0.0018545385386926356, 
    -0.0017824908525862716, -0.0016911455560735642, -0.0015822111927192434, 
    -0.0014584699727928072, -0.0013236824019849528, -0.0011824316939504918, 
    -0.0010398589207966608, -0.00090125270505070408, -0.00077147942578520575, 
    -0.00065431264340534375, -0.00055177139509047666, 
    -0.00046358017671188178, -0.00038687055219970419, 
    -0.00031620766788163025, -0.00024397532688182638, 
    -0.00016109127769338376, -5.8008029548261764e-05, 7.4103844349091247e-05, 
    0.00024212133639246082, 0.00044981864681331005, 0.00069696264811358155, 
    0.00097878309919905717, 0.0012859316141823659, 0.0016049941009454493, 
    0.0019195172720465881, 0.0022114841388040777, 0.0024630510360833364, 
    0.0026583412074205255, 0.0027850604912312495, 0.0028356948800924795, 
    0.0028081426733232097, 0.0027056840211402366, 0.0025363372380383005, 
    0.0023116989894322836, 0.0020454936730395271, 0.0017520553451704549, 
    0.0014449627082114543, 0.0011360253236681517, 0.00083472371024192365, 
    0.00054812508388558923, 0.00028122381236943267, 3.7563494462824986e-05, 
    -0.00018000942856260383, -0.0003686766000915393, -0.00052519931998085839, 
    -0.0006458065811884645, -0.00072645400147301786, -0.00076340954788260999, 
    -0.00075404980558283451, -0.00069770611105637718, 
    -0.00059636068332165543, -0.00045505784723750246, 
    -0.00028188073852877934, -8.7510246624975671e-05, 0.00011560594789447904, 
    0.00031435380493503076, 0.0004961360091290636, 0.00064999033230911146, 
    0.00076748339024613305, 0.00084332115048500527, 0.00087561169507561847, 
    0.00086582964897866717, 0.00081850861019611035, 0.00074073201803741512, 
    0.00064147289889253032, 0.00053082439185240572, 0.00041916191712571677, 
    0.00031628823785291474, 0.0002306121543696187, 0.00016843108088888308, 
    0.00013339395953570514, 0.00012623358553687748, 0.00014483320068695441, 
    0.00018463376502238072, 0.00023933294735637852, 0.00030174745308620917, 
    0.00036463677956297618, 0.00042134891928735874, 0.00046619970808272813, 
    0.00049458323511533512, 0.00050292238109638486, 0.00048855528930779333, 
    0.00044969493733546776, 0.0003855120985073613, 0.00029635745244188595, 
    0.00018405188768523122, 5.2133995250526805e-05, -9.408571188799131e-05, 
    -0.00024774246255192923, -0.00040094638698512451, 
    -0.00054553516874190607, -0.0006739403510191579, -0.00077996049307969546, 
    -0.0008593078638345317, -0.00090982641872320181, -0.00093136230840693435, 
    -0.00092534480713680827, -0.00089421954681344297, 
    -0.00084084673579033406, -0.00076797257484161399, -0.0006778885712872988, 
    -0.00057230803921274557, -0.00045247774549957755, 
    -0.00031948032642653551, -0.00017466710752152883, 
    -2.0108628975698254e-05, 0.00014103527246902048, 0.00030431913448764433, 
    0.00046401643381800841, 0.00061338261405683337, 0.000745108638214768, 
    0.00085195625743606461, 0.00092747218727813477, 0.00096668509593412642, 
    0.000966677889015692, 0.00092691884679876706, 0.00084929773259081705, 
    0.00073784346649976456, 0.00059820013534072551, 0.00043695589632943601, 
    0.00026093675962042063, 7.6596365227248574e-05, -0.00011042522334221161, 
    -0.00029552020079470786, -0.00047512260971106741, 
    -0.00064657430818953023, -0.0008079169372925025, -0.00095770007502185507, 
    -0.0010948440280461906, -0.0012185856550372153, -0.0013285151032428001, 
    -0.0014246725270452613, -0.0015076663583058899, -0.0015787296759507538, 
    -0.0016396412556573302, -0.0016924965262391171, -0.0017393278261553522, 
    -0.0017816783667605602, -0.0018202298055643726, -0.0018545500185086548, 
    -0.0018830668652426673, -0.0019032471026980567, -0.0019119789964588225, 
    -0.001906075645686152, -0.0018828204911714376, -0.0018404570698613441, 
    -0.0017785457660809871, -0.0016981226297216692, -0.0016016544210986482, 
    -0.0014927881912984704, -0.0013759799010145373, -0.0012560739025175326, 
    -0.0011379218904414145, -0.0010260877730573, -0.0009246370391833501, 
    -0.00083700234624914784, -0.00076587425451287458, 
    -0.00071309267036943468, -0.00067953626425293519, 
    -0.00066502307126258898, -0.00066827023309040234, 
    -0.00068692770088749902, -0.00071775900968603019, 
    -0.00075692801849524172, -0.00080039869068749051, 
    -0.00084439363871907668, -0.00088581843664974416, 
    -0.00092260879800465899, -0.00095388763186758803, 
    -0.00097991112600228606, -0.0010017710697923282, -0.0010209217032648575, 
    -0.0010386293718092523, -0.0010554683546002079, -0.0010710139888533865, 
    -0.0010838132201937774, -0.0010916460888888879, -0.0010919949328665561, 
    -0.0010825990084340693, -0.001061938010367848, -0.0010295509917733572, 
    -0.00098617428642519414, -0.00093370424825628948, -0.0008750727834371234, 
    -0.00081404444644403917, -0.00075499719700364591, 
    -0.00070267036332851817, -0.00066191130958941123, 
    -0.00063743825823504114, -0.00063362690310728891, 
    -0.00065429763658220337, -0.00070246980098489565, 
    -0.00078006382853618497, -0.00088758196967731568, -0.001023818366721486, 
    -0.0011856762778211297, -0.0013681736907495354, -0.0015646741382368502, 
    -0.001767348043541595, -0.0019677856895622329, -0.0021576835926745454, 
    -0.0023294781881608205, -0.0024768576163989183, -0.0025950934330331342, 
    -0.0026811771547581328, -0.0027338096040330057, -0.0027532561884577268, 
    -0.0027411359796417562, -0.0027001513732856589, -0.0026338061719453697, 
    -0.0025461313816375493, -0.0024414583373991877, -0.002324249064929289, 
    -0.0021990229638707381, -0.0020703251139061792, -0.0019427539909184677, 
    -0.0018209459950526098, -0.0017095020834158843, -0.0016128145088503496, 
    -0.0015347911906503382, -0.0014785253034240839, -0.0014459652242793614, 
    -0.0014376302224428656, -0.0014524577217755223, -0.0014877725058243219, 
    -0.0015394073331554418, -0.0016019476397806627, -0.0016691047360904473, 
    -0.0017341673635373803, -0.0017905394736326193, -0.0018323139923719799, 
    -0.0018548503605888473, -0.0018552921091739328, -0.0018329584114422006, 
    -0.0017895398404882664, -0.0017290254666920825, -0.0016573587320569919, 
    -0.0015818214145517549, -0.0015102340867393074, -0.0014500554701602046, 
    -0.001407522289609631, -0.0013869251862778642, -0.0013901267728644103, 
    -0.0014163766892083941, -0.0014624404988482311, -0.0015230474374882126, 
    -0.0015915650297560733, -0.0016608068713360325, -0.0017238442118094337, 
    -0.0017746907273296277, -0.001808768811596408, -0.0018230884791678244, 
    -0.0018161580622350416, -0.0017876665424484376, -0.0017380335135621248, 
    -0.001667950294970277, -0.0015780207416495062, -0.0014685868212644369, 
    -0.0013397754948345523, -0.0011917428314854154, -0.0010250838545644771, 
    -0.00084128352618756982, -0.00064312543933066964, 
    -0.00043493408023122948, -0.00022257067391305945, 
    -1.3142151618474937e-05, 0.00018554528731061655, 0.00036569695098998239, 
    0.00052028159740829605, 0.00064368690787476232, 0.00073216831063576803, 
    0.00078402617811781981, 0.00079951604591786099, 0.00078054409242383387, 
    0.00073023012767698954, 0.00065244542149558787, 0.00055139286128436658, 
    0.00043129274205622653, 0.00029619766338589092, 0.00014991136483668763, 
    -4.0240863073633209e-06, -0.00016230204029307418, 
    -0.00032183511503402698, -0.00047978250252502473, 
    -0.00063362968804423967, -0.00078132369674735924, 
    -0.00092144635454933805, -0.0010533720110392814, -0.0011773654706980811, 
    -0.0012945757756934408, -0.0014068894707737522, -0.0015166603913708979, 
    -0.0016263263371281659, -0.001737968574974632, -0.001852890672860757, 
    -0.0019712763055079029, -0.0020919977655956927, -0.0022126129268436644, 
    -0.0023295578099110461, -0.0024385273034395172, -0.0025350096788802861, 
    -0.002614864609775953, -0.0026748941562658992, -0.0027132876309443471, 
    -0.0027298669944389956, -0.0027261189438503989, -0.0027049861888737907, 
    -0.0026704924544711638, -0.0026272601272345187, -0.0025799963847330256, 
    -0.0025330309966626005, -0.0024899635593484434, -0.0024534701328591448, 
    -0.0024252790867292091, -0.0024063048541524616, -0.0023968737527256135, 
    -0.0023969841233515113, -0.0024065033590323797, -0.0024252817615394574, 
    -0.0024530783451238093, -0.0024893591038515307, -0.0025329132077251534, 
    -0.002581422761424001, -0.0026310743710250199, -0.0026763432759413209, 
    -0.0027100634861875871, -0.0027238155836111595, -0.0027086094202558321, 
    -0.0026557421964504735, -0.0025577280149810797, -0.0024091016359785384, 
    -0.0022069802574999488, -0.0019513014465989641, -0.0016447517977479743, 
    -0.0012924693824977378, -0.00090160633912324348, -0.00048086913448786521, 
    -4.0073093777064653e-05, 0.00041026921684099969, 0.00085935148230622139, 
    0.0012964754588545263, 0.0017114405769248328, 0.0020949112074154464, 
    0.002438725004765305, 0.0027361301740646826, 0.0029819284066485499, 
    0.0031725306561003145, 0.0033059426177176154, 0.0033816719676266114, 
    0.0034005937998121101, 0.0033647623127364833, 0.003277222803792963, 
    0.0031417948564906157, 0.0029629012801516636, 0.0027454291033231115, 
    0.0024946526756106035, 0.0022162177852579129, 0.0019161205276378677, 
    0.001600665336081429, 0.0012763564787411255, 0.00094971287243366797, 
    0.00062706105267217483, 0.00031433345288759892, 1.689681884745379e-05, 
    -0.00026057158477144711, -0.00051417131811710851, 
    -0.00074084861994235419, -0.00093847708764170255, -0.0011059437869057986, 
    -0.0012432776169909875, -0.0013517910725466872, -0.001434201477774487, 
    -0.0014946510049722072, -0.0015385854098623059, -0.001572448803786565, 
    -0.0016031891677264125, -0.0016376487444091945, -0.0016819024954782733, 
    -0.0017406221018320806, -0.0018165612911286038, -0.0019101860567401479, 
    -0.0020195029775314601, -0.0021400810470883292, -0.0022652881385730292, 
    -0.002386725140931645, -0.0024948901155222494, -0.0025800169647552957, 
    -0.0026330599543868071, -0.0026467130957659813, -0.002616326190596918, 
    -0.0025406101251335411, -0.0024219888483925636, -0.002266530377772458, 
    -0.0020834106048004683, -0.0018839851598036828, -0.0016806158721907832, 
    -0.001485447771015529, -0.0013093345817144103, -0.0011610538958294954, 
    -0.0010468375224800736, -0.00097023186994140136, -0.00093221315919387302, 
    -0.0009315666808868753, -0.00096539079863368002, -0.0010297072605017247, 
    -0.0011200543398684789, -0.0012319645418657449, -0.001361225506326111, 
    -0.0015039377551194775, -0.001656371113334987, -0.0018147278925754796, 
    -0.0019748767623679118, -0.0021321371546559162, -0.0022811547665100118, 
    -0.0024159098605468451, -0.0025298633091331377, -0.0026162447106942953, 
    -0.0026684672278444862, -0.0026806189125974365, -0.0026479913088893851, 
    -0.0025675601166581159, -0.0024383849519810058, -0.0022618478384406129, 
    -0.0020417132237106777, -0.0017839927581125036, -0.0014966272149641423, 
    -0.0011890366949790314, -0.0008716026555872637, -0.00055513624942514364, 
    -0.00025038311191498571, 3.239183758948299e-05, 0.00028371739757167833, 
    0.00049511650335395648, 0.00065922219247295424, 0.00076980146540514018, 
    0.00082177190847813962, 0.00081122892760095036, 0.00073558158016436806, 
    0.0005938057074772378, 0.00038680494192499599, 0.00011783548612828186, 
    -0.00020710719535164208, -0.00057903465421540014, 
    -0.00098593483519844182, -0.0014130296446050437, -0.0018433402839064992, 
    -0.0022585823989880851, -0.0026403190985719088, -0.0029712834304814373, 
    -0.0032367526890013675, -0.0034257680264687994, -0.0035321038736626916, 
    -0.0035548061515045105, -0.0034982286408594674, -0.0033715619312209228, 
    -0.0031878868051902491, -0.0029628783049678734, -0.0027133364899658311, 
    -0.0024557169199819328, -0.0022048106294265814, -0.0019726989211131529, 
    -0.0017680234197188787, -0.0015955819080418045, -0.0014562540688550722, 
    -0.0013472614258120815, -0.0012627718722892629, -0.0011948505637966267, 
    -0.0011346751256891521, -0.0010738564491220386, -0.0010056714155534357, 
    -0.00092601536522166517, -0.00083396349171084897, 
    -0.00073193402790149324, -0.000625450048313113, -0.00052258283676107856, 
    -0.00043317373447965903, -0.00036782485300911088, 
    -0.00033679656556040194, -0.00034883352633131154, 
    -0.00041004915146428513, -0.00052298793809700322, 
    -0.00068600742064646003, -0.00089310550197005184, -0.0011342472271817174, 
    -0.0013961920267107142, -0.0016637382461440911, -0.0019212174657477824, 
    -0.0021540445420361576, -0.0023500904799607274, -0.0025007049593047947, 
    -0.0026012475324504632, -0.0026511086001325566, -0.0026532336400579616, 
    -0.0026133209756162928, -0.0025388475344865361, -0.002438135944479274, 
    -0.0023196349206155331, -0.0021915119925322848, -0.00206153491187716, 
    -0.0019371681172818506, -0.0018257124047617872, -0.0017343659328270524, 
    -0.0016701132239691379, -0.0016394509920377679, -0.0016479506215695144, 
    -0.0016997737360054212, -0.0017971994594544142, -0.0019402280411659123, 
    -0.002126339198972523, -0.0023504304191647256, -0.0026049490554974886, 
    -0.0028802643078531288, -0.0031652317104045639, -0.0034479602989557346, 
    -0.0037166491367564974, -0.0039603847072405569, -0.004169793350763798, 
    -0.0043374178333128142, -0.0044578331114142715, -0.0045275115270096769, 
    -0.0045445630982435701, -0.0045084067103390449, -0.0044194747025826991, 
    -0.0042789968492595518, -0.004088859969168919, -0.003851579370379003, 
    -0.0035703269954549702, -0.0032490492566813307, -0.0028926398568734171, 
    -0.0025071269371688023, -0.0020998344871351726, -0.0016794766309715769, 
    -0.001256104516999472, -0.00084090504503412419, -0.00044577937054359964, 
    -8.2762993378088532e-05, 0.00023674903760735231, 0.00050284687321629142, 
    0.00070800085142015017, 0.00084783932414692119, 0.00092177095168093288, 
    0.00093328284282082302, 0.00088990354904522036, 0.0008027472786883669, 
    0.00068566545497868192, 0.00055410798221751118, 0.00042377748940115883, 
    0.00030924561139673455, 0.00022267837415077308, 0.00017279795839166576, 
    0.00016419778707660036, 0.00019708280252560468, 0.00026743869742050085, 
    0.00036760586506162814, 0.00048717966693609697, 0.00061414977686943839, 
    0.00073615984740194799, 0.00084181798367051236, 0.00092190396380213149, 
    0.00097041278364985977, 0.00098531421657983864, 0.00096894051796513503, 
    0.00092792317912223884, 0.00087262443545670554, 0.00081609186181043933, 
    0.00077258613435386117, 0.00075586987275973508, 0.00077747566711635805, 
    0.00084518027103390914, 0.00096193277664984587, 0.0011253859312662547, 
    0.0013280525031043812, 0.0015580454230332769, 0.0018002974300594828, 
    0.0020380691548058704, 0.0022545659877715543, 0.0024344806834315034, 
    0.0025653083004854704, 0.002638276531134479, 0.0026488338536167751, 
    0.0025966660019935898, 0.0024852945591636393, 0.0023213384443273319, 
    0.0021135826886665393, 0.0018720196524135073, 0.0016070247024351917, 
    0.0013287682868026551, 0.0010469114581194063, 0.00077053202975688466, 
    0.00050819798023098476, 0.0002681286405438665, 5.8306018492005087e-05, 
    -0.00011349468699087229, -0.00023979972465093581, 
    -0.00031364949489361572, -0.00032894654592187465, -0.0002808828865555662, 
    -0.0001664367286704588, 1.5162671000925213e-05, 0.00026204446863293672, 
    0.00056949228331988004, 0.00092998175866115123, 0.001333461227957636, 
    0.0017678791719562459, 0.0022198261274755157, 0.0026752135233100299, 
    0.0031198592846618058, 0.0035399024535631846, 0.0039220246122225961, 
    0.0042535356208648172, 0.0045224080722965718, 0.0047173852255922161, 
    0.0048282332767017912, 0.0048461793341394999, 0.0047645039287886283, 
    0.0045792025576076624, 0.0042896161626809872, 0.0038988976478486993, 
    0.0034142457180873944, 0.0028468073638668471, 0.0022112584759843503, 
    0.0015250164970981371, 0.00080717353314947553, 7.7235743586748966e-05, 
    -0.00064617135120543753, -0.0013464720034739876, -0.0020100272575277211, 
    -0.0026266628606528546, -0.00318979144285279, -0.0036961925344251921, 
    -0.0041454945241531952, -0.0045395133828607754, -0.0048815056289636585, 
    -0.005175449759388647, -0.0054254487230386726, -0.0056352788141659322, 
    -0.0058081121758949339, -0.0059464302353395984, -0.0060520920445869724, 
    -0.0061264980927059074, -0.0061708170516749927, -0.0061861915403438996, 
    -0.0061738975648906588, -0.0061354310783223454, -0.0060725218421710586, 
    -0.0059871054753741267, -0.0058812677079091678, -0.0057571789548840685, 
    -0.0056171043813524578, -0.0054634464408885013, -0.0052988719099181332, 
    -0.0051264435879188964, -0.0049497081453378049, -0.004772704022284047, 
    -0.0045998340471119208, -0.0044356213815073828, -0.00428436171792357, 
    -0.0041497209717014857, -0.0040343371314979747, -0.0039394772841362955, 
    -0.0038648315687468899, -0.0038084467445409259, -0.0037668547175404043, 
    -0.0037353489454262285, -0.003708393939166733, -0.0036801362344921307, 
    -0.0036449666606620766, -0.0035980425169755792, -0.0035357661778204199, 
    -0.0034561198844739994, -0.0033588199434961014, -0.0032452771310619265, 
    -0.0031183374257486031, -0.0029818671212612454, -0.0028402063935006302, 
    -0.0026976028282149887, -0.0025576934864455585, -0.0024231062525577928, 
    -0.002295242564174892, -0.0021742759049071395, -0.0020593211498703304, 
    -0.001948768776914696, -0.0018406960461827314, -0.0017333161706696895, 
    -0.0016253686113260701, -0.0015164264846201569, -0.0014070183320285879, 
    -0.0012985455217416376, -0.0011929156577586309, -0.0010919516587760743, 
    -0.00099664377110172779, -0.00090637748352133136, 
    -0.00081834116465096484, -0.00072725533015488434, 
    -0.00062555576684228148, -0.00050405783414238573, 
    -0.00035303798751639125, -0.00016356305031654889, 7.1102526254957564e-05, 
    0.00035424793575077886, 0.00068479303386324028, 0.0010568584573009405, 
    0.0014599018462276836, 0.001879420415492877, 0.0022981471283163267, 
    0.0026975769222960869, 0.003059676280653117, 0.0033685610889542705, 
    0.0036119401786199163, 0.0037821843851362658, 0.0038768739640662503, 
    0.0038987682757744405, 0.0038552094572601326, 0.0037570855650724791, 
    0.0036175070650539894, 0.0034504129868049077, 0.0032692756067310516, 
    0.0030860229534183914, 0.0029102656894023403, 0.0027488527285711452, 
    0.0026058015444737188, 0.0024825445102833778, 0.0023784406784860732, 
    0.0022914425085978482, 0.0022187728815204629, 0.00215755231873393, 
    0.0021053245949315797, 0.0020604588888731086, 0.0020224429505154213, 
    0.0019920591638095935, 0.0019714049414231885, 0.0019637335517126995, 
    0.0019730717082994858, 0.002003645209105601, 0.0020591560918545521, 
    0.0021419952740631188, 0.0022525051872942146, 0.0023884413968385601, 
    0.0025446708876022783, 0.0027132206383901404, 0.0028836925603616418, 
    0.0030440449648549287, 0.0031816533819621498, 0.0032845608007245489, 
    0.0033427557739196517, 0.00334929007373907, 0.003301098922760308, 
    0.0031993958040955461, 0.0030495991028118125, 0.0028608317505366869, 
    0.0026450642211081564, 0.0024159940569175825, 0.0021878351503284081, 
    0.0019741421109066271, 0.0017868319659961308, 0.0016354292859544579, 
    0.0015266276723478786, 0.0014640956104299172, 0.0014485492747107597, 
    0.0014780104137639225, 0.0015482537894508013, 0.0016533608386523791, 
    0.001786279289365932, 0.001939348390108394, 0.0021046887574021236, 
    0.0022744429555227575, 0.0024408482795521495, 0.0025961741670214576, 
    0.0027325780018550667, 0.0028419772412852625, 0.0029160414882900289, 
    0.0029463982010802009, 0.0029251061954177317, 0.0028452969203531116, 
    0.0027019538888191259, 0.002492629993380509, 0.0022180041525640495, 
    0.0018821862529142292, 0.0014926812671251048, 0.0010600401172571408, 
    0.00059721875982250044, 0.00011869542661439039, -0.00036053048583334292, 
    -0.00082595833894497019, -0.0012645195646089104, -0.0016653173755992756, 
    -0.0020200366893253644, -0.0023230087960395881, -0.0025708934481964616, 
    -0.0027620666297347067, -0.0028958131357613116, -0.0029715357565332215, 
    -0.0029881399264750424, -0.0029437447704622143, -0.0028357402353841243, 
    -0.0026612029124456153, -0.0024175519885343494, -0.0021033272805698559, 
    -0.0017189469638555371, -0.0012673317495131176, -0.00075430292065263008, 
    -0.00018873544356228119, 0.00041752833613510073, 0.0010499995831251148, 
    0.0016920156230646403, 0.0023253778279226692, 0.002931135894167756, 
    0.0034905161811673718, 0.0039859575048176591, 0.0044022125249767556, 
    0.0047274509921435325, 0.0049542084673870734, 0.0050800760863041828, 
    0.0051080229076969847, 0.005046287732359829, 0.0049078123979445689, 
    0.0047092637812716385, 0.0044697036252610567, 0.0042090185793714615, 
    0.003946277621319415, 0.0036981582395566879, 0.0034776795333548486, 
    0.0032933153488187566, 0.0031486269169820505, 0.0030423196076879615, 
    0.0029688269231559353, 0.0029192168965957587, 0.0028824323350390775, 
    0.002846666747352762, 0.0028007161770269577, 0.0027351506888619714, 
    0.0026431600367940772, 0.0025210256479452982, 0.0023681910961381586, 
    0.0021869951198616711, 0.0019821778463382849, 0.0017602602037206428, 
    0.0015288884833021671, 0.0012962366223723445, 0.0010704947686552399, 
    0.00085948018579014361, 0.00067035869825278038, 0.0005094908059640271, 
    0.00038236073680391458, 0.00029355958256130241, 0.00024673799106344368, 
    0.00024446716963386718, 0.00028798707106965143, 0.00037683193086290135, 
    0.00050842947656074965, 0.00067771240594229347, 0.00087694885722697723, 
    0.0010958537419093564, 0.0013221153283452637, 0.0015422648027413912, 
    0.001742855908849439, 0.001911787657253011, 0.0020395443616811181, 
    0.0021201665000035097, 0.002151804635840855, 0.002136666439462879, 
    0.0020804149828237703, 0.0019910488669091821, 0.0018774451478345041, 
    0.0017478077184841006, 0.0016082930173008448, 0.0014620402700043326, 
    0.0013088321263690021, 0.0011454380959624716, 0.00096663525501350248, 
    0.0007666753400796917, 0.00054094376522966425, 0.00028746751521662491, 
    7.9942270165613671e-06, -0.00029152777654268235, -0.00060112525250706982, 
    -0.00090757626070709881, -0.0011956428998968324, -0.0014495815520508351, 
    -0.0016547259083228045, -0.0017989431447731335, -0.0018737959984744257, 
    -0.0018752897532852617, -0.0018041409456731894, -0.0016655521931225419, 
    -0.0014685683412045574, -0.0012250870912026899, -0.0009486484997000981, 
    -0.00065316863229740224, -0.00035175189430251645, 
    -5.5699135976412926e-05, 0.00022613260825020157, 0.00048760041343142428, 
    0.00072515046077385357, 0.00093738696718127367, 0.0011244780232126852, 
    0.0012875326020552044, 0.001428119094064818, 0.0015479745778491324, 
    0.0016488919202474459, 0.0017326077690915887, 0.001800632005507717, 
    0.0018539011002481076, 0.0018924190717806494, 0.001915011645559976, 
    0.0019194398102741913, 0.0019029936783463526, 0.001863459864938482, 
    0.0018001321860615601, 0.0017144516593786605, 0.001609901275976563, 
    0.0014911662387582494, 0.0013628341006265852, 0.00122813778330169, 
    0.0010881433281698177, 0.00094160168290909041, 0.00078547328532308479, 
    0.00061593573143984637, 0.00042974311231694108, 0.00022564347386948402, 
    5.6252609870323882e-06, -0.00022425331232759569, -0.0004536628922893305, 
    -0.00066847371970469118, -0.0008519139505018499, -0.00098620706078376649, 
    -0.001054404010409062, -0.0010422227077499691, -0.00093969147846453816, 
    -0.00074246234883555457, -0.00045267851055330881, 
    -7.9269754172878678e-05, 0.00036240112315253899, 0.00085161404607837982, 
    0.0013639886927652241, 0.0018736055302118091, 0.00235524074737834, 
    0.0027864062330881026, 0.0031488893268777395, 0.0034297039829121185, 
    0.0036214011517105306, 0.003721829487303333, 0.0037334989159031095, 
    0.0036627236840782651, 0.0035186529616327493, 0.003312305591215287, 
    0.003055651440325016, 0.0027607166474228964, 0.0024387809248609463, 
    0.0020996798889567031, 0.0017513229180524234, 0.001399503028233615, 
    0.0010479868336805925, 0.00069888806134182978, 0.00035326878155137636, 
    1.1863282641327767e-05, -0.00032418608048025545, -0.00065268087999852055, 
    -0.00096994920249097983, -0.0012706914965915229, -0.0015482103114133879, 
    -0.0017950232132858566, -0.0020038772831816715, -0.0021690403642313019, 
    -0.0022876394241832733, -0.0023607852601268201, -0.0023941971578761508, 
    -0.0023981716473036713, -0.0023868335775651117, -0.0023767386382956401, 
    -0.0023850269504714591, -0.0024273268322255884, -0.0025157249221488772, 
    -0.002657037875863764, -0.0028515982806478725, -0.0030927829409607213, 
    -0.0033673121533833294, -0.0036563540063391277, -0.0039373033085365588, 
    -0.0041860691594860821, -0.0043795406264320932, -0.0044979148278015907, 
    -0.0045266275336853434, -0.0044575652473447776, -0.0042894840184051165, 
    -0.0040276719362812045, -0.0036829484356017731, -0.0032702085049452342, 
    -0.0028067128393021168, -0.0023102906832784568, -0.0017977367310332308, 
    -0.0012835967071152512, -0.00077961954365120994, -0.0002949427106146559, 
    0.0001631043853362305, 0.0005878605197598511, 0.00097242687920768569, 
    0.0013092502526721077, 0.001590428142775031, 0.0018085572849743459, 
    0.0019578430215204498, 0.002035232250619978, 0.0020413629574124125, 
    0.0019812837463625047, 0.0018647993423326437, 0.0017063050356895312, 
    0.0015239656351388406, 0.0013382638000775202, 0.0011700286265252458, 
    0.0010381711006196403, 0.0009575567381748584, 0.00093724689479208177, 
    0.00097943848353027703, 0.0010792117246491608, 0.0012251242098312251, 
    0.0014005596923516177, 0.0015856849844128847, 0.001759750986801805, 
    0.0019034606356752167, 0.0020011309151835121, 0.0020423862111903458, 
    0.0020231459112549587, 0.0019458575751805129, 0.0018188867312709585, 
    0.0016551790322223373, 0.00147032424483312, 0.001280317899569183, 
    0.001099370029269581, 0.00093800413864651645, 0.00080173961135960909, 
    0.00069050712076072838, 0.00059882363923238562, 0.00051665225295058727, 
    0.0004307919362491073, 0.00032660363175182567, 0.00018987349342414612, 
    8.5537990583220012e-06, -0.00022575095089775622, -0.00051682640084139975, 
    -0.00086346568835208605, -0.0012597478002544136, -0.0016958998139547758, 
    -0.0021595325273267257, -0.0026370561379558135, -0.0031150114483764848, 
    -0.003581101577040979, -0.0040247739882697427, -0.0044373272735192338, 
    -0.0048115283507767373, -0.0051409436853198385, -0.0054192283126088901, 
    -0.0056395918114511721, -0.0057946025670791729, -0.0058764704088112756, 
    -0.0058778162966613692, -0.0057927334355720008, -0.0056180737455507708, 
    -0.0053546843355143986, -0.0050083276408038578, -0.004590171717994293, 
    -0.0041167075937306756, -0.0036090227120832755, -0.0030915330866609901, 
    -0.0025902623173629548, -0.0021308114997221693, -0.0017362431804244683, 
    -0.0014251156111003789, -0.0012098290319147061, -0.0010955290727941666, 
    -0.0010796934232611074, -0.0011525411484241846, -0.001298224622007954, 
    -0.0014967518754850568, -0.0017262165693529901, -0.0019650648449164618, 
    -0.0021941074170990335, -0.0023980425232632049, -0.0025665110587665295, 
    -0.0026947131423902455, -0.0027835308429441713, -0.0028392052867457322, 
    -0.0028724788861389629, -0.0028972057423451085, -0.0029285647952194929, 
    -0.0029810883627039123, -0.0030667794680432972, -0.0031935358192367322, 
    -0.0033640684042783174, -0.0035753829360748624, -0.0038189013342504094, 
    -0.0040812067167800663, -0.0043453920710513913, -0.0045929506919943517, 
    -0.0048059731195535162, -0.0049694684271076916, -0.0050733908438926429, 
    -0.0051140825909007735, -0.0050948221986884326, -0.0050253745139033018, 
    -0.0049205386752390352, -0.004798147483368596, -0.004676718495186292, 
    -0.0045733266331345335, -0.0045019240693068754, -0.0044722347508925012, 
    -0.004489271227347635, -0.0045534096735225672, -0.0046609815539991857, 
    -0.004805188243145274, -0.0049772243815141264, -0.00516746695970238, 
    -0.0053664704492215783, -0.005565666393910121, -0.0057577009056733143, 
    -0.005936431391679947, -0.0060967267740992233, -0.0062341784972419611, 
    -0.0063448965112405178, -0.0064253683513741996, -0.0064723877273980459, 
    -0.0064831010362404696, -0.0064551135753208389, -0.0063866970343919452, 
    -0.0062770568900009632, -0.0061266403373749076, -0.0059373537814712777, 
    -0.0057127089027785233, -0.0054578959680339802, -0.0051797862906182834, 
    -0.0048869955542943074, -0.0045899315781857521, -0.0043007626744481125, 
    -0.0040331666497195945, -0.0038017565247024519, -0.0036211580286261073, 
    -0.0035047583775491237, -0.0034633335057040809, -0.0035036693824346998, 
    -0.0036274492264282334, -0.0038305909709699455, -0.0041031803456631263, 
    -0.0044301407228099056, -0.004792550867911651, -0.005169467873442103, 
    -0.0055400927069116255, -0.0058859148772923984, -0.0061925707130643113, 
    -0.0064510530915839921, -0.0066581225509262446, -0.0068159598049713273, 
    -0.0069311554661642934, -0.0070134175033169637, -0.0070741441164198738, 
    -0.0071251143194046183, -0.0071773692441809379, -0.0072402321702740779, 
    -0.0073205753496617537, -0.0074221903438184567, -0.0075454241491596805, 
    -0.0076870295632438706, -0.0078403381801693799, -0.0079957680450120465, 
    -0.008141573334319455, -0.0082648607681850058, -0.0083527094552667148, 
    -0.008393310576673977, -0.0083770628480952184, -0.0082974489233579272, 
    -0.0081516337150107886, -0.0079406252284499514, -0.007669028675980123, 
    -0.0073443527243776128, -0.0069760418980921203, -0.0065743138109524597, 
    -0.006149078366906942, -0.0057090811147413861, -0.005261330148653264, 
    -0.0048109325982342646, -0.0043612484603396144, -0.0039143077274316302, 
    -0.003471335786595219, -0.0030332016482299429, -0.0026005874153584622, 
    -0.0021739780639281957, -0.0017533798299047098, -0.0013380271360061557, 
    -0.00092624595917011423, -0.00051551109602791323, 
    -0.00010276163378284161, 0.00031516534807292005, 0.00074126001092588367, 
    0.0011781669584290701, 0.0016283132664245399, 0.0020940948515967128, 
    0.0025780332404503523, 0.0030828406048330182, 0.0036112215050088502, 
    0.0041656024907916582, 0.0047476202564353757, 0.0053575521436373596, 
    0.0059937145313595126, 0.0066520084220970154, 0.0073256256898224723, 
    0.0080051611058394138, 0.0086789981621671116, 0.0093339979715189002, 
    0.0099561922274658335, 0.010531539332226848, 0.011046486149621568, 
    0.011488379145168879, 0.011845775624135956, 0.01210863056999345, 
    0.012268464865184629, 0.012318564386307691, 0.012254183816331855, 
    0.012072816255279126, 0.011774410806385463, 0.011361580634503158, 
    0.010839706038357233, 0.010216834125361828, 0.0095034803188825401, 
    0.0087121257500413166, 0.0078566407483431962, 0.0069516602086766464, 
    0.0060120685360403334, 0.0050526697744478193, 0.0040881735949994539, 
    0.0031332908909801199, 0.0022029594132246233, 0.0013124810811237593, 
    0.00047743249211343607, -0.00028676670762632362, -0.0009655534407309479, 
    -0.0015461859850891904, -0.0020187708043591722, -0.0023772213819931061, 
    -0.0026198736220792089, -0.0027496718813207911, -0.0027738197501459192, 
    -0.0027029964924568536, -0.0025502786927979458, -0.0023300860438870744, 
    -0.0020573413579686737, -0.0017469559066723146, -0.0014136542840030835, 
    -0.001071926266516217, -0.00073605082663113412, -0.00041988796163538284, 
    -0.00013644989221062162, 0.00010283676603495559, 0.00028903240799305557, 
    0.00041663673025202553, 0.0004843878286567086, 0.00049567643336243493, 
    0.0004583991061557776, 0.0003842619076948114, 0.00028741271206175604, 
    0.00018271087526503413, 8.3890425001738851e-05, 2.0880188703079484e-06, 
    -5.511753436517164e-05, -8.3910480949839851e-05, -8.3859743837228545e-05, 
    -5.7269056699846834e-05, -8.2457686557140109e-06, 5.8149637048853199e-05, 
    0.00013681915443337689, 0.00022353538183143455, 0.00031576198178554779, 
    0.00041335348365007164, 0.0005188973282709775, 0.00063747963141072247, 
    0.00077585200618784163, 0.00094081005743984762, 0.0011373672238607514, 
    0.001366825019648992, 0.0016255138548277716, 0.001904426153050597, 
    0.0021898486293183165, 0.0024647001813995514, 0.0027101580773057944, 
    0.0029070383771787342, 0.0030367413614233343, 0.0030821952297008081, 
    0.0030288725602308987, 0.0028663026465185625, 0.0025893956143419675, 
    0.002198935367606313, 0.0017010079273378131, 0.0011056833572587182, 
    0.00042549635577870341, -0.00032580482816246147, -0.0011339753220704657, 
    -0.0019844382098134195, -0.0028620721694747769, -0.0037509458300279434, 
    -0.004634123514869414, -0.0054939484550986439, -0.0063126192594344073, 
    -0.0070730300967208068, -0.0077598625242176486, -0.0083607424072572566, 
    -0.0088674128369068943, -0.0092766278860967766, -0.0095905171140182703, 
    -0.0098163905245707023, -0.0099657639721404973, -0.010052922847711046, 
    -0.010092987258613906, -0.010099998216328595, -0.010085000779424492, 
    -0.010054627113914291, -0.010010219622814211, -0.0099475275602767428, 
    -0.0098569706995593094, -0.0097242279118745865, -0.0095310368116886847, 
    -0.0092563277466052932, -0.0088777356084251483, -0.0083737475729649732, 
    -0.0077262138533905683, -0.0069230863256794948, -0.005960733484108199, 
    -0.0048455091127267459, -0.0035940208847403451, -0.0022323929562149984, 
    -0.00079458626508717824, 0.00067951471988627352, 0.0021461459943834349, 
    0.0035595309440827139, 0.0048738033085062487, 0.0060451065913419604, 
    0.007034335539189719, 0.0078096656778460219, 0.0083490934249095504, 
    0.008642242675328508, 0.0086912753034850236, 0.0085105799774112447, 
    0.0081254970803233302, 0.0075701634592654022, 0.006884713092980544, 
    0.0061124959388196695, 0.0052974895646460372, 0.0044820347408003284, 
    0.0037052150941376517, 0.003001694527879645, 0.0024010412865355301, 
    0.0019273723216331928, 0.0015992107840683189, 0.0014291843830043709, 
    0.0014234558370164853, 0.0015810972658122486, 0.0018934202587439081, 
    0.0023439506345654636, 0.0029093202386792139, 0.0035609240861660604, 
    0.0042669479883915302, 0.0049944143167092179, 0.0057108626741323382, 
    0.0063857307390045234, 0.0069915897470349438, 0.0075051220285039903, 
    0.0079079215266969274, 0.0081867618273817038, 0.0083336037184385953, 
    0.0083453880586147732, 0.0082240494299196925, 0.0079769358628369678, 
    0.0076172289192901936, 0.0071644093247452282, 0.0066436356142378092, 
    0.0060839680212814015, 0.0055150224290313604, 0.0049624337243099224, 
    0.0044432381512656662, 0.0039620375118499069, 0.0035093199067687676, 
    0.0030627717018581165, 0.0025914711299907223, 0.0020620164907027114, 
    0.0014450728399666218, 0.00072077612462010234, -0.00011802627239483546, 
    -0.001064253904299733, -0.002096103645567973, -0.0031769457617412539, 
    -0.0042552441050800419, -0.005266060993246187, -0.0061348828193914778, 
    -0.0067839153917333304, -0.0071401982878658756, -0.0071435648507650242, 
    -0.0067532592239324873, -0.0059520078094644231, -0.004746937151964949, 
    -0.0031680214500347729, -0.0012648915706169488, 0.00089750894910191814, 
    0.0032432621755163859, 0.0056897214146715913, 0.0081512998095517649, 
    0.010542424889268908, 0.012780360916618331, 0.014787003147940018, 
    0.016491242479307801, 0.017831084761367688, 0.01875641943398168, 
    0.019232137533256626, 0.019240926371805054, 0.018785074506611394, 
    0.017886446827475228, 0.016583693432962041, 0.014927820322572357, 
    0.01297614117186225, 0.010786857468893938, 0.0084149794241831812, 
    0.0059105100168745147, 0.0033195198144983446, 0.00068634991570464237, 
    -0.0019434105852175537, -0.0045203505221381021, -0.0069902140633877393, 
    -0.0092954842316866817, -0.011378587715175355, -0.013186582998878836, 
    -0.01467650667439257, -0.015818965395795036, -0.016600080533322313, 
    -0.017021994593606132, -0.017103308739416907, -0.016880716803436113, 
    -0.016409747272349121, -0.015764388352184393, -0.015031792196088651, 
    -0.01430265712417848, -0.013657934913500388, -0.013156406857009645, 
    -0.012824476040772397, -0.012650863886178247, -0.012588574881623408, 
    -0.012563025318288359, -0.012485041795052025, -0.012264119613451686, 
    -0.011824247862123587, -0.01111458469270581, -0.010119776030136137, 
    -0.0088647847800283341, -0.0074157639484152948, -0.005874311062562987 ;

 Fqt-F =
  // Fqt-F(0, 0-1999)
    1, 0.99983779032138842, 0.99935247732892418, 0.9985480218385705, 
    0.997430947728428, 0.99601018783675077, 0.99429688146883977, 
    0.99230413397229322, 0.9900467495476748, 0.98754094859609165, 
    0.98480407964832251, 0.98185433493938024, 0.97871047752977869, 
    0.97539158348587351, 0.97191680439144645, 0.96830515118414395, 
    0.96457529937292252, 0.96074541758105614, 0.95683301794480302, 
    0.95285482613698624, 0.94882667437897195, 0.94476341408091102, 
    0.94067884979982797, 0.93658569407068759, 0.93249554220725994, 
    0.92841886512124816, 0.9243650172562331, 0.92034225575552131, 
    0.91635776528173452, 0.91241769488799684, 0.90852720164097178, 
    0.90469050120663141, 0.90091092589560151, 0.89719098413235598, 
    0.89353242294473245, 0.88993629112277606, 0.88640299976156289, 
    0.88293238424825105, 0.87952376429337509, 0.87617600343083168, 
    0.87288756757657415, 0.86965658637709919, 0.86648091100087388, 
    0.86335817395812076, 0.86028584507904582, 0.85726128553155678, 
    0.85428179564730078, 0.85134465917491176, 0.8484471805472984, 
    0.84558671710663458, 0.84276070898884448, 0.83996670130449869, 
    0.83720236486089783, 0.83446551343227549, 0.83175411495804019, 
    0.82906630249668312, 0.82640037917047293, 0.82375482145415568, 
    0.82112828055394338, 0.81851957871038306, 0.81592770693166916, 
    0.81335181640251608, 0.81079120910249336, 0.80824532765770285, 
    0.80571373835494831, 0.8031961201173331, 0.80069224839203135, 
    0.79820198083701366, 0.79572524111587561, 0.7932620040392776, 
    0.79081228139346182, 0.78837610868096963, 0.78595353383396982, 
    0.78354460595833941, 0.78114936732307927, 0.77876784645286479, 
    0.77640004966208187, 0.7740459582816992, 0.7717055198706293, 
    0.76937864627656105, 0.76706520828280089, 0.76476503241563254, 
    0.76247790064084253, 0.76020354886732322, 0.75794166710738975, 
    0.75569190487449034, 0.75345387607901182, 0.75122716924840249, 
    0.74901135562564014, 0.74680600401445807, 0.74461069140599567, 
    0.74242501406944961, 0.74024859874185611, 0.73808110736064947, 
    0.73592224600960787, 0.73377176872189176, 0.73162948373105896, 
    0.72949525772776025, 0.72736901840332169, 0.72525075609696521, 
    0.72314052158316455, 0.72103842579126021, 0.71894463397974273, 
    0.71685936383628734, 0.71478288091687403, 0.71271549299280357, 
    0.71065754596564934, 0.70860941615055073, 0.7065715082901487, 
    0.70454424972893248, 0.70252808664216138, 0.70052347737813903, 
    0.69853088890210646, 0.69655078853239738, 0.69458364070715872, 
    0.69262989898359117, 0.69069000143239812, 0.68876436356172011, 
    0.68685337563044269, 0.68495739392668098, 0.68307673967635252, 
    0.68121169407130078, 0.67936249672296667, 0.67752934346752047, 
    0.6757123816960966, 0.67391170817106727, 0.67212736430599662, 
    0.67035933349658294, 0.66860754064385752, 0.66687185195687049, 
    0.66515207541965848, 0.66344796413612672, 0.66175921850245434, 
    0.66008549102947822, 0.65842638748126392, 0.65678147281129207, 
    0.65515027613617483, 0.65353229538040924, 0.65192700356442834, 
    0.65033385534860633, 0.64875229283372626, 0.64718175126063215, 
    0.64562166631490892, 0.64407147895454797, 0.6425306402223423, 
    0.64099861589026796, 0.63947489148548053, 0.63795897568289384, 
    0.63645040114081308, 0.63494872851571105, 0.63345354711060275, 
    0.63196447537255018, 0.63048116402263732, 0.62900329265952237, 
    0.62753057167304971, 0.62606274110557336, 0.62459957023032564, 
    0.62314085284221843, 0.62168640725237012, 0.62023607098436451, 
    0.61878970318283777, 0.61734717650823745, 0.61590837867692216, 
    0.61447320967879726, 0.61304158098906625, 0.6116134127254248, 
    0.61018863344150864, 0.60876717872468511, 0.60734899276196308, 
    0.60593402939394192, 0.60452225654971325, 0.60311365709606857, 
    0.60170822759412979, 0.60030597452851087, 0.59890690982495187, 
    0.59751104485527895, 0.59611838561604513, 0.5947289272103381, 
    0.59334265381208184, 0.59195953557663761, 0.59057952946854297, 
    0.58920257968017409, 0.58782861912436724, 0.58645757102304108, 
    0.58508935255510564, 0.58372387923806124, 0.58236106481838823, 
    0.58100082617748627, 0.5796430860886268, 0.57828777438644396, 
    0.57693483083127528, 0.5755842051401675, 0.57423585786078446, 
    0.57288975976107726, 0.57154589362194996, 0.57020425275651776, 
    0.56886484319507236, 0.56752768278279186, 0.56619280363117397, 
    0.56486025263370598, 0.56353009165090306, 0.56220239784639492, 
    0.56087726264433424, 0.55955478847381168, 0.55823508679035772, 
    0.5569182743707124, 0.55560447165200522, 0.55429379803982304, 
    0.55298637483310076, 0.55168232062766687, 0.55038175565378944, 
    0.54908480204653176, 0.54779158272420458, 0.54650222402600235, 
    0.5452168544024073, 0.54393560680102182, 0.54265861695418594, 
    0.54138602615295028, 0.54011798220010632, 0.538854641016555, 
    0.53759616742280003, 0.53634273583259851, 0.53509453167487941, 
    0.53385174793343804, 0.53261458696017383, 0.53138325410960618, 
    0.53015795551424993, 0.52893889160582253, 0.52772625033271725, 
    0.52652020188910575, 0.52532088887951012, 0.52412841802287591, 
    0.5229428515727893, 0.52176419913734073, 0.52059241182030225, 
    0.51942737858044108, 0.51826893057282963, 0.51711684166760619, 
    0.51597084247394487, 0.51483062529257007, 0.51369585687988739, 
    0.51256618720227631, 0.51144125613428826, 0.51032070015536801, 
    0.50920415717552658, 0.50809127119170006, 0.50698169166490836, 
    0.50587507852201741, 0.50477109955212773, 0.50366942967374295, 
    0.50256975005854954, 0.50147174848488452, 0.50037511980543126, 
    0.49927956665369849, 0.49818480396620474, 0.49709056275830377, 
    0.49599659402013757, 0.49490267535609833, 0.49380861501908646, 
    0.49271425558204307, 0.49161947597694278, 0.49052419249766049, 
    0.48942835636821752, 0.48833195357023451, 0.48723500200610587, 
    0.48613755110433499, 0.4850396776495251, 0.48394148358219286, 
    0.48284309715697721, 0.4817446674520125, 0.48064636198024807, 
    0.47954836079204816, 0.47845085052037212, 0.47735401855201953, 
    0.47625804527897136, 0.47516309691766184, 0.47406932033973997, 
    0.47297684132949552, 0.47188576081437805, 0.47079615516442935, 
    0.46970807677125831, 0.46862155425991714, 0.46753659402127118, 
    0.4664531787580608, 0.46537126923714284, 0.46429080178287246, 
    0.46321168764506909, 0.46213381777546209, 0.46105706575547367, 
    0.45998129857045789, 0.45890638333260847, 0.4578321963046923, 
    0.45675862912014209, 0.45568559899677058, 0.45461304768212113, 
    0.45354094610437989, 0.45246929337668607, 0.45139811683997205, 
    0.45032747174952681, 0.44925744168431281, 0.44818813747371211, 
    0.44711969497602116, 0.44605227782791934, 0.44498607214049601, 
    0.44392128570157358, 0.44285814625396419, 0.4417968982492953, 
    0.44073779831179527, 0.43968110782106457, 0.43862708725642879, 
    0.43757598867151792, 0.43652804904605341, 0.43548348593908254, 
    0.43444249540051072, 0.43340525167377647, 0.4323719079582381, 
    0.43134259921350188, 0.43031744601632604, 0.42929655715666476, 
    0.42828003362803518, 0.42726797308439612, 0.42626047331183448, 
    0.42525763368716313, 0.42425955672127019, 0.42326634854017664, 
    0.42227811507860885, 0.42129495887149138, 0.42031697814994307, 
    0.41934426232391669, 0.41837689137940531, 0.41741493639917077, 
    0.41645845543618232, 0.41550749308783291, 0.41456207937456069, 
    0.41362222849695529, 0.41268793638299861, 0.41175918023075686, 
    0.41083591425648924, 0.40991806768094124, 0.40900554188979499, 
    0.40809820809481878, 0.40719590447873927, 0.4062984374179609, 
    0.40540558651969266, 0.40451710862389506, 0.4036327464962568, 
    0.40275223491221385, 0.40187531255551201, 0.40100172676686252, 
    0.40013124316176119, 0.39926365096483279, 0.39839877279457175, 
    0.3975364699756459, 0.39667664330669106, 0.39581923456977719, 
    0.39496422062793346, 0.39411160628605707, 0.39326141761038708, 
    0.39241369640841939, 0.39156849522953574, 0.39072587552586452, 
    0.38988590392362371, 0.3890486501045709, 0.38821418293740079, 
    0.38738256961792722, 0.38655387173805117, 0.38572814948695344, 
    0.38490545700147771, 0.38408584832834791, 0.38326937359775493, 
    0.38245608267529957, 0.38164602451922708, 0.38083924787363127, 
    0.38003580037482854, 0.3792357315570124, 0.37843908870287946, 
    0.37764591655796192, 0.37685625443343423, 0.37607013309186649, 
    0.37528757414504599, 0.3745085858674041, 0.37373316375947496, 
    0.37296129094158204, 0.37219293573620355, 0.37142804631154108, 
    0.37066654651758024, 0.36990832716051791, 0.36915323741774586, 
    0.36840108053131881, 0.36765161482399183, 0.36690456211680317, 
    0.36615962281926834, 0.36541649042249713, 0.36467486741056926, 
    0.36393447411596735, 0.36319505563170174, 0.36245638422288845, 
    0.36171826513441541, 0.36098053544867509, 0.36024306457383409, 
    0.3595057555832038, 0.35876854039477724, 0.35803137848177757, 
    0.35729425085020255, 0.3565571551237956, 0.35582010254816732, 
    0.35508311369195306, 0.35434621482397788, 0.35360943292137709, 
    0.35287279771540686, 0.3521363366930958, 0.35140007863266287, 
    0.35066405474414114, 0.3499283016674819, 0.349192868832915, 
    0.34845782054466212, 0.34772323767459179, 0.34698921553550144, 
    0.34625586132246039, 0.34552329023812339, 0.34479162316260148, 
    0.34406098118421197, 0.34333148694115107, 0.34260325912583356, 
    0.34187641160934612, 0.34115104892289555, 0.34042726514025734, 
    0.33970514121659434, 0.33898474670365047, 0.338266142075902, 
    0.33754938406828128, 0.33683453175881301, 0.3361216472128068, 
    0.3354107975690227, 0.33470205364964806, 0.33399548392919992, 
    0.33329115394299774, 0.33258912289295534, 0.33188944179124369, 
    0.33119215486151643, 0.33049730300357827, 0.32980492602124317, 
    0.32911507058301437, 0.32842779334281486, 0.32774316454851732, 
    0.32706127002598218, 0.32638220915525429, 0.3257060964564607, 
    0.32503305463679721, 0.32436321160170639, 0.32369669235938164, 
    0.32303361229466121, 0.32237407073441748, 0.32171814167182389, 
    0.32106587058524588, 0.32041727224667932, 0.31977233153252627, 
    0.31913100667210653, 0.31849323450926481, 0.31785893437399981, 
    0.31722801331037398, 0.31660036983308221, 0.31597590026947314, 
    0.31535450132128962, 0.31473607569054474, 0.31412053665646533, 
    0.31350781111080822, 0.31289784094656764, 0.31229058476709576, 
    0.31168601390225648, 0.31108411001384562, 0.31048485859185537, 
    0.30988824422779804, 0.3092942456127834, 0.30870283292073364, 
    0.30811396748325937, 0.30752760092914661, 0.30694367737539413, 
    0.30636213788717381, 0.30578292306708776, 0.3052059752452379, 
    0.3046312446401257, 0.30405869253565421, 0.30348829251911669, 
    0.30292003332136402, 0.30235391769813441, 0.30178996241805911, 
    0.30122819709735499, 0.30066866143706444, 0.30011140359309707, 
    0.29955647597236584, 0.29900393346269016, 0.29845383365060829, 
    0.29790623592657745, 0.2973612055421207, 0.29681881788540099, 
    0.29627916021346767, 0.29574233370591119, 0.29520845228351922, 
    0.2946776399330312, 0.29415002669098195, 0.2936257430805676, 
    0.29310491385829479, 0.29258765200321546, 0.29207406098324529, 
    0.29156423343211502, 0.29105825297046362, 0.29055619664637278, 
    0.29005813841203815, 0.28956415113138312, 0.28907431237806924, 
    0.28858870497218242, 0.288107417615801, 0.28763054205427191, 
    0.28715817036095259, 0.2866903883140377, 0.28622727063731507, 
    0.28576887531003187, 0.2853152360428805, 0.28486636364319484, 
    0.28442224418165951, 0.28398283976436473, 0.28354809037355516, 
    0.28311791262929975, 0.28269219904699022, 0.28227081375438023, 
    0.28185358981959346, 0.2814403224180072, 0.28103076722186898, 
    0.28062464128734665, 0.28022162408705642, 0.27982136537308494, 
    0.27942349137180189, 0.27902761234572893, 0.27863332930487972, 
    0.27824023861692104, 0.27784793848809558, 0.27745603380391543, 
    0.27706414548419733, 0.27667191748642367, 0.27627902326869597, 
    0.27588516981829969, 0.27549009790152712, 0.27509357780578708, 
    0.27469540725905639, 0.27429540296782678, 0.27389339561887183, 
    0.27348922666154057, 0.27308274415275541, 0.27267380347339326, 
    0.27226226438354939, 0.27184799037345636, 0.27143084803194617, 
    0.27101070434394059, 0.27058742728128482, 0.2701608854992068, 
    0.26973094632889716, 0.26929748201811649, 0.26886037082004299, 
    0.26841950106411877, 0.26797477731055164, 0.26752612158420253, 
    0.2670734768332344, 0.26661680623542766, 0.26615608925321155, 
    0.26569131864798384, 0.26522249728995073, 0.26474963048011679, 
    0.26427272560556619, 0.26379178360235389, 0.26330679747092911, 
    0.2628177500903508, 0.26232461177626898, 0.26182734177258488, 
    0.2613258923904056, 0.2608202099713805, 0.26031024247928647, 
    0.25979594221602098, 0.25927727381975146, 0.25875422086683186, 
    0.25822678892626189, 0.25769501191074112, 0.25715895403919176, 
    0.25661871435596501, 0.25607442938014946, 0.25552627573739045, 
    0.25497447271526497, 0.2544192830275317, 0.25386101146340306, 
    0.25330000318038176, 0.25273663753469111, 0.2521713232354732, 
    0.25160448864629859, 0.25103657832708559, 0.25046804548896173, 
    0.24989934678732567, 0.24933094008791248, 0.24876328389765273, 
    0.2481968346088427, 0.24763204522219423, 0.24706936075490799, 
    0.24650921596708503, 0.24595202830420451, 0.24539819937111049, 
    0.24484810746607591, 0.24430210902081401, 0.24376053889435817, 
    0.24322371328613582, 0.24269193208521248, 0.24216548134706542, 
    0.2416446352027426, 0.24112965655307439, 0.24062079428655278, 
    0.24011827941967678, 0.23962232358392993, 0.23913311532986273, 
    0.23865081835745039, 0.23817556932086947, 0.23770747756212166, 
    0.23724662245595166, 0.2367930550291712, 0.23634679903925829, 
    0.23590785193400646, 0.2354761889981038, 0.23505176770256508, 
    0.23463453065305864, 0.23422440693917021, 0.23382131340487916, 
    0.23342515405457617, 0.23303581514187036, 0.23265316133459016, 
    0.2322770314282584, 0.23190723674692015, 0.23154355696511075, 
    0.23118574517344309, 0.23083352777179619, 0.2304866088964567, 
    0.23014467557778029, 0.22980740250624249, 0.2294744589347236, 
    0.22914551099826933, 0.22882022604728336, 0.22849827625173452, 
    0.2281793412255014, 0.22786310984387614, 0.22754927995889368, 
    0.22723756204253137, 0.22692767842100001, 0.22661936706451069, 
    0.22631238330258896, 0.22600649993984512, 0.22570150953940438, 
    0.22539722653926061, 0.22509348549116606, 0.22479014416000898, 
    0.22448707775422697, 0.22418418269371354, 0.22388137062655294, 
    0.22357856627527761, 0.22327570191700491, 0.22297271571764496, 
    0.2226695481798743, 0.22236614005691979, 0.22206243005763424, 
    0.22175835502183641, 0.22145384914479105, 0.2211488438656197, 
    0.22084326903046317, 0.22053705303175275, 0.22023012376749251, 
    0.21992241124201295, 0.21961385148032284, 0.21930439088105047, 
    0.21899399168891523, 0.21868263462711543, 0.21837032137300508, 
    0.21805707463424573, 0.2177429375765344, 0.21742797065861197, 
    0.21711225023361935, 0.21679586551008764, 0.21647891378286616, 
    0.21616149348746963, 0.21584369847579288, 0.21552561394517566, 
    0.21520730986717468, 0.21488884142977224, 0.21457024988214435, 
    0.21425156680049937, 0.21393281586769936, 0.2136140138493878, 
    0.21329517034036291, 0.21297628737246266, 0.21265735460013946, 
    0.2123383478923839, 0.2120192283611706, 0.21169994313989501, 
    0.21138042387142505, 0.21106058987670218, 0.21074034796435784, 
    0.2104195974844863, 0.21009823223514659, 0.20977614739448178, 
    0.20945324392084536, 0.2091294319057399, 0.20880463471890878, 
    0.2084787897222169, 0.20815184905651241, 0.20782377958620907, 
    0.20749456049621937, 0.20716418506025935, 0.2068326593514718, 
    0.20650000182212458, 0.20616624322450197, 0.20583142605416457, 
    0.20549560218631283, 0.20515882768743457, 0.20482115931573272, 
    0.20448264898300195, 0.20414333425083075, 0.20380323639957318, 
    0.20346235370867324, 0.20312066460657052, 0.20277812792868211, 
    0.20243468970546244, 0.20209028905317494, 0.20174486704609623, 
    0.20139837382172054, 0.20105077594422144, 0.20070205906603072, 
    0.20035223215142101, 0.20000132451405872, 0.19964938551837152, 
    0.19929648285848184, 0.19894269873608825, 0.19858812817234833, 
    0.19823287861876829, 0.19787706628634266, 0.19752081071566557, 
    0.19716423332553559, 0.19680744969487687, 0.19645056816292333, 
    0.19609368507405431, 0.19573688621825061, 0.1953802502194128, 
    0.1950238537487653, 0.19466777817558059, 0.19431211656267866, 
    0.19395697671012813, 0.1936024809835668, 0.19324876822983103, 
    0.19289599174155639, 0.19254431760126012, 0.19219391924189233, 
    0.19184497535552775, 0.191497666777872, 0.19115216953397846, 
    0.19080864897367356, 0.1904672597043261, 0.1901281387146066, 
    0.18979140435546094, 0.1894571505562774, 0.18912544285909524, 
    0.1887963159822155, 0.18846976802203308, 0.18814575768748726, 
    0.18782420143831127, 0.18750496936701128, 0.18718788496784078, 
    0.1868727274002922, 0.18655923512906358, 0.18624710741805503, 
    0.18593601223452916, 0.18562559176636625, 0.18531547078997895, 
    0.18500526358198682, 0.18469458381759721, 0.18438305119235046, 
    0.18407029829221397, 0.18375597887505848, 0.1834397728899736, 
    0.18312139101366331, 0.18280058022561449, 0.1824771223146561, 
    0.18215083978213503, 0.18182159402797224, 0.18148928503605066, 
    0.18115385423143282, 0.18081528101160071, 0.18047358564738775, 
    0.18012882954648976, 0.179781116650923, 0.17943059758676777, 
    0.17907746810586717, 0.17872197127528092, 0.17836439323913822, 
    0.17800505824209109, 0.1776443201223035, 0.17728255467862825, 
    0.17692015091798355, 0.17655750050783373, 0.17619498666102465, 
    0.17583297678718632, 0.17547181222198752, 0.17511180112558292, 
    0.17475321336923461, 0.17439627638935018, 0.17404117080880233, 
    0.17368803563973126, 0.17333696663914952, 0.17298802203258648, 
    0.17264122332183135, 0.17229656064790944, 0.17195399171818931, 
    0.1716134444461542, 0.17127481369397643, 0.17093796122447438, 
    0.17060271654011239, 0.17026887843908609, 0.16993621344088666, 
    0.16960446072660318, 0.16927333471805503, 0.16894252898235212, 
    0.16861172419607659, 0.16828059204180346, 0.1679488012728122, 
    0.1676160247461361, 0.1672819454588611, 0.16694626523502298, 
    0.16660871479299807, 0.16626906136939987, 0.16592711506954522, 
    0.16558273539283194, 0.16523583236725861, 0.16488637080687668, 
    0.16453436969085564, 0.16417990041506822, 0.16382308984283236, 
    0.16346411959016249, 0.16310322376754499, 0.16274068910584066, 
    0.1623768541847492, 0.16201210313601244, 0.161646862093065, 
    0.16128159165357098, 0.16091677893580725, 0.16055292994882867, 
    0.16019055952768868, 0.15983018114862041, 0.15947230136542973, 
    0.1591174107950572, 0.15876598159830974, 0.1584184587487607, 
    0.15807525856790369, 0.15773676314446752, 0.15740331638429503, 
    0.15707521699799737, 0.15675271383157383, 0.15643600215221495, 
    0.15612522140142787, 0.15582045576078318, 0.15552173526402285, 
    0.15522904024270046, 0.15494230529901937, 0.15466142635551353, 
    0.15438626480978271, 0.15411665450458265, 0.15385240455501129, 
    0.15359330343912422, 0.15333912257487128, 0.15308961578195743, 
    0.15284452502680165, 0.15260357809134761, 0.15236649114403983, 
    0.15213296841032534, 0.15190270652893703, 0.15167539641520739, 
    0.1514507292226451, 0.15122839762952767, 0.15100809959950581, 
    0.15078954212407883, 0.15057244062550817, 0.1503565217903326, 
    0.15014152094244496, 0.14992718145788955, 0.14971325605744989, 
    0.14949950416853883, 0.14928569180607035, 0.14907159400131689, 
    0.14885699323268328, 0.1486416829783043, 0.14842546980202798, 
    0.14820817823963803, 0.14798965253498783, 0.14776976161518512, 
    0.14754840265392624, 0.14732550556944693, 0.14710103368710717, 
    0.14687498659278045, 0.14664739891302911, 0.14641834301703435, 
    0.14618792797280264, 0.14595629745127628, 0.1457236297107781, 
    0.14549013296663299, 0.14525604382749105, 0.14502162135126859, 
    0.14478714194639045, 0.14455289193846524, 0.14431916161064862, 
    0.14408623961587291, 0.14385440668496874, 0.14362393031811316, 
    0.14339505973541766, 0.14316802627606043, 0.14294303692506025, 
    0.14272027346645336, 0.14249988546614825, 0.14228198975176262, 
    0.14206666683451172, 0.14185395937990625, 0.1416438749935004, 
    0.14143638806414235, 0.1412314422293538, 0.14102895466711773, 
    0.14082882064748431, 0.14063091622666715, 0.1404351036067501, 
    0.14024123462389587, 0.14004915761079773, 0.13985871951455242, 
    0.13966977339283698, 0.13948217943706367, 0.13929580916306003, 
    0.13911055004476691, 0.13892630437777903, 0.13874299191299932, 
    0.13856054936074916, 0.138378931875593, 0.13819810894282056, 
    0.13801806278704992, 0.13783878699331065, 0.13766028374554526, 
    0.13748255915431487, 0.13730562410377692, 0.1371294901194364, 
    0.13695416626169549, 0.13677965713563914, 0.13660595936270215, 
    0.13643305952751714, 0.1362609318900386, 0.13608953618540789, 
    0.13591881365368072, 0.13574868268926971, 0.13557903635481947, 
    0.13540974201983891, 0.135240637147961, 0.1350715301934928, 
    0.1349022043610407, 0.13473241869178515, 0.13456191869493184, 
    0.13439044351887736, 0.13421773371213919, 0.13404353922666495, 
    0.13386762975580518, 0.13368979492884317, 0.13350984744739861, 
    0.13332762607448731, 0.13314299228448065, 0.13295583283084489, 
    0.13276605411505712, 0.13257358217505974, 0.1323783627766838, 
    0.13218036106884981, 0.13197956262032889, 0.1317759730101013, 
    0.13156962119121313, 0.13136056053652859, 0.13114886843258122, 
    0.13093464629347162, 0.13071801512698056, 0.13049911232902603, 
    0.13027808569163271, 0.13005508791358084, 0.1298302715667024, 
    0.12960378955896107, 0.12937579053833748, 0.12914642160697931, 
    0.12891582411786806, 0.12868413292042008, 0.12845147440486832, 
    0.12821796367147456, 0.12798369841714721, 0.12774875839171368, 
    0.12751320473176017, 0.12727707939460839, 0.12704040558932539, 
    0.12680319281469699, 0.12656543635952022, 0.12632712235213817, 
    0.1260882279104715, 0.12584872900879779, 0.12560859663440782, 
    0.12536780385746116, 0.12512632505236204, 0.12488414316709921, 
    0.1246412505889315, 0.12439765471199252, 0.12415338119005002, 
    0.12390847485355957, 0.12366299686473736, 0.12341702078649452, 
    0.12317062463847477, 0.12292388390600918, 0.12267686425822995, 
    0.12242961441334724, 0.12218216433536105, 0.1219345255025449, 
    0.12168668817502987, 0.12143862435419121, 0.12119029141809398, 
    0.12094163589955563, 0.12069259662026971, 0.12044311027554586, 
    0.1201931157894342, 0.11994255610275988, 0.11969138222608541, 
    0.11943955408707557, 0.11918704279664807, 0.11893382836673898, 
    0.11867990314871246, 0.11842526933416016, 0.11816993726801212, 
    0.11791392391747166, 0.11765725002509068, 0.11739993659872898, 
    0.11714200201636624, 0.11688345685852565, 0.116624302290427, 
    0.11636452730000492, 0.11610410287954888, 0.11584298271977603, 
    0.11558110224775635, 0.1153183786511022, 0.11505471370549207, 
    0.11478999787948138, 0.1145241219822503, 0.11425698133633558, 
    0.11398848902635564, 0.113718582796466, 0.11344723414514436, 
    0.11317445415700417, 0.11290029508656825, 0.11262485081049502, 
    0.11234825201691753, 0.11207066181450741, 0.11179227184279293, 
    0.11151329523241055, 0.11123395871386423, 0.1109544995914493, 
    0.11067516166250622, 0.11039619216359779, 0.11011784167435573, 
    0.10984036135968155, 0.10956400597527921, 0.10928903284644001, 
    0.1090157025625208, 0.10874427350952676, 0.10847499813288704, 
    0.1082081192409266, 0.10794386441396393, 0.10768244287127296, 
    0.10742404209697284, 0.10716882702751712, 0.10691694118809913, 
    0.10666851129995394, 0.10642364670141759, 0.10618244116155816, 
    0.1059449761595856, 0.10571131927580768, 0.10548152349702203, 
    0.10525562432852746, 0.10503363562451995, 0.10481554706840968, 
    0.10460132103151183, 0.10439088998652955, 0.1041841543911504, 
    0.10398097951280931, 0.10378120055361428, 0.10358462133253796, 
    0.10339102207221194, 0.10320016632154161, 0.10301181050968995, 
    0.10282571427851864, 0.10264164875235751, 0.10245940126703607, 
    0.10227878048102376, 0.10209961342520224, 0.10192174218135025, 
    0.10174502010386689, 0.10156930628397576, 0.10139446297856003, 
    0.10122035457568608, 0.10104684149620094, 0.10087378242282585, 
    0.10070103822798675, 0.10052846927257834, 0.10035593825408841, 
    0.10018331509737557, 0.1000104800392614, 0.09983732951492004, 
    0.09966377725890975, 0.099489761393265361, 0.099315242702169695, 
    0.099140205336321202, 0.098964652559187211, 0.09878860880553153, 
    0.09861211723036499, 0.098435241325443693, 0.098258059421391028, 
    0.098080670480542143, 0.097903186083935972, 0.097725736061452267, 
    0.097548463440453023, 0.09737152459015265, 0.097195089475464208, 
    0.097019339316817083, 0.096844465009565922, 0.096670662169243041, 
    0.096498131448014196, 0.096327070307637208, 0.096157668326768198, 
    0.095990101999467212, 0.095824532128065548, 0.09566109555048001, 
    0.095499906024287304, 0.095341047632294396, 0.09518457588665849, 
    0.095030518159989696, 0.094878874068075214, 0.094729618367541207, 
    0.094582704706057855, 0.094438069380168535, 0.09429563776742661, 
    0.094155324939968352, 0.094017042195750855, 0.093880699544954052, 
    0.093746207662762843, 0.093613480519526351, 0.093482435782370851, 
    0.093352997803260007, 0.093225092977557031, 0.093098652312030766, 
    0.092973611817188773, 0.092849910188918486, 0.09272749051903631, 
    0.092606301460049653, 0.092486297647624532, 0.092367436557411489, 
    0.092249682686600123, 0.092133006713013041, 0.092017386299734633, 
    0.091902809772760941, 0.091789274357254799, 0.091676790271911612, 
    0.091565375750344277, 0.091455060738297927, 0.091345884309687195, 
    0.09123789006383759, 0.091131123886348697, 0.091025626898342024, 
    0.090921434572310666, 0.090818569344030153, 0.090717043867417135, 
    0.090616857766245174, 0.090517997997135599, 0.090420441080808517, 
    0.090324154503807971, 0.090229100658603095, 0.090135242753644693, 
    0.090042550554886538, 0.089951009688683373, 0.089860624133490871, 
    0.089771421024562592, 0.089683453477958378, 0.089596798767616906, 
    0.089511555257957079, 0.08942784129660937, 0.089345785342414122, 
    0.08926552148622259, 0.089187179524976706, 0.089110877156044446, 
    0.089036711924736667, 0.08896474998653052, 0.088895016843146477, 
    0.088827499814228841, 0.088762142316239551, 0.088698850596302725, 
    0.088637502234097373, 0.088577955343977305, 0.088520056817422546, 
    0.088463656101254798, 0.088408609051979531, 0.088354785697992738, 
    0.088302075759494489, 0.088250389673395185, 0.088199662427270301, 
    0.088149847469128184, 0.088100920499111376, 0.08805287110442285, 
    0.088005693338078256, 0.087959380600463238, 0.087913917035678094, 
    0.087869267125207984, 0.087825376004885811, 0.087782162912856412, 
    0.087739523607552272, 0.087697332952975368, 0.087655449974212693, 
    0.087613726432679839, 0.087572010118893276, 0.087530148556483833, 
    0.087487993586699786, 0.087445402899206603, 0.087402239661468567, 
    0.087358372901700079, 0.087313674635516175, 0.087268021670822968, 
    0.08722129511756592, 0.087173377319369222, 0.087124157132170629, 
    0.087073525922587214, 0.087021375520614591, 0.08696760399201757, 
    0.086912108093811752, 0.086854791563091574, 0.086795562366638671, 
    0.086734333554148071, 0.086671029712258527, 0.086605587445504159, 
    0.086537956490883888, 0.086468101301612282, 0.086396001402864714, 
    0.086321656340400774, 0.086245088385797308, 0.086166345915240999, 
    0.086085503694750168, 0.086002669916367125, 0.085917987966897744, 
    0.085831634698922216, 0.085743819800710899, 0.085654784622711241, 
    0.085564796684122826, 0.085474145615664535, 0.085383133468578412, 
    0.085292065283947949, 0.085201241806334926, 0.085110948767527256, 
    0.085021454226203441, 0.084933000497324454, 0.08484580244037862, 
    0.084760039787454888, 0.084675858475904489, 0.084593364023373682, 
    0.084512627121649822, 0.084433687561597429, 0.084356566254511198, 
    0.08428126695482549, 0.084207784398059787, 0.084136107350677614, 
    0.084066219578215903, 0.083998099938854459, 0.083931724657699922, 
    0.08386706471630434, 0.083804087868320221, 0.083742753600038994, 
    0.083683009591383861, 0.083624783108511749, 0.083567977675626251, 
    0.083512466279139067, 0.083458093213905238, 0.083404677077626027, 
    0.083352014959359483, 0.08329988778051152, 0.083248067404577936, 
    0.083196322276065368, 0.083144424667108516, 0.083092149348107588, 
    0.083039279933180152, 0.082985606917151136, 0.082930928650258418, 
    0.082875052872968577, 0.082817800494728977, 0.082759010795037918, 
    0.082698543189990703, 0.082636282403663747, 0.082572142021090048, 
    0.082506067066051111, 0.082438034575683133, 0.082368049498253007, 
    0.082296142562039057, 0.082222367732186261, 0.082146792603075572, 
    0.08206949662862642, 0.081990563036596673, 0.081910078951865015, 
    0.081828133620382423, 0.081744809155213233, 0.081660181527750272, 
    0.081574315449180049, 0.081487260068349873, 0.08139905339147907, 
    0.081309724530495342, 0.081219303007551036, 0.081127826472003645, 
    0.081035354850164443, 0.080941980185942994, 0.080847832674161513, 
    0.080753088096485168, 0.080657967034579378, 0.080562731680129562, 
    0.080467682194509532, 0.080373151050059793, 0.080279496960453986, 
    0.080187103028455886, 0.080096367385239786, 0.080007700759509207, 
    0.079921519558704204, 0.079838243432784825, 0.079758287926745025, 
    0.079682060247514383, 0.079609952167626605, 0.079542335578863116, 
    0.079479558287466445, 0.079421937878937754, 0.079369757829124366, 
    0.079323258813762162, 0.079282635731621698, 0.079248030926855062, 
    0.079219529293678329, 0.079197159806596307, 0.079180897405395467, 
    0.079170664500105792, 0.07916634202037863, 0.079167774639481589, 
    0.079174780833607461, 0.079187155908636106, 0.07920468052787763, 
    0.079227121442528289, 0.079254233521783679, 0.079285754920416757, 
    0.079321408187734296, 0.079360894199632714, 0.07940389307185744, 
    0.079450065111086349, 0.079499051612785865, 0.079550478570328528, 
    0.079603958816433992, 0.079659090244381781, 0.079715456235407697, 
    0.079772628988281247, 0.079830171116303042, 0.079887636496310324, 
    0.07994457718193354, 0.080000544776420379, 0.080055093670442723, 
    0.080107780287146282, 0.080158173327444251, 0.080205849690320949, 
    0.080250406980534664, 0.080291468986829151, 0.080328698398351828, 
    0.080361807689605616, 0.080390565313953985, 0.080414803431065149, 
    0.080434420230322115, 0.080449376362119199, 0.08045968802530766, 
    0.08046541820792924, 0.080466664961363357, 0.080463552235398889, 
    0.080456223616630393, 0.080444835540785659, 0.080429563977189783, 
    0.080410604091628063, 0.08038817548339719, 0.080362520568313153, 
    0.080333905112066326, 0.080302616783175573, 0.080268958703758289, 
    0.08023324045899223, 0.080195772526364215, 0.080156857833693293, 
    0.080116782373765225, 0.08007581333677033, 0.080034197118109093, 
    0.079992165811678284, 0.079949941922866669, 0.079907744504727637, 
    0.079865793383122358, 0.079824311020836494, 0.079783523866054654, 
    0.079743658680747426, 0.079704940169533098, 0.079667586545325728, 
    0.079631805916512102, 0.079597788446618772, 0.079565700551818774, 
    0.07953567568912577, 0.079507812167627617, 0.079482168112543439, 
    0.079458760471362244, 0.079437568091497407, 0.079418532802300365, 
    0.079401567352146971, 0.079386555491683816, 0.079373355589702807, 
    0.079361805317579373, 0.079351721604760728, 0.079342904954933582, 
    0.079335141922789454, 0.079328211155812636, 0.079321887515935177, 
    0.079315945744357089, 0.079310157399473641, 0.079304287999209633, 
    0.079298091026451453, 0.0792913008523492, 0.079283623476011728, 
    0.079274727064883102, 0.079264233916749, 0.079251718472701266, 
    0.079236705703769575, 0.079218675580425515, 0.079197069262772229, 
    0.07917129819055857, 0.079140761928128286, 0.079104867899204956, 
    0.079063050118133665, 0.079014789707552782, 0.078959632973344004, 
    0.078897202625076504, 0.078827207819538669, 0.078749448732458635, 
    0.078663819305998625, 0.078570301254172442, 0.078468954655880635, 
    0.078359908082999558, 0.078243348295414433, 0.07811950127596097, 
    0.077988625638222564, 0.077851001366218364, 0.07770692053978985, 
    0.077556683229602894, 0.077400591242322347, 0.077238950289367198, 
    0.077072070439615503, 0.07690026890315306, 0.076723876687029458, 
    0.076543245047035316, 0.076358751369140859, 0.07617080579732799, 
    0.075979854702032446, 0.075786375846947293, 0.0755908761051126, 
    0.075393883306655834, 0.075195939007634133, 0.074997586628718915, 
    0.074799362660899579, 0.074601788686312981, 0.074405365228681145, 
    0.074210565005020324, 0.074017825778898316, 0.07382754747261687, 
    0.073640090021863128, 0.073455774677589791, 0.07327489103755036, 
    0.073097707989088948, 0.072924485996809146, 0.072755490370220097, 
    0.072590992380392239, 0.072431260411414802, 0.072276548912052013, 
    0.072127084415384263, 0.071983043646910952, 0.071844545454177164, 
    0.071711639479988959, 0.07158430765611945, 0.071462464691893213, 
    0.071345965551193741, 0.071234617700771857, 0.071128201214189557, 
    0.071026484512053373, 0.07092923975291017, 0.070836259357249631, 
    0.070747365804527382, 0.070662414805293269, 0.070581301889042325, 
    0.070503952867784353, 0.070430322485455998, 0.070360386454608903, 
    0.070294138019362365, 0.070231585812323166, 0.070172752778262584, 
    0.070117676631997597, 0.070066402314332268, 0.070018980646042422, 
    0.069975458193578977, 0.069935864439320983, 0.069900204440112773, 
    0.069868448619408066, 0.069840540041693391, 0.069816385569550249, 
    0.069795863559338672, 0.069778823482519889, 0.06976509232770628, 
    0.069754478972484532, 0.06974677699023546, 0.069741768114885777, 
    0.069739217991702046, 0.069738886137975742, 0.069740511312033016, 
    0.069743816849451329, 0.069748509903144337, 0.069754283558154356, 
    0.06976081790199766, 0.069767782765847094, 0.069774842964538966, 
    0.06978166668494995, 0.069787927183981857, 0.069793314460020933, 
    0.069797536112450001, 0.069800327581960891, 0.069801451981667276, 
    0.069800705980563621, 0.069797917328485296, 0.069792943835653293, 
    0.069785675704494329, 0.069776035646979748, 0.069763981232132469, 
    0.069749508250245368, 0.069732653130367042, 0.069713498099327087, 
    0.069692166112415355, 0.069668813361960458, 0.069643627287942295, 
    0.069616807510940987, 0.069588558676301662, 0.069559086906960582, 
    0.069528593278288392, 0.069497264174518944, 0.06946527969908467, 
    0.069432811680373199, 0.06940002523787113, 0.069367079542026575, 
    0.069334127912636254, 0.069301323072237894, 0.069268812633582227, 
    0.069236743576608403, 0.069205256914821781, 0.069174488732488285, 
    0.069144568462007922, 0.069115618824145339, 0.069087752691608911, 
    0.069061077339942503, 0.06903568821142983, 0.069011677704856514, 
    0.068989130611415594, 0.06896812776597222, 0.068948745308294021, 
    0.068931060988549328, 0.068915144296017083, 0.068901053259091474, 
    0.068888825475023133, 0.068878469191954783, 0.068869961361695778, 
    0.068863244432570664, 0.068858231342871584, 0.068854810486216861, 
    0.068852860480440856, 0.068852258741104524, 0.068852889563877417, 
    0.068854649763783568, 0.068857444381028338, 0.068861180122181495, 
    0.068865766591059321, 0.06887110529457087, 0.06887708948877895, 
    0.068883592525658163, 0.068890464291320896, 0.068897518949974493, 
    0.068904530425487623, 0.068911221850840629, 0.06891727341742937, 
    0.068922325562026918, 0.068925985126609274, 0.068927835741457388, 
    0.068927447013848162, 0.068924391501353252, 0.068918247598468194, 
    0.068908613438971963, 0.06889511261445283, 0.068877397983116248, 
    0.068855161049704974, 0.068828136926991759, 0.068796110066936672, 
    0.068758925293459811, 0.068716498155086472, 0.068668826090977297, 
    0.068616008115116214, 0.068558249994431816, 0.068495861093427854, 
    0.068429224371876568, 0.068358758964059851, 0.068284870489558044, 
    0.068207924074978471, 0.068128245681679689, 0.068046132233158863, 
    0.067961874293181443, 0.067875773366660577, 0.06778815654733418, 
    0.067699386894093411, 0.067609865329026242, 0.067520034835205966, 
    0.067430382202397721, 0.067341435153890933, 0.067253760082332817, 
    0.067167958522083793, 0.06708465219489744, 0.06700447991360188, 
    0.066928080600116985, 0.066856080164274509, 0.066789082564248523, 
    0.066727662878275779, 0.066672366673318523, 0.066623708858553177, 
    0.066582177916645058, 0.066548235153552571, 0.066522314601179647, 
    0.066504825413965449, 0.066496141242949267, 0.066496600367759853, 
    0.066506494451959275, 0.06652606493109646, 0.066555492850092893, 
    0.066594896460834024, 0.066644330663471182, 0.066703783896601573, 
    0.066773184660134044, 0.066852400447412724, 0.066941249921785448, 
    0.067039516233991334, 0.067146952783077501, 0.067263303769532296, 
    0.067388312679333026, 0.067521739883363838, 0.067663365536131878, 
    0.067813000742764112, 0.067970487762857384, 0.068135695735987836, 
    0.068308526531955016, 0.068488904269465162, 0.068676778480824097, 
    0.068872117900164981, 0.069074912222758009, 0.069285165586636013, 
    0.069502900175058793, 0.069728150841605357, 0.069960965485395016, 
    0.070201404919629104, 0.07044954030370533, 0.070705450969406752, 
    0.070969231967199467, 0.071240994205245364, 0.071520862067351296, 
    0.071808973956991484, 0.072105471905621235, 0.072410492485293923, 
    0.072724155710735996, 0.073046547847067045, 0.073377712379384175, 
    0.073717643645314912, 0.07406628221301817, 0.074423516592410338, 
    0.074789176875914201, 0.075163042366391514, 0.075544835915778014, 
    0.075934230207006362, 0.076330847160927889, 0.076734259515596481, 
    0.077143993379571951, 0.077559533572158113, 0.07798032997802401, 
    0.078405794305514864, 0.078835301334359745, 0.079268180721986325, 
    0.079703715843173109, 0.080141147840490215, 0.080579679903861973, 
    0.081018501674610846, 0.081456799544013483, 0.081893772361570777, 
    0.082328643813230962, 0.082760672463213517, 0.083189157036762162, 
    0.08361343361192812, 0.084032877311875115, 0.084446903088190084, 
    0.084854956349031091, 0.085256512239696741, 0.085651069267716554, 
    0.08603814692692241, 0.086417286841410035, 0.086788051202867103, 
    0.087150032730145946, 0.087502859232682237, 0.087846200517318784, 
    0.088179780929528079, 0.088503372808592759, 0.088816794523068981, 
    0.089119902946119739, 0.089412592512146186, 0.08969477128116396, 
    0.089966359626229245, 0.090227281286053951, 0.090477449994880416, 
    0.090716778885377991, 0.090945179928413986, 0.091162574033953142, 
    0.091368906079063797, 0.091564151978576439, 0.091748328384590211, 
    0.091921504858541697, 0.092083806616993516, 0.092235416315953778, 
    0.092376582280849495, 0.092507619920349157, 0.092628913020615586, 
    0.092740919226475788, 0.092844168028632407, 0.092939250198286902, 
    0.093026812096066364, 0.093107533996192302, 0.093182115388091957, 
    0.093251255396320135, 0.093315623276852125, 0.09337585167706354, 
    0.093432520616098289, 0.0934861467419007, 0.093537202294784239, 
    0.093586112277849715, 0.09363328191918055, 0.093679097752293189, 
    0.0937239407812685, 0.093768181358486052, 0.093812149396875988, 
    0.09385612033766122, 0.093900293687206815, 0.093944772951968528, 
    0.093989563603034718, 0.09403456556167103, 0.094079577099769884, 
    0.094124290298814806, 0.094168310438002861, 0.094211175981359779, 
    0.094252389373204057, 0.094291442104612724, 0.094327851658334308, 
    0.094361176792598631, 0.094391029569440954, 0.094417081087238341, 
    0.094439057901649262, 0.094456737118972484, 0.094469933082739724, 
    0.094478477692122462, 0.09448222280824424, 0.094481018071631145, 
    0.094474708544698818, 0.094463136680057722, 0.094446146527402519, 
    0.094423607605100129, 0.094395431260888243, 0.094361598789337323, 
    0.094322185746213746, 0.09427738524216743, 0.094227532942690179, 
    0.094173097463550681, 0.094114683941516578, 0.094053023182575621, 
    0.093988961139495703, 0.093923444698471345, 0.093857495051154594, 
    0.093792209329762455, 0.093728732478698132, 0.093668243292028844, 
    0.093611931104213217, 0.093560961852920996, 0.09351645491386007, 
    0.093479457492616574, 0.09345091437578773, 0.09343164418469449, 
    0.093422330319123559, 0.09342349966663048, 0.093435510068039559, 
    0.09345854851630836, 0.093492628204607395, 0.093537593637579519, 
    0.093593118903053232, 0.093658725953065833, 0.093733787836611696, 
    0.093817554316240725, 0.09390915029576373, 0.094007610111214002, 
    0.094111879726843164, 0.094220846437895592, 0.094333350325485746, 
    0.094448207974445642, 0.094564217787564644, 0.094680169612238407, 
    0.094794863189827452, 0.094907092341293242, 0.095015682113077357, 
    0.095119508996596491, 0.095217534454928601, 0.095308837001273364, 
    0.09539264400102189, 0.095468357206838522, 0.09553557113956275, 
    0.09559408649663298, 0.095643918495657634, 0.09568529189807766, 
    0.095718621500433518, 0.095744487798018404, 0.095763580856887895, 
    0.095776642887955232, 0.095784393757181646, 0.095787471488554918, 
    0.095786372716227558, 0.095781418034642921, 0.095772736598552746, 
    0.095760256482218725, 0.095743729521300738, 0.095722769584866363, 
    0.095696881531678879, 0.095665500001295728, 0.095628019563538641, 
    0.095583814270396611, 0.095532253208567189, 0.095472725677966885, 
    0.095404654584078277, 0.095327524009964013, 0.095240882262851212, 
    0.095144341033850013, 0.095037580530703533, 0.09492033447272584, 
    0.094792383109725376, 0.094653555357628219, 0.094503722415550037, 
    0.094342802180663488, 0.09417077334872577, 0.093987678257545559, 
    0.093793637432736152, 0.093588847045701293, 0.093373577031443444, 
    0.09314817000437127, 0.092913025711162972, 0.092668614566282864, 
    0.09241547018086041, 0.09215419473176055, 0.091885464847658652, 
    0.091610028266470814, 0.091328692339948531, 0.091042321033746973, 
    0.090751810101539557, 0.090458057252856286, 0.090161935344265379, 
    0.089864293919856328, 0.089565902642055273, 0.089267438680632027, 
    0.088969457620942369, 0.088672365931261668, 0.088376409843027429, 
    0.088081683611827138, 0.087788145145043753, 0.087495643045117408, 
    0.087203934989381782, 0.086912713858998042, 0.08662164620474358, 
    0.086330397937568817, 0.086038643833478534, 0.085746075504673433, 
    0.085452429938762328, 0.085157466692736355, 0.08486097487142609, 
    0.084562761509294745, 0.084262636068440103, 0.083960401055815551, 
    0.083655851161450065, 0.083348750047040163, 0.083038840776931896, 
    0.082725838575761934, 0.082409412309684238, 0.082089205181527236, 
    0.081764830251680284, 0.081435863182582321, 0.081101859484757954, 
    0.080762344308408021, 0.080416850495701742, 0.080064914279883992, 
    0.079706097903589013, 0.079339983122053565, 0.078966173271187323, 
    0.078584302809095563, 0.078194039850207744, 0.077795095312857512, 
    0.077387262202815846, 0.076970447762921168, 0.076544712342881516, 
    0.076110280729165911, 0.075667581011010288, 0.075217255456523913, 
    0.074760139763356118, 0.074297274422294474, 0.073829892861729515, 
    0.073359337320722168, 0.072887060010373303, 0.072414510872590723, 
    0.071943108075298065, 0.071474138747054883, 0.071008711498696128, 
    0.070547710963832583, 0.070091741490803813, 0.069641128538402458, 
    0.069195879076603795, 0.068755732070122658, 0.068320161343934122, 
    0.067888422932907311, 0.067459617683668135, 0.067032721844967544, 
    0.066606658416869705, 0.066180320044942925, 0.065752633136900163, 
    0.065322560065202193, 0.064889069298658841, 0.064451151378907098, 
    0.064007759154231209, 0.063557810915299148, 0.063100158983294824, 
    0.062633578905602325, 0.062156768677466216, 0.061668333346125724, 
    0.061166847101558224, 0.060650853666282645, 0.060118917028776017, 
    0.059569682183237195, 0.059001949041604815, 0.058414693224495572, 
    0.057807165904125386, 0.057178895325994225, 0.056529754081154925, 
    0.055859916317390214, 0.055169844630396023, 0.054460289666794282, 
    0.053732306177950245, 0.052987205584632421, 0.052226543439328386, 
    0.051452083103388696, 0.050665740824736148, 0.04986953838150756, 
    0.04906553105676361, 0.048255756743650957, 0.047442208192071469, 
    0.046626882617586983, 0.045811844933708136, 0.044999246344148404, 
    0.044191448328587429, 0.043391131474799241, 0.042601287679879397, 
    0.041825274334368723, 0.041066633787785363, 0.040328930886199738, 
    0.039615676171970579, 0.038930297258220489, 0.038276092674559704, 
    0.037656287971575948, 0.03707406535913528, 0.036532513149935358, 
    0.036034774196212357, 0.03558385846393361, 0.035182697254181453, 
    0.03483402108962496, 0.034540256970190392, 0.034303415763273601, 
    0.034125072490306205, 0.034006174491211398, 0.033947015697592342, 
    0.033947029057569564, 0.034004967157740956, 0.034118988573319138, 
    0.034286875454945388,
  // Fqt-F(1, 0-1999)
    1, 0.9994840397665119, 0.997941456186896, 0.99538818742700441, 
    0.9918504270609948, 0.98736390348575465, 0.98197293445963629, 
    0.97572930901168742, 0.96869105260657351, 0.96092113322520589, 
    0.95248615786570467, 0.94345510521503406, 0.93389813177877967, 
    0.92388547157748013, 0.91348645231816916, 0.90276863403600827, 
    0.89179706986427965, 0.88063369393592172, 0.86933682788771405, 
    0.85796079585361862, 0.84655564907986569, 0.83516698736136452, 
    0.82383587148445492, 0.81259881749215701, 0.80148786102934444, 
    0.79053068185150632, 0.77975077618189692, 0.76916766624577815, 
    0.75879712952971801, 0.74865145888796236, 0.73873973818802152, 
    0.72906812508206353, 0.71964014389468756, 0.71045696716386419, 
    0.70151769115572604, 0.69281959918832847, 0.68435840617754762, 
    0.67612849217695037, 0.66812312109369998, 0.66033464618991022, 
    0.65275470266766511, 0.64537439682612974, 0.63818447614700002, 
    0.63117549551229246, 0.6243379632419217, 0.61766247448599731, 
    0.61113982443657622, 0.60476110403877692, 0.59851777707894016, 
    0.59240174094913201, 0.58640537691879879, 0.5805215808041152, 
    0.574743787395529, 0.56906598493156113, 0.5634827128400991, 
    0.55798905758677797, 0.55258063399945312, 0.54725356163153782, 
    0.54200443597900017, 0.53683028995610249, 0.53172855968363864, 
    0.52669704033444043, 0.52173384394152422, 0.51683736143538705, 
    0.51200621609503827, 0.50723923534816073, 0.5025354185889257, 
    0.49789391044524051, 0.49331397548547173, 0.48879497266929178, 
    0.4843363324300668, 0.47993752951511531, 0.47559806145949757, 
    0.4713174191923698, 0.46709506535907797, 0.46293040878234282, 
    0.4588227808610319, 0.45477141968917018, 0.45077544931513852, 
    0.4468338730464711, 0.44294556480996772, 0.43910926693453972, 
    0.43532359897753264, 0.43158706474362857, 0.4278980639486869, 
    0.42425491456397857, 0.42065587162739076, 0.41709915679045778, 
    0.41358298206881805, 0.41010558268620562, 0.40666524600002052, 
    0.40326033603945677, 0.39988932386238096, 0.39655080443418517, 
    0.39324352451006328, 0.38996639926732413, 0.38671853285058982, 
    0.38349923582486856, 0.38030803165127752, 0.37714466080466758, 
    0.37400907728471666, 0.37090144564833089, 0.36782212756803068, 
    0.36477167038496017, 0.36175079012254147, 0.35876035077246743, 
    0.3558013431150342, 0.35287485682877012, 0.3499820600083508, 
    0.34712417099426507, 0.34430243387258869, 0.34151809103407438, 
    0.33877236310945896, 0.33606642390772573, 0.33340138463938124, 
    0.33077827314552838, 0.32819802150893412, 0.32566145050806372, 
    0.32316926443457705, 0.32072203840363744, 0.31832021898999674, 
    0.31596411812063435, 0.31365391536686843, 0.31138965747973041, 
    0.3091712523525792, 0.30699846872428177, 0.30487092773359503, 
    0.30278810156676988, 0.30074931040774999, 0.29875372291739533, 
    0.2968003535855912, 0.29488806895468461, 0.29301559201537325, 
    0.29118151109766327, 0.28938428580264297, 0.28762226145046682, 
    0.28589368208149701, 0.2841967059452879, 0.28252942229406069, 
    0.28088987311673103, 0.27927607054928566, 0.27768601917656954, 
    0.27611773965566483, 0.27456929249961204, 0.273038793984554, 
    0.27152443938771115, 0.27002451880304507, 0.26853743494123089, 
    0.26706171000654405, 0.26559600094012165, 0.26413910412604624, 
    0.26268995860302191, 0.26124765069431422, 0.25981140664364799, 
    0.25838059297166699, 0.25695470643608237, 0.25553336533650917, 
    0.25411629343758207, 0.25270331042789224, 0.25129431147596193, 
    0.24988925955682392, 0.24848815953244299, 0.24709104747744595, 
    0.2456979764386672, 0.24430900784191292, 0.24292420174454726, 
    0.24154361480958308, 0.24016729933099346, 0.23879530997140505, 
    0.23742771535071702, 0.23606461359910824, 0.23470614466561016, 
    0.23335249569990207, 0.23200390130426621, 0.23066063574902546, 
    0.22932300259085303, 0.22799132250871079, 0.22666592065904556, 
    0.22534712177740363, 0.22403523932550318, 0.22273057058859863, 
    0.22143338825363518, 0.22014393954430697, 0.2188624403133046, 
    0.21758907684836731, 0.21632401051241745, 0.2150673803738255, 
    0.21381930878029443, 0.2125799083135525, 0.21134928814822929, 
    0.21012755703874833, 0.20891482600126912, 0.20771121193186429, 
    0.20651683425295483, 0.20533181799350556, 0.20415628913656833, 
    0.20299037298700287, 0.2018341882054972, 0.20068784531020059, 
    0.19955144565985578, 0.19842507511508975, 0.19730880491992445, 
    0.19620268902207699, 0.19510675956957135, 0.19402102338004246, 
    0.1929454591085184, 0.19188001750919634, 0.190824613849605, 
    0.18977913839760438, 0.18874345068426818, 0.18771739035930016, 
    0.18670078390017786, 0.18569344956394407, 0.18469520556100463, 
    0.1837058744370984, 0.18272529308182431, 0.1817533167108796, 
    0.18078982703830107, 0.17983474103192673, 0.17888801453802206, 
    0.17794964594579687, 0.17701967367795257, 0.17609817736555877, 
    0.17518526668651821, 0.17428107822110592, 0.17338576192494426, 
    0.17249946954543321, 0.17162234018955266, 0.17075448293174711, 
    0.1698959679655363, 0.16904680945429462, 0.16820695399134872, 
    0.16737627106524541, 0.1665545426187372, 0.16574145793233197, 
    0.16493661158939618, 0.16413950718625736, 0.16334955651132349, 
    0.16256609502731223, 0.16178838966188747, 0.16101565457805073, 
    0.16024706977198841, 0.1594817983570764, 0.15871900278997389, 
    0.15795785930419584, 0.15719756886828049, 0.15643736270286743, 
    0.15567651045995337, 0.15491432356942056, 0.15415015619432845, 
    0.15338340652623114, 0.15261351778694621, 0.15183997870149515, 
    0.15106232443505371, 0.1502801426363809, 0.1494930772909881, 
    0.14870083448771898, 0.14790319231340754, 0.1471000058279201, 
    0.14629120933860962, 0.14547681732300435, 0.14465692314712519, 
    0.14383168689483958, 0.14300132880628169, 0.1421661168118355, 
    0.14132635694964604, 0.14048237766821822, 0.13963451975917307, 
    0.13878313074013948, 0.13792855492902778, 0.13707112719640044, 
    0.1362111655077852, 0.13534896747909267, 0.13448480590838718, 
    0.13361892545548182, 0.13275154360885352, 0.13188285342929065, 
    0.13101303188198773, 0.13014225018378028, 0.12927068374626846, 
    0.12839852458502346, 0.12752599285955182, 0.12665334885712709, 
    0.1257808994992568, 0.12490900742971704, 0.12403808837317438, 
    0.12316861090204652, 0.12230109574840502, 0.12143610707743059, 
    0.12057425193331511, 0.11971617153739915, 0.11886253153336142, 
    0.11801401669507326, 0.11717132758844617, 0.11633517209988051, 
    0.11550626154544158, 0.11468529961677965, 0.11387297952446301, 
    0.11306997653413095, 0.1122769414831349, 0.11149449674015668, 
    0.11072322615812404, 0.10996367399473461, 0.10921633336476143, 
    0.10848163615326184, 0.10775994838531615, 0.10705155916821374, 
    0.10635667476999956, 0.10567540977773043, 0.10500778760541264, 
    0.10435373611669843, 0.10371309392092928, 0.10308561703888959, 
    0.10247098847781277, 0.10186883182878927, 0.10127872372544071, 
    0.10070020856310577, 0.10013281092061056, 0.099576045719515005, 
    0.099029427993514677, 0.098492483916557336, 0.097964755033725703, 
    0.097445804808339323, 0.096935220684160564, 0.096432617830323378, 
    0.095937636495771944, 0.095449939029397329, 0.094969208356935675, 
    0.094495146740109059, 0.094027474239702813, 0.093565935518785268, 
    0.093110295858118489, 0.092660349646021462, 0.092215916455395744, 
    0.09177684613780368, 0.091343012578765634, 0.090914311208301499, 
    0.090490649516337535, 0.090071937895469315, 0.089658083123763346, 
    0.089248980601777397, 0.088844506001607718, 0.088444515442714408, 
    0.088048847199212243, 0.087657322349928832, 0.087269758612118692, 
    0.086885971875431248, 0.086505793776210663, 0.086129075995252213, 
    0.085755695629038842, 0.085385559228624508, 0.085018600911801107, 
    0.084654782869965112, 0.084294087634919371, 0.083936517560866092, 
    0.083582097051202786, 0.083230870544961519, 0.082882904282432696, 
    0.082538281141879444, 0.08219709240092718, 0.081859428418258801, 
    0.081525366551175815, 0.081194961664016421, 0.080868234221633722, 
    0.080545162051930394, 0.080225670360778725, 0.079909632297094357, 
    0.079596859014139626, 0.079287102354283753, 0.078980051770431478, 
    0.078675340037831831, 0.078372548870357217, 0.078071215983010242, 
    0.077770841956579226, 0.077470901691534963, 0.077170848460707944, 
    0.07687012417726706, 0.076568163711423318, 0.076264404316952472, 
    0.075958300915570445, 0.075649331928483776, 0.0753370137035278, 
    0.075020905710671257, 0.074700620184010177, 0.074375814090708592, 
    0.074046187139276257, 0.073711471459867464, 0.073371420339948784, 
    0.073025802119889599, 0.072674392521275319, 0.072316969703169157, 
    0.071953312301965694, 0.071583200532605182, 0.071206424372037752, 
    0.070822798722704278, 0.070432177310497432, 0.070034465325250359, 
    0.069629633697591647, 0.069217723804705339, 0.068798853001307433, 
    0.068373213750531847, 0.067941070048721533, 0.067502755183712654, 
    0.067058664390572856, 0.066609246653220572, 0.066155001153845261, 
    0.065696471477369192, 0.065234237656392871, 0.064768910195025745, 
    0.064301131994332392, 0.063831569907167138, 0.063360919063358556, 
    0.062889895797414358, 0.06241923884255654, 0.061949704764105419, 
    0.061482060927080584, 0.061017072656996241, 0.060555486019412415, 
    0.060098013584600665, 0.059645317400124014, 0.059197998694867124, 
    0.058756585331228475, 0.05832152860641112, 0.057893194880396952, 
    0.057471860348129358, 0.057057708371174076, 0.056650827675955528, 
    0.056251212423295706, 0.055858769149564724, 0.055473325386893757, 
    0.055094645870430441, 0.054722449027312305, 0.054356418296871475, 
    0.053996212813891303, 0.053641474559224737, 0.053291829068000444, 
    0.052946888501436647, 0.052606257073010344, 0.052269535086733203, 
    0.051936331698367789, 0.051606277448351563, 0.051279037640989664, 
    0.050954329530970441, 0.050631932310851446, 0.050311695502556521, 
    0.049993543746637961, 0.049677472789695941, 0.049363544919236529, 
    0.049051879845489005, 0.048742642119403309, 0.04843602916155635, 
    0.048132257545603227, 0.047831556864189807, 0.04753416275729401, 
    0.047240314109370365, 0.04695025423499774, 0.046664228970509335, 
    0.046382484509402029, 0.046105270335701935, 0.045832831814932605, 
    0.045565409047152165, 0.04530323374898429, 0.045046528526675782, 
    0.044795504462650799, 0.04455036147823789, 0.044311287445619359, 
    0.044078458698190486, 0.043852032421997582, 0.043632145913778085, 
    0.043418904950177563, 0.043212381730365075, 0.043012608741333384, 
    0.042819576020785115, 0.04263323291414383, 0.042453494427177295, 
    0.042280250747954468, 0.042113377434369534, 0.041952748223656328, 
    0.041798247869044985, 0.041649782166991091, 0.041507286888974607, 
    0.041370734638247419, 0.041240137580041185, 0.041115548482467387, 
    0.040997058502126787, 0.040884792011784361, 0.040778901147602055, 
    0.040679556907963432, 0.040586943565326002, 0.040501245775255726, 
    0.040422643966005575, 0.040351303490238209, 0.040287369865686158, 
    0.040230962093780208, 0.040182169266097918, 0.040141050052058119, 
    0.040107632400380441, 0.040081909754501384, 0.04006384183290216, 
    0.040053354417278433, 0.040050341864760974, 0.040054660884186875, 
    0.040066131573121694, 0.040084528704051874, 0.040109582500242394, 
    0.040140975682192194, 0.040178343131122077, 0.04022128130231329, 
    0.040269358943258407, 0.040322132448941797, 0.04037915957340428, 
    0.040440010035022143, 0.040504273411984718, 0.040571560649950704, 
    0.040641508014996441, 0.040713774287147481, 0.040788037013737025, 
    0.040863986369809147, 0.04094131924164035, 0.041019734219824987, 
    0.041098924851151367, 0.041178576458343795, 0.041258361731579693, 
    0.041337936632530263, 0.041416942197604958, 0.041495000408856404, 
    0.04157171355290426, 0.041646661894502661, 0.041719400670142529, 
    0.04178945894900208, 0.041856333529378599, 0.041919490313490036, 
    0.041978365316800589, 0.042032366018626414, 0.042080878091062028, 
    0.042123269940383609, 0.04215890078666959, 0.042187127032970242, 
    0.042207311502337093, 0.042218834299569553, 0.042221104790911124, 
    0.042213572300761323, 0.042195738784944918, 0.042167170141881427, 
    0.042127504390596773, 0.042076459661130217, 0.04201384266735355, 
    0.041939559124389535, 0.041853614739894809, 0.041756124755153758, 
    0.041647310084681227, 0.041527491432092813, 0.04139707880568147, 
    0.04125655682331008, 0.041106466237917381, 0.040947388074009529, 
    0.040779925980168115, 0.040604696273524768, 0.040422318711138314, 
    0.040233414823055258, 0.040038599452847712, 0.039838474416363477, 
    0.039633623801208752, 0.039424603580749701, 0.039211933048254988, 
    0.038996088527252004, 0.0387774956158905, 0.038556522450299772, 
    0.038333482423921705, 0.038108626269532458, 0.037882144092074702, 
    0.037654163359282899, 0.037424749515747702, 0.037193906075230584, 
    0.036961578973853236, 0.036727660633663756, 0.036491995167497744, 
    0.036254383272363862, 0.036014594553918006, 0.035772378812498958, 
    0.035527474765892311, 0.03527962778310257, 0.035028600777351239, 
    0.034774191681485316, 0.034516246877107533, 0.034254671817295856, 
    0.033989445802372509, 0.033720628169053156, 0.033448364017703146, 
    0.033172884166104415, 0.032894502128203683, 0.032613610362365202, 
    0.03233066909624592, 0.032046201347967096, 0.031760780892326118, 
    0.031475021263433975, 0.031189567161476653, 0.030905083642544431, 
    0.030622246358366211, 0.030341728627111608, 0.030064190934133608, 
    0.029790273226389719, 0.029520585565422058, 0.029255707780618909, 
    0.028996180437305428, 0.028742505161612197, 0.028495145548814702, 
    0.028254528749896979, 0.028021048903807928, 0.027795070842598558, 
    0.027576930196886198, 0.027366931564613218, 0.027165347873221935, 
    0.026972416153183944, 0.026788341018296493, 0.026613292203853733, 
    0.026447407920936909, 0.02629079642231966, 0.026143542168712817, 
    0.026005705886393986, 0.02587732689977245, 0.025758424777639066, 
    0.025648998540323115, 0.025549025928856078, 0.025458464816168206, 
    0.025377247131122535, 0.025305276547164881, 0.025242427159836996, 
    0.025188539831482847, 0.025143419421260187, 0.025106836737272271, 
    0.025078528350437231, 0.025058203331536556, 0.025045546667435071, 
    0.025040230027056409, 0.025041917799074921, 0.025050271005458563, 
    0.025064953225128288, 0.025085631487748533, 0.025111981223208683, 
    0.025143684459173102, 0.025180431796000054, 0.025221926668491802, 
    0.025267885354968253, 0.025318039080542993, 0.025372135603834271, 
    0.025429936024826429, 0.025491217262762645, 0.025555772419184438, 
    0.025623411118305035, 0.025693960400260018, 0.025767268862161481, 
    0.025843209743083632, 0.02592168566152139, 0.026002632429413745, 
    0.026086017056326322, 0.026171837553304565, 0.026260117177406714, 
    0.026350895679968907, 0.026444216255458137, 0.02654011690865726, 
    0.026638620161815955, 0.026739727660429508, 0.02684341547996601, 
    0.026949636307928276, 0.027058318417250097, 0.027169374020855529, 
    0.027282699953646537, 0.02739818336259725, 0.027515700335988193, 
    0.027635123479635929, 0.027756322115952858, 0.027879169837133393, 
    0.028003544372246156, 0.028129332172714596, 0.028256431878704805, 
    0.028384758752622034, 0.02851425240093931, 0.028644879356483108, 
    0.02877663842037112, 0.028909557418443262, 0.029043691933642445, 
    0.029179111416977908, 0.029315894049955788, 0.029454111122386679, 
    0.029593822159638617, 0.029735075981010037, 0.029877916092289073, 
    0.03002239344280936, 0.030168570459377826, 0.030316524147042025, 
    0.030466341848275031, 0.03061811061574812, 0.030771904625969678, 
    0.03092777048638734, 0.031085723282061582, 0.031245742002816285, 
    0.031407767873825494, 0.031571705689526129, 0.031737424685788357, 
    0.031904764655507852, 0.032073537644823472, 0.03224353852769829, 
    0.032414548269454856, 0.03258634013146712, 0.032758681780205898, 
    0.032931336523136387, 0.033104059969962324, 0.033276598734164921, 
    0.033448681974604523, 0.033620020476725437, 0.033790297364439378, 
    0.033959165715791766, 0.034126243076846641, 0.034291109917544013, 
    0.034453308690390261, 0.034612341693405144, 0.034767675300543449, 
    0.034918741597162802, 0.035064940963558361, 0.035205650558762326, 
    0.035340229923054439, 0.035468031329915252, 0.035588409939002863, 
    0.035700732817764591, 0.035804396094200976, 0.035898836867833607, 
    0.035983548006882436, 0.036058090810861351, 0.036122101906989057, 
    0.036175299248439707, 0.036217483959574373, 0.036248540795748678, 
    0.036268432887776786, 0.036277200708140785, 0.036274957047256903, 
    0.036261884787337752, 0.036238237920294986, 0.036204335517782273, 
    0.036160562425784325, 0.036107364018933032, 0.036045246431344637, 
    0.035974768370528133, 0.03589653486546894, 0.035811189494950539, 
    0.035719405153506634, 0.035621870712547458, 0.03551927510156451, 
    0.035412294690672821, 0.035301577237765766, 0.035187727565948242, 
    0.035071304343673865, 0.034952814922957258, 0.034832714900111229, 
    0.034711409755054053, 0.034589260148431437, 0.034466582789413752, 
    0.034343649051428254, 0.034220688992035717, 0.03409789156734952, 
    0.033975405451020575, 0.033853337567680664, 0.033731750561879714, 
    0.033610664570496586, 0.03349004972662302, 0.033369832840769796, 
    0.033249893465572965, 0.033130062217307008, 0.033010122382298945, 
    0.032889816564636742, 0.032768849938251063, 0.032646893667952204, 
    0.032523592434591658, 0.032398565161174384, 0.032271415767825801, 
    0.032141734029767582, 0.032009110529172338, 0.031873142927473452, 
    0.031733446510900064, 0.031589665600459858, 0.031441483559932822, 
    0.031288634531765946, 0.031130910766878673, 0.030968171195624401, 
    0.030800347878574556, 0.030627449062731526, 0.030449560541896577, 
    0.030266845343074496, 0.03007953994656315, 0.02988794807568397, 
    0.029692429104007517, 0.029493389811220436, 0.029291272898841963, 
    0.029086546770524135, 0.028879696007910769, 0.028671218465927847, 
    0.02846161608821253, 0.02825138542787492, 0.028041014866677677, 
    0.027830970207734892, 0.02762169172395627, 0.027413582069224712, 
    0.027207005414862904, 0.027002279241890345, 0.026799673222952007, 
    0.026599408948150847, 0.026401658565269298, 0.026206541353863778, 
    0.026014128473861701, 0.025824438796249724, 0.025637442683972625, 
    0.025453057848250943, 0.025271155057392365, 0.025091556422726022, 
    0.024914044651407286, 0.02473835727382, 0.024564191912437767, 
    0.024391207480635623, 0.024219024156473035, 0.024047225830518326, 
    0.023875360181442616, 0.023702942848513282, 0.023529460561426546, 
    0.023354382310531031, 0.023177164173984671, 0.022997257920568535, 
    0.022814120787573288, 0.022627225787447358, 0.022436071403139177, 
    0.02224019250535671, 0.022039171736397609, 0.021832646559197373, 
    0.021620324941821027, 0.021401996457156909, 0.02117754671507047, 
    0.020946975138292308, 0.0207104022945232, 0.020468082786845438, 
    0.020220410510335653, 0.019967919088456722, 0.019711273175023369, 
    0.019451263700706774, 0.019188788177663799, 0.018924834400686597, 
    0.018660459837774382, 0.018396764446979439, 0.018134868743304354, 
    0.017875888868818916, 0.01762091531050761, 0.01737099462242625, 
    0.017127110387403756, 0.016890167284574445, 0.016660979012912885, 
    0.016440257424153941, 0.016228602827753871, 0.016026495602851142, 
    0.015834290767895463, 0.015652212285469102, 0.015480352227416913, 
    0.015318670065727224, 0.015166998253926284, 0.015025053340575658, 
    0.014892445408294099, 0.014768692715999418, 0.014653237024684958, 
    0.014545456270888196, 0.014444682021048635, 0.014350209260154933, 
    0.014261311086142299, 0.014177249747026562, 0.014097290661210094, 
    0.014020710524250486, 0.013946815640370121, 0.01387494911748508, 
    0.013804507625382602, 0.013734950136098774, 0.013665808797900653, 
    0.013596695366100696, 0.013527307463705495, 0.013457431653618002, 
    0.01338694529348995, 0.013315815788629923, 0.013244093181283331, 
    0.013171906226545413, 0.013099452841794949, 0.013026989350595944, 
    0.012954818286779708, 0.012883274549408212, 0.012812714323229965, 
    0.012743501544730846, 0.012675997321524045, 0.012610555069131153, 
    0.012547516270024978, 0.012487203999655215, 0.012429920565266294, 
    0.012375947944822798, 0.012325551342050493, 0.012278978159017625, 
    0.012236465948390276, 0.012198245642987876, 0.012164547234487396, 
    0.012135605800097668, 0.012111664000403588, 0.012092974732985444, 
    0.012079798537506308, 0.012072400577186599, 0.01207103998310639, 
    0.012075958398626905, 0.012087364613423508, 0.012105425168130428, 
    0.012130253046535658, 0.012161906402765635, 0.012200389473211094, 
    0.012245651530425162, 0.012297596575276376, 0.012356087046278335, 
    0.012420956599958427, 0.012492008195100339, 0.012569024600806037, 
    0.012651773057093942, 0.012740012486783567, 0.012833497943437525, 
    0.012931988483193381, 0.013035242847701387, 0.013143026853808866, 
    0.013255109892861874, 0.013371256142106089, 0.013491221845343867, 
    0.013614748697159293, 0.013741560003083048, 0.013871358988306985, 
    0.0140038337802807, 0.014138656341710092, 0.014275494734334156, 
    0.014414021147524849, 0.0145539171507454, 0.01469488965330535, 
    0.014836675442203223, 0.014979048279070444, 0.015121822508198943, 
    0.015264853385912653, 0.015408034339821268, 0.01555129442536927, 
    0.015694587908839593, 0.015837887786097481, 0.015981176629472592, 
    0.016124428607811409, 0.016267604381944831, 0.016410633286897958, 
    0.016553408220317797, 0.016695776164407278, 0.016837532763765973, 
    0.016978416264693527, 0.017118104082886339, 0.017256215284409619, 
    0.017392315714154415, 0.01752591750860601, 0.017656484286573033, 
    0.017783436883915732, 0.017906161797300441, 0.018024021439949807, 
    0.018136372042457792, 0.018242582032939839, 0.018342051142042005, 
    0.018434231768268569, 0.018518643641444905, 0.018594888548850105, 
    0.018662661425570822, 0.01872175570477827, 0.018772068922398664, 
    0.01881359862672085, 0.018846435010265013, 0.018870754611196999, 
    0.01888681100494569, 0.018894926000774071, 0.018895471057633485, 
    0.01888886761861969, 0.018875575024435657, 0.018856086831086916, 
    0.018830925618079114, 0.018800636959844852, 0.018765786868638015, 
    0.018726952680673398, 0.018684718697487009, 0.01863967604894861, 
    0.018592417507981521, 0.018543540720913122, 0.018493649461121392, 
    0.018443346357552369, 0.01839323659857978, 0.018343917727712853, 
    0.018295971253963296, 0.018249946650400053, 0.018206353194052959, 
    0.018165646645912952, 0.018128222037682856, 0.018094404047542187, 
    0.018064447525730994, 0.018038528173369393, 0.018016747940517896, 
    0.017999130535887725, 0.017985624896100966, 0.017976105419581275, 
    0.017970379987801505, 0.017968191310560502, 0.017969223247595961, 
    0.01797310075385361, 0.017979396295693315, 0.017987634912375743, 
    0.017997292900914015, 0.018007802683630912, 0.018018560105811515, 
    0.01802892785004543, 0.01803824619582519, 0.018045838576864804, 
    0.018051017212246254, 0.018053097057837642, 0.018051405017874906, 
    0.018045289142236833, 0.018034131905567571, 0.0180173668057481, 
    0.017994484719585768, 0.017965048099159116, 0.017928696110745587, 
    0.01788514960134226, 0.017834210735222511, 0.01777575956504775, 
    0.017709747349076911, 0.017636188626895692, 0.017555153647748307, 
    0.01746675459737361, 0.017371139902487353, 0.017268483021570916, 
    0.01715897555607826, 0.017042825481745467, 0.016920252601996734, 
    0.016791486998705349, 0.016656771423099195, 0.016516360028581145, 
    0.016370518872645144, 0.016219519062256032, 0.01606363859992295, 
    0.01590315536702884, 0.015738343435618786, 0.015569471087784781, 
    0.015396798660332627, 0.015220587621349948, 0.015041096293004078, 
    0.014858587635314387, 0.014673326176937044, 0.014485579256234829, 
    0.014295614270669187, 0.014103696517391049, 0.013910078310611496, 
    0.013714988856128216, 0.013518627873107149, 0.013321162511610066, 
    0.013122725756633542, 0.012923424736927888, 0.012723352554464568, 
    0.012522608336764605, 0.012321311702337849, 0.012119622015352662, 
    0.011917741109768317, 0.01171592751417673, 0.011514499945153868, 
    0.011313844320922289, 0.011114411263707982, 0.01091671773500805, 
    0.010721342672606564, 0.010528916488708209, 0.010340111507828886, 
    0.010155626053071271, 0.0099761699187421466, 0.0098024441952784015, 
    0.0096351280378978964, 0.0094748605565137881, 0.0093222257605143181, 
    0.0091777427831666557, 0.0090418546927662335, 0.0089149257769144709, 
    0.0087972429735132009, 0.008689013586880779, 0.0085903775984824439, 
    0.0085014181535643212, 0.0084221739729504769, 0.0083526539899009735, 
    0.0082928524622554733, 0.0082427628027996452, 0.0082023870526348602, 
    0.0081717460504509391, 0.0081508806835322925, 0.0081398459517613743, 
    0.0081387023068746588, 0.0081475063767483293, 0.0081662991892519701, 
    0.008195103081248746, 0.0082339121134022055, 0.0082826892786771293, 
    0.0083413632733931077, 0.0084098242057394322, 0.008487918403858959, 
    0.0085754459738812492, 0.0086721556220632837, 0.0087777489831604039, 
    0.0088918823020882332, 0.0090141699706695663, 0.009144193907354806, 
    0.009281514164390367, 0.0094256756887480392, 0.0095762210078271532, 
    0.0097326937660253236, 0.0098946465648982219, 0.010061643647454925, 
    0.010233259168057559, 0.010409070924660936, 0.010588652129324765, 
    0.010771564155989987, 0.010957350464362962, 0.011145529663001259, 
    0.011335592653352305, 0.011526997869236192, 0.011719178947787054, 
    0.011911546434504757, 0.012103495968139985, 0.01229441865084778, 
    0.012483714543685688, 0.012670804399504767, 0.012855138777603952, 
    0.013036217515434356, 0.013213596931158594, 0.013386902354259825, 
    0.013555836414044047, 0.013720187977741704, 0.013879830070752419, 
    0.014034723022208821, 0.014184904616951594, 0.014330491635706035, 
    0.014471670091465105, 0.014608689178466994, 0.014741855763165956, 
    0.014871522393680914, 0.014998075679811772, 0.015121920722753104, 
    0.015243471036341666, 0.015363130170492692, 0.015481276985615421, 
    0.015598253014470631, 0.015714351292227428, 0.015829809321370562, 
    0.015944810259305876, 0.016059485322215954, 0.016173922946975675, 
    0.016288181775560656, 0.016402297996210513, 0.016516301392920926, 
    0.01663022548725827, 0.01674411454564613, 0.016858026407587032, 
    0.016972033573379636, 0.017086219538290863, 0.017200679340816847, 
    0.017315515023319503, 0.017430825878429167, 0.017546708513472134, 
    0.017663251534948986, 0.017780532666761228, 0.017898621556238913, 
    0.018017576861191858, 0.018137450258409241, 0.018258283400233524, 
    0.018380109656163057, 0.018502948500056102, 0.018626802852623817, 
    0.01875165041430215, 0.018877436518380794, 0.01900406823921762, 
    0.019131413923665238, 0.019259300098455265, 0.019387523616879003, 
    0.019515856275570721, 0.019644057765100854, 0.019771889059737639, 
    0.019899120391303121, 0.020025542776243632, 0.020150968512757442, 
    0.020275228634549999, 0.020398178436824236, 0.020519686627387589, 
    0.02063963743469456, 0.020757931527035992, 0.020874483320575163, 
    0.020989230803077567, 0.02110213648526434, 0.021213190413828572, 
    0.021322419249613509, 0.021429880391066112, 0.021535663191414738, 
    0.021639879953918369, 0.021742660956426144, 0.021844145158027389, 
    0.021944476323746864, 0.022043797830473038, 0.022142249311443672, 
    0.022239966957442462, 0.022337075466344617, 0.022433686988608599, 
    0.022529894710230276, 0.022625769145938029, 0.022721349267748433, 
    0.022816636977043326, 0.022911592313045476, 0.023006121074589003, 
    0.023100068201525305, 0.023193217540520457, 0.023285288160680113, 
    0.023375940198167574, 0.023464784590303264, 0.023551399477292199, 
    0.023635346180500182, 0.0237161871895827, 0.023793505341669803, 
    0.023866919151325963, 0.023936102229282892, 0.024000787656667667, 
    0.024060789404194732, 0.02411600762253497, 0.024166439783217652, 
    0.024212180031635524, 0.024253420087258292, 0.024290443174480668, 
    0.024323613764639426, 0.024353363563054856, 0.024380175230144536, 
    0.024404565683920992, 0.024427078021162917, 0.024448272025248415, 
    0.024468717329468467, 0.024488992181396014, 0.024509682404956181, 
    0.024531381769515644, 0.024554690932432264, 0.024580210505183674, 
    0.024608540373294286, 0.024640269778716636, 0.024675972617905263, 
    0.024716197620751026, 0.024761468717461634, 0.024812288066178693, 
    0.024869131687054825, 0.024932446601408417, 0.025002639081064801, 
    0.025080060443231082, 0.02516498667681347, 0.025257602954917198, 
    0.025357991242826856, 0.02546612418984991, 0.025581857572680132, 
    0.025704931564895981, 0.025834972865802733, 0.025971495961056114, 
    0.026113914766238731, 0.02626154564653687, 0.026413614114357088, 
    0.026569260722011451, 0.02672754666742265, 0.026887460894537606, 
    0.027047917269206405, 0.027207762522220624, 0.027365780582360201, 
    0.02752070109678794, 0.027671213610330012, 0.027815987689660988, 
    0.027953698678421918, 0.028083055942674694, 0.028202830489941915, 
    0.028311887687755624, 0.028409208953865606, 0.028493912318245211, 
    0.028565260063524386, 0.028622662802706339, 0.028665673932828636, 
    0.028693974661820474, 0.028707353909504459, 0.028705691343402995, 
    0.028688937427190239, 0.028657100457408817, 0.02861023093423587, 
    0.028548418560444669, 0.028471781972827237, 0.028380463247748903, 
    0.028274630583796107, 0.028154477617764944, 0.028020229209823055, 
    0.027872143373497374, 0.027710519733092551, 0.027535708997738884, 
    0.027348125953170307, 0.027148254117334309, 0.026936652104657708, 
    0.026713951166273675, 0.026480846408598324, 0.026238080417167877, 
    0.025986419890820851, 0.02572662825745024, 0.025459440874404771, 
    0.025185544590083639, 0.024905561673437594, 0.024620045172792291, 
    0.024329477176208727, 0.024034280609459873, 0.023734825849204607, 
    0.023431446295758811, 0.023124456387203649, 0.022814164630614323, 
    0.022500891352567522, 0.022184965497233325, 0.021866733239044495, 
    0.021546550460372207, 0.021224785134299849, 0.020901810300668965, 
    0.020578002579924582, 0.020253737306958966, 0.019929392491631205, 
    0.019605344270875631, 0.019281963536356694, 0.018959623147824338, 
    0.018638692413557475, 0.018319540769699258, 0.018002536872349706, 
    0.017688046985470246, 0.017376434791105597, 0.017068054874656464, 
    0.01676325635310838, 0.016462374024258614, 0.01616572706865059, 
    0.015873612287269682, 0.01558630138143027, 0.015304045141285635, 
    0.015027079431672695, 0.014755629438596349, 0.014489914390692752, 
    0.014230148381427721, 0.013976550145867061, 0.013729336994608418, 
    0.013488725694776986, 0.013254925902607661, 0.013028141411740773, 
    0.012808571442883535, 0.012596418070747411, 0.012391885664425379, 
    0.01219519287128361, 0.012006576498907573, 0.011826300592533154, 
    0.011654657932865695, 0.011491970040827054, 0.01133858697919384, 
    0.011194877051804471, 0.011061227400260294, 0.01093802383825869, 
    0.010825637630731293, 0.010724418202913337, 0.010634671710821051, 
    0.01055665324317777, 0.010490557635056517, 0.010436507163454503, 
    0.010394551043710724, 0.010364658360293605, 0.01034671944210558, 
    0.010340542553970008, 0.010345855814313458, 0.010362316995457612, 
    0.010389514405048476, 0.010426977624745063, 0.010474188992673434, 
    0.010530592803764227, 0.010595599121370142, 0.010668589377880084, 
    0.010748919590539658, 0.010835917808306455, 0.010928886672527576, 
    0.011027096895884983, 0.011129790595689564, 0.011236187559632861, 
    0.011345489402245704, 0.011456892410643417, 0.011569589974835348, 
    0.01168278400896793, 0.011795692871828864, 0.011907552455045045, 
    0.012017613312584089, 0.01212513804392344, 0.012229396574785828, 
    0.012329665787576228, 0.01242522842880058, 0.012515382950112758, 
    0.012599465486288024, 0.012676870078512471, 0.012747071772756375, 
    0.012809641223064208, 0.012864249260805091, 0.012910667026209058, 
    0.012948759322889206, 0.01297847255392932, 0.012999822815785623, 
    0.013012890542364156, 0.013017809283026292, 0.013014759729025075, 
    0.013003974449165991, 0.0129857333482733, 0.012960361224299916, 
    0.012928233782041304, 0.012889769901183517, 0.012845425717184016, 
    0.012795692944114839, 0.012741081504382018, 0.012682103571208286, 
    0.012619265932297594, 0.012553051303795413, 0.012483911486294319, 
    0.012412251274733372, 0.012338425474963041, 0.012262731239461247, 
    0.012185407769519365, 0.012106634612098086, 0.012026531536630015, 
    0.011945155934877794, 0.011862499679557182, 0.011778484486653428, 
    0.011692954918529183, 0.011605676412153076, 0.011516325201555882, 
    0.011424485332996811, 0.011329640580550556, 0.011231179048875817, 
    0.011128393264843127, 0.011020495665063702, 0.010906637413969297, 
    0.010785928043066223, 0.010657456738893728, 0.010520310451356336, 
    0.01037358413732138, 0.010216395623676666, 0.010047896797038693, 
    0.0098672912109675198, 0.0096738530010007304, 0.0094669528366870277, 
    0.0092460702762590212, 0.009010816088044115, 0.0087609363122207896, 
    0.0084963178598438799, 0.0082169904292887959, 0.0079231352458750664, 
    0.007615086797415193, 0.0072933440664143473, 0.0069585680353991177, 
    0.0066115923384305894, 0.0062534186577982943, 0.005885216676324868, 
    0.0055083058088265377, 0.0051241445458604234, 0.0047343089053767506, 
    0.0043404654397237365, 0.0039443451289936093, 0.0035477218324459852, 
    0.0031523786411201964, 0.0027600739482026449, 0.0023725081431829795, 
    0.0019912944735645216, 0.0016179329018506509, 0.0012537922966775023, 
    0.00090010224268788374, 0.00055794845015001303, 0.00022828203209470678, 
    -8.8086764627550536e-05, -0.00039048877924688905, 
    -0.00067839887428346158, -0.00095143748006610608, -0.0012093591581210565, 
    -0.001452039988864602, -0.0016794618158172123, -0.0018916993602937995, 
    -0.0020889066863719781, -0.0022713094939626763, -0.0024392004850990502, 
    -0.0025929456582774141, -0.002732983945732851, -0.002859822194733669, 
    -0.0029740300054915915, -0.0030762344120865278, -0.0031671068042404037, 
    -0.0032473411044230665, -0.0033176407186942931, -0.0033787055220839343, 
    -0.003431214722993051, -0.0034758121108941541, -0.0035131051869880742, 
    -0.0035436436690931983, -0.003567921685852583, -0.003586369876384366, 
    -0.0035993537756689011, -0.0036071680075996774, -0.0036100503162789996, 
    -0.0036081851288592781, -0.0036017224128224168, -0.0035907866001311526, 
    -0.0035754930922951419, -0.0035559559588768629, -0.0035322867440615181, 
    -0.0035045863351913439, -0.0034729408232464275, -0.0034374042011864033, 
    -0.0033980013068263589, -0.0033547253183351723, -0.0033075385659622181, 
    -0.0032563881897628706, -0.0032012081780826949, -0.0031419410300930319, 
    -0.0030785489138346503, -0.003011025772562782, -0.0029394080371203677, 
    -0.0028637810977577009, -0.0027842872811549343, -0.002701119558328966, 
    -0.002614519354677102, -0.002524757440673387, -0.0024321295048079718, 
    -0.0023369458180802403, -0.0022395150055845754, -0.0021401363125576143, 
    -0.002039090176339073, -0.0019366327325842638, -0.0018329875383960496, 
    -0.0017283460590879225, -0.001622865558949086, -0.0015166699000470471, 
    -0.0014098617095516931, -0.0013025181680212221, -0.0011947101114513517, 
    -0.00108650267013262, -0.00097796315594289303, -0.0008691817669225127, 
    -0.00076026992683884726, -0.00065137062875598897, 
    -0.00054265759061975264, -0.00043431806783901755, 
    -0.00032655501103322237, -0.00021956167772493916, 
    -0.00011350235538952393, -8.4954576665006911e-06, 9.5405516969122254e-05, 
    0.00019822845712169179, 0.00030009122370704112, 0.00040120638944927804, 
    0.00050188452614334501, 0.00060253153244039636, 0.00070364483282967481, 
    0.00080581148362303835, 0.00090968783968626665, 0.0010159956134048347, 
    0.0011254925345854838, 0.0012389643240594199, 0.0013572028297842145, 
    0.0014809849986917585, 0.0016110560034543523, 0.0017481123074477209, 
    0.001892784451363307, 0.0020456138666147001, 0.0022070413153780725, 
    0.0023773963965057414, 0.0025568953841190729, 0.0027456347293587698, 
    0.0029435991325148956, 0.003150642588770112, 0.0033664850185604199, 
    0.0035906977722333505, 0.0038226914567228041, 0.0040617318832601688, 
    0.0043069382130005076, 0.0045573137029959344, 0.0048117722526804562, 
    0.0050691662744545441, 0.0053283009801300789, 0.0055879705653927364, 
    0.0058469677130742886, 0.0061041026337595675, 0.0063582172284754575, 
    0.0066081847201514138, 0.0068529120847402279, 0.0070913418556921284, 
    0.0073224584245901031, 0.0075452869738357013, 0.0077589084786945555, 
    0.0079624541938586313, 0.0081551227044117415, 0.0083361777492500164, 
    0.0085049635629953994, 0.0086609067780078347, 0.0088035214433422986, 
    0.0089324110319454648, 0.0090472823354375322, 0.0091479493789534978, 
    0.0092343481354705548, 0.0093065483847571562, 0.0093647704991403173, 
    0.0094093893852473312, 0.0094409395892176493, 0.0094601133219103378, 
    0.0094677478460713678, 0.009464817067130666, 0.0094524066182334263, 
    0.0094316732944216847, 0.0094037980081848587, 0.0093699323069823971, 
    0.0093311527764767237, 0.0092884406581959216, 0.0092426890146019101, 
    0.00919471541195091, 0.0091452873148695438, 0.0090951210125559279, 
    0.0090448993197830389, 0.0089952641616241977, 0.0089468333057915253, 
    0.0089002085899301496, 0.0088559832367164464, 0.0088147434973918984, 
    0.0087770716189874923, 0.0087435478007687525, 0.0087147428727942181, 
    0.0086912258092187011, 0.0086735699155769935, 0.0086623518549036986, 
    0.0086581611841927524, 0.0086615839399540526, 0.0086731903349429509, 
    0.0086935165701693025, 0.0087230353296750742, 0.0087621458383284785, 
    0.0088111516775651478, 0.0088702581690187337, 0.0089395717379019291, 
    0.0090191091731410596, 0.0091088023945680632, 0.0092085050949792385, 
    0.0093179853639144099, 0.009436923830753596, 0.0095649154813258093, 
    0.0097014648948624133, 0.0098459921690120852, 0.0099978464003576666, 
    0.010156343634566276, 0.010320807024856719, 0.010490601837583364, 
    0.01066517638226426, 0.010844086031197351, 0.01102701747209341, 
    0.011213791589621321, 0.011404358668538259, 0.011598802889496308, 
    0.011797309264385353, 0.012000148109596147, 0.01220763998320795, 
    0.012420139489302876, 0.012638014042708926, 0.012861620625762807, 
    0.013091310333798982, 0.013327417003790948, 0.013570254425016512, 
    0.013820131887840419, 0.014077349373615456, 0.014342207279135384, 
    0.014615022203298978, 0.014896133560533395, 0.015185900767707507, 
    0.015484704069890561, 0.015792909984412819, 0.016110855941680435, 
    0.016438801928055646, 0.016776900040449634, 0.017125156787995258, 
    0.017483407971488792, 0.017851304094480408, 0.01822831305133055, 
    0.018613722437767672, 0.019006650031471364, 0.019406085388207428, 
    0.019810905446535618, 0.020219923285481122, 0.020631911536714773, 
    0.021045645373534143, 0.021459926426245442, 0.021873615263414952, 
    0.022285649320941237, 0.022695054101509536, 0.023100951706291572, 
    0.023502551962085512, 0.023899158786625366, 0.024290162359676931, 
    0.024675022203451545, 0.025053251536909345, 0.025424401783876716, 
    0.0257880480211139, 0.02614377682463884, 0.026491189143074311, 
    0.02682988933687043, 0.027159484611125811, 0.027479581697677558, 
    0.027789779013510946, 0.02808967062007792, 0.02837883069672437, 
    0.028656810743542732, 0.028923132647252939, 0.029177290416640821, 
    0.029418745696382805, 0.029646925090634393, 0.029861215764110077, 
    0.030060969701560004, 0.030245516715483152, 0.030414153316731907, 
    0.030566161958937882, 0.030700803996208281, 0.030817348170338613, 
    0.030915061069860611, 0.030993237877167509, 0.031051211439276891, 
    0.031088372172640672, 0.03110419443597269, 0.031098264831605014, 
    0.031070298830356991, 0.031020182413171418, 0.030947978934820021, 
    0.030853943689753263, 0.03073853187541643, 0.030602385438872566, 
    0.030446331575990741, 0.030271378331152614, 0.030078696827690678, 
    0.029869614452396647, 0.02964560029724041, 0.029408255169811073, 
    0.029159305972120655, 0.028900584182336413, 0.028634008351628805, 
    0.028361557318281851, 0.028085250638867448, 0.027807101533063844, 
    0.027529090447369897, 0.027253119931599155, 0.026980984535496952, 
    0.026714348136264516, 0.026454730993166493, 0.026203512406365665, 
    0.025961920970555719, 0.025731025002605365, 0.025511725843668408, 
    0.025304712990312742, 0.025110449439510216, 0.024929152964751622, 
    0.024760770873455067, 0.024605019968830862, 0.024461410977575721, 
    0.024329290722210059, 0.024207897014448875, 0.024096402761809695, 
    0.023993963582490785, 0.02389976313883042, 0.023813023607651095, 
    0.023733030423601257, 0.023659150127245402, 0.023590829927705972, 
    0.023527618592309965, 0.023469163867640697, 0.023415225829491609, 
    0.02336568954213954, 0.023320562551843019, 0.023279978955802427, 
    0.023244210980426349, 0.0232136617019933, 0.023188847535798036, 
    0.023170374215303404, 0.023158898511364587, 0.023155085976852091, 
    0.023159568199623632, 0.023172929462693458, 0.023195670623988286, 
    0.023228235960559639, 0.023270990903734967, 0.023324246137413834, 
    0.023388264395728296, 0.023463269688186482, 0.023549434210271645, 
    0.023646870021081876, 0.02375563406211461, 0.023875716850431675, 
    0.024007031897469576, 0.0241494202241593, 0.024302636802320487, 
    0.024466356569021332, 0.024640176450736202, 0.024823609075811916, 
    0.025016110329512318, 0.02521709099099393, 0.025425931167224202, 
    0.025642017539636824, 0.02586477080187851, 0.026093665985320515, 
    0.026328275021179674, 0.026568272815864144, 0.026813440458652808, 
    0.027063665597674803, 0.027318915266299371, 0.027579239683727552, 
    0.027844752801986856, 0.028115625265708807, 0.028392087921548084, 
    0.028674422956172604, 0.028963001213111954, 0.029258280088942077, 
    0.029560831917739273, 0.029871360906252947, 0.030190700913365731, 
    0.030519834192177634, 0.030859862994051534, 0.031211992381440831, 
    0.031577475152112212, 0.031957560734961143, 0.032353425106925689, 
    0.032766112042937431, 0.033196490461721753, 0.03364519281060991, 
    0.034112580896610879, 0.03459869798897653, 0.035103263733094685, 
    0.035625694229848091, 0.036165127373317715, 0.036720456074251694, 
    0.037290381285705311, 0.037873428958363403, 0.038467974992569612, 
    0.0390722610507978, 0.039684409481184943, 0.040302428484743795, 
    0.040924242025541756, 0.041547730441937283, 0.042170749017156901, 
    0.04279117698172924, 0.043406935317065701, 0.044016010906501403, 
    0.044616461513454254, 0.045206414138958047, 0.045784057343866244, 
    0.046347644750310078, 0.046895469081128044, 0.04742587251314774, 
    0.047937230946172242, 0.048427954772014885, 0.048896506648764666, 
    0.049341396228677156, 0.049761195558575173, 0.050154566260271351, 
    0.050520239231950065, 0.050857040567638429, 0.051163880978003125, 
    0.051439754065662667, 0.051683709380446502, 0.051894837187303526, 
    0.052072242394117396, 0.052215028857488036, 0.052322284793148793, 
    0.052393090080155087, 0.05242654817433904, 0.052421829659640755, 
    0.05237826527607925, 0.052295377768547119, 0.052172940724968322, 
    0.052010971819499263, 0.051809729771033319, 0.051569617180427296, 
    0.05129113408383254, 0.050974788226642441, 0.050621027305044974, 
    0.050230204549505345, 0.049802593416682701, 0.049338437864016961, 
    0.048837990184838455, 0.0483015545298097, 0.047729525765062467, 
    0.047122405540258198, 0.046480835439971738, 0.045805623265678767, 
    0.045097760014395631, 0.044358485032707402, 0.043589252689592337, 
    0.042791785694045209, 0.041968020791068331, 0.04112008607659836, 
    0.040250237587302978, 0.039360783599748386, 0.038454051399191835, 
    0.037532300198669689, 0.036597673609869888, 0.035652163756020989, 
    0.034697578404437011, 0.033735504650552015, 0.032767306445474563, 
    0.031794126048756241, 0.030816888580997209, 0.029836342948040308, 
    0.028853112651064057, 0.027867846694809382, 0.026881274815675153, 
    0.02589430695213174, 0.024908020676014123, 0.02392369881331859, 
    0.022942750462818504, 0.021966786523840463, 0.020997557190089226, 
    0.020037034457191266, 0.019087475542910771, 0.018151480877103582, 
    0.017232057165977716, 0.016332629834188275, 0.015457036608445225, 
    0.014609505642927529, 0.013794508995000201, 0.013016677002417147, 
    0.012280642182893615, 0.011590924429284145, 0.010951806890043495, 
    0.010367278147884219, 0.0098409759491659594, 0.0093761962119823447, 
    0.0089758982178381221, 0.0086426891967191811, 0.0083788571448272821, 
    0.0081864219594741643, 0.0080671358297155545, 0.0080225694550819012, 
    0.0080541923209773957, 0.0081634086432880917, 0.008351665535267741, 
    0.0086204053243296164, 0.0089710565797380057, 0.0094048998319381863, 
    0.0099229682928079835, 0.01052593832739156, 0.01121400177216922, 
    0.011986796774434455, 0.012843358963814847, 0.013782105439678279, 
    0.014800870563440285, 0.015897000274756226, 0.017067449897479225, 
    0.01830901011022892, 0.019618404496758311, 0.02099248265415115, 
    0.022428308146232184, 0.023923346298538296, 0.025475443906757392, 
    0.027082821786497489, 0.028744033167403846, 0.030457743084217101, 
    0.032222659120302755, 0.034037348126266735, 0.035900099812994704, 
    0.037808716383466404, 0.039760289253882357, 0.041751053903483881, 
    0.043776347791465241, 0.045830508205847283, 0.047907016378126124, 
    0.04999859973715283, 0.052097455957971599, 0.054195625839272323, 
    0.056285207534939832, 0.058358564607504111, 0.060408512575119956, 
    0.062428331841567312, 0.064412080875784539, 0.066354561169631232, 
    0.068251533251144969, 0.070099575538042788, 0.071896239301113843, 
    0.073639611852444123, 0.075328217699625749, 0.076960708433663746, 
    0.078535496316745224, 0.080050475320087106, 0.081502758609768286, 
    0.082888494060690016, 0.084202605966384209, 0.085438819252028633, 
    0.086589723511505415, 0.087647305388950589, 0.088602986501719772, 
    0.089448249158531015, 0.090174806037478072, 0.090775124659376996, 
    0.091242942613303235, 0.09157393561092915,
  // Fqt-F(2, 0-1999)
    1, 0.99898754410228308, 0.99596355310686779, 0.99096810864983109, 
    0.98406678892612764, 0.97534853284593592, 0.96492285275606471, 
    0.95291656630811217, 0.93947023093701709, 0.92473445935892484, 
    0.90886627814567933, 0.89202566456363963, 0.87437237283660962, 
    0.85606311031145998, 0.8372491202454645, 0.81807418126856601, 
    0.79867301632370935, 0.77917010572151624, 0.75967886721729838, 
    0.74030116311457239, 0.72112711188273937, 0.70223515341032938, 
    0.68369233445082178, 0.66555477149557807, 0.64786825109118784, 
    0.6306689324897552, 0.61398411520737139, 0.59783304533206938, 
    0.58222772303552361, 0.56717372274844069, 0.55267099764530647, 
    0.53871465214121783, 0.52529568613041588, 0.51240167901614164, 
    0.50001741966837754, 0.48812547916950627, 0.47670671966369815, 
    0.46574075600216625, 0.45520636468801384, 0.44508185200067457, 
    0.43534538060034406, 0.42597527195185275, 0.41695025904437855, 
    0.40824971734620075, 0.39985384479563713, 0.39174380634230721, 
    0.38390183906401815, 0.3763113185843574, 0.36895679597485914, 
    0.36182400871148163, 0.35489987497774905, 0.34817246147295633, 
    0.34163094608407973, 0.33526556758115877, 0.32906755712176966, 
    0.32302906601313147, 0.31714308134153379, 0.3114033341957218, 
    0.30580420838747246, 0.30034064485340095, 0.29500805821629472, 
    0.28980225475665, 0.28471936552010002, 0.27975579404682283, 
    0.27490816493827896, 0.27017329742578389, 0.26554817885671672, 
    0.26102994476639552, 0.25661586523565322, 0.25230332302193198, 
    0.24808980088232516, 0.24397285451505352, 0.23995009767062739, 
    0.23601916907978987, 0.2321777117867071, 0.22842334578389581, 
    0.22475364257513603, 0.22116610911729756, 0.21765816765020779, 
    0.21422715168647988, 0.2108703007029569, 0.2075847637856594, 
    0.20436761632461023, 0.20121587417742182, 0.19812651612943086, 
    0.19509651315360782, 0.19212285142953539, 0.18920256683134329, 
    0.18633277494425965, 0.18351070466176039, 0.18073373329512565, 
    0.17799941097828581, 0.1753054925982081, 0.17264995566112445, 
    0.17003102506768739, 0.16744718567210939, 0.16489719906235348, 
    0.16238011693481669, 0.15989528277256201, 0.15744232782347095, 
    0.15502116440435842, 0.15263197708379669, 0.15027520235182665, 
    0.14795151064665721, 0.14566178283896689, 0.14340708247239825, 
    0.14118862456583783, 0.13900774090585924, 0.13686584862716838, 
    0.13476441074777834, 0.13270490027458623, 0.13068875751361814, 
    0.12871735743344395, 0.12679197205866494, 0.12491374416221467, 
    0.12308365904447752, 0.12130252753246996, 0.11957097064781863, 
    0.11788942099700057, 0.11625811654715203, 0.11467711319816984, 
    0.11314629018691578, 0.11166536598510252, 0.11023391443402621, 
    0.10885137048187853, 0.10751704482076045, 0.10623012576128112, 
    0.10498968609024033, 0.10379468323845729, 0.10264396078991037, 
    0.10153624129696821, 0.10047012925499874, 0.099444106543284463, 
    0.098456535792735389, 0.097505661187218332, 0.096589619530935117, 
    0.095706452495946767, 0.094854123246043073, 0.094030533685001097, 
    0.093233553577074038, 0.092461034227438885, 0.0917108375733139, 
    0.090980855314391471, 0.090269033734004092, 0.089573384789853369, 
    0.088892006686402639, 0.088223094707440053, 0.087564956997796164, 
    0.086916016941165686, 0.086274824216452078, 0.085640061351381747, 
    0.085010546030089063, 0.084385238118701841, 0.083763233221462008, 
    0.083143768072920815, 0.082526208755128602, 0.081910043805249175, 
    0.081294861152220052, 0.080680329176132104, 0.080066163619848377, 
    0.079452105035694165, 0.078837881254584297, 0.078223188082442774, 
    0.077607670310094204, 0.076990922157286992, 0.076372488789155271, 
    0.075751888447272292, 0.075128638673526857, 0.074502291016301903, 
    0.073872471447598717, 0.073238923883291507, 0.072601544439282184, 
    0.071960406696324697, 0.071315773364797067, 0.070668090319796248, 
    0.0700179721769396, 0.069366176900647447, 0.068713574403311925, 
    0.068061115953228682, 0.067409797778998665, 0.066760622899943112, 
    0.06611456861519216, 0.065472558847062906, 0.064835438400031031, 
    0.064203962385438879, 0.063578792191474512, 0.062960495039266803, 
    0.062349549197323204, 0.061746354385249849, 0.061151241428799047, 
    0.060564485250401701, 0.05998631500879275, 0.059416926824691602, 
    0.05885649015450263, 0.05830515748345666, 0.057763068477058192, 
    0.057230353662035896, 0.056707133865853306, 0.056193520410118963, 
    0.055689617506081653, 0.055195516241022952, 0.05471129661621553, 
    0.054237025123842625, 0.05377275475452175, 0.053318521482181351, 
    0.052874346471905247, 0.05244023817834402, 0.052016187582724284, 
    0.051602180019482226, 0.051198190573708426, 0.050804195733254398, 
    0.0504201768163276, 0.05004612501020058, 0.049682040652164229, 
    0.049327931892894326, 0.048983810553623899, 0.048649688802276929, 
    0.048325572933612407, 0.04801146166423835, 0.047707338952367208, 
    0.047413170976183625, 0.047128895958043704, 0.046854421778716814, 
    0.046589608602845674, 0.04633426360388232, 0.046088126482847783, 
    0.045850858565878977, 0.045622032221143832, 0.045401122799175631, 
    0.045187506998649367, 0.044980463911111324, 0.044779177387711006, 
    0.044582745692494818, 0.044390190411945744, 0.044200469864021104, 
    0.044012488724974951, 0.043825119006712279, 0.043637207499760869, 
    0.043447599663472905, 0.043255152718564664, 0.043058753407874031, 
    0.042857336155040886, 0.042649900895861438, 0.042435521843785934, 
    0.042213359281368268, 0.041982664045061284, 0.041742783438212923, 
    0.041493162462391493, 0.04123334586738104, 0.040962976761813701, 
    0.040681789437749388, 0.040389607262812786, 0.040086339195655143, 
    0.039771971788129808, 0.039446567751060861, 0.039110261329450828, 
    0.038763257746988591, 0.038405837167348571, 0.03803835768212762, 
    0.037661258959332117, 0.037275065722108841, 0.036880382188890962, 
    0.036477886129584282, 0.036068312697943757, 0.035652435277675025, 
    0.035231044104577974, 0.034804922306613667, 0.034374819913052287, 
    0.033941435482172912, 0.033505398355654095, 0.033067253107529851, 
    0.032627440800018497, 0.032186292326538808, 0.031744015969691924, 
    0.031300689671206604, 0.030856262484234731, 0.030410562375393736, 
    0.029963308182625298, 0.029514134604651535, 0.029062620180006479, 
    0.028608324843044149, 0.02815082669910323, 0.027689766991162403, 
    0.027224886520848986, 0.026756064311389993, 0.026283342319645804, 
    0.025806945388259169, 0.025327286973665916, 0.024844963897235818, 
    0.024360751884632048, 0.023875582572218963, 0.023390516120731519, 
    0.022906718585341233, 0.022425435026318299, 0.021947964623517509, 
    0.021475633312661922, 0.021009764726082514, 0.020551659767770212, 
    0.020102567789292081, 0.019663663257518511, 0.019236021372312111, 
    0.018820594023421865, 0.018418190596829188, 0.018029461956498193, 
    0.017654879239972335, 0.017294732569518304, 0.016949121845687493, 
    0.016617958121169084, 0.016300962768387099, 0.015997678661357841, 
    0.015707484514899006, 0.01542962989271573, 0.015163273382324366, 
    0.014907528686729114, 0.014661507655310095, 0.014424361614312941, 
    0.014195315628914931, 0.013973689633973914, 0.013758911335916066, 
    0.013550525443929104, 0.013348196119189746, 0.013151698811474006, 
    0.01296091817929257, 0.012775833950203904, 0.012596510184144132, 
    0.012423079405594303, 0.012255727601164156, 0.01209467860498626, 
    0.011940179356588016, 0.011792485634706648, 0.011651855994868652, 
    0.01151853991302464, 0.011392774903278625, 0.011274776234643851, 
    0.011164736491640834, 0.011062814106717157, 0.010969133371991228, 
    0.010883771841786299, 0.010806754999361205, 0.010738049142966043, 
    0.010677556415385279, 0.010625107689956172, 0.010580462779137502, 
    0.010543319035701602, 0.010513312688773393, 0.010490035333663779, 
    0.010473038317289995, 0.010461851774062388, 0.010455992366846058, 
    0.010454972098865206, 0.010458309819749909, 0.010465540247752781, 
    0.010476225957150852, 0.010489962919691412, 0.010506394000878539, 
    0.010525220839845867, 0.01054620995837903, 0.010569200687253366, 
    0.010594105590541712, 0.010620904822939821, 0.010649634842596893, 
    0.010680373189945436, 0.010713219382236891, 0.010748269357285505, 
    0.01078559065878326, 0.010825193780623268, 0.010867010013121682, 
    0.010910859343467741, 0.010956433533456669, 0.011003277803447982, 
    0.011050784605959372, 0.011098193352621159, 0.011144597942388075, 
    0.011188957975600716, 0.011230118941405907, 0.011266834049167548, 
    0.011297791446554125, 0.011321644104245333, 0.011337048277303139, 
    0.01134270271049796, 0.011337384530567401, 0.011319981075256018, 
    0.011289507150262086, 0.011245124836796258, 0.011186140749053303, 
    0.011112002336083305, 0.011022286105562695, 0.010916678322030686, 
    0.010794971697563122, 0.010657058446535358, 0.010502945672153072, 
    0.010332772014277614, 0.010146831151860001, 0.009945587860761199, 
    0.0097296826098977971, 0.0094999317141011841, 0.0092573168844187152, 
    0.0090029749299527055, 0.0087381764337256564, 0.0084643102639685511, 
    0.0081828545468164687, 0.007895350743919392, 0.0076033784063996432, 
    0.0073085290712660289, 0.0070123779452738759, 0.0067164641501826858, 
    0.0064222673796353888, 0.0061311905312165984, 0.005844547503616967, 
    0.0055635585841242894, 0.0052893432130285099, 0.005022924155955742, 
    0.0047652231560111691, 0.0045170638073272172, 0.0042791631211798959, 
    0.0040521244986173478, 0.0038364232395936581, 0.003632391410406124, 
    0.0034402106389713723, 0.0032599000362049674, 0.0030913170203830109, 
    0.0029341630785802131, 0.0027879938088303051, 0.0026522361338869589, 
    0.0025262068119865267, 0.0024091362392591881, 0.0023001928712089088, 
    0.0021985128306169573, 0.0021032273426936474, 0.0020134893460296366, 
    0.001928502576039051, 0.0018475448384871916, 0.0017699833083020438, 
    0.0016952882521037737, 0.0016230360471725324, 0.0015528999783491829, 
    0.0014846377261994864, 0.001418074656436885, 0.0013530883454900228, 
    0.0012895927218347565, 0.0012275284722957137, 0.0011668546880212389, 
    0.0011075473458737372, 0.001049594268235198, 0.00099299722064634215, 
    0.00093777425503309701, 0.00088396371349201382, 0.00083162512794662325, 
    0.00078084574611350665, 0.00073173997654937839, 0.00068444538242976808, 
    0.00063911977770366509, 0.00059593647393045611, 0.00055508068784432111, 
    0.00051675129530449936, 0.00048115742106623598, 0.00044852057618389985, 
    0.00041906216895174376, 0.00039299394473350162, 0.00037050080107851923, 
    0.00035172095405157085, 0.00033672573121727842, 0.0003255061581150583, 
    0.00031796085172546885, 0.00031389202661659811, 0.00031300439195835529, 
    0.00031491404486818828, 0.00031915342307972975, 0.00032518959915513537, 
    0.00033243804367216973, 0.00034028712424975436, 0.00034811783455114781, 
    0.00035533063246112129, 0.00036137211361746824, 0.00036576521438540406, 
    0.0003681348507087337, 0.00036822586217913897, 0.00036591813126223032, 
    0.000361228427947215, 0.00035430559824897403, 0.00034541615013842077, 
    0.0003349228890112286, 0.00032325658191380199, 0.00031088573896324563, 
    0.00029828541952034882, 0.00028590690542113222, 0.00027415260686778909, 
    0.00026335590348553194, 0.00025376650396626103, 0.00024553409888683687, 
    0.00023870462754310798, 0.00023321193205020282, 0.00022888138186622848, 
    0.00022542608334697958, 0.00022244987279141715, 0.00021945275352966155, 
    0.00021584309702196231, 0.00021094640659040538, 0.00020402563529617576, 
    0.00019430448827898838, 0.00018099327927087016, 0.00016330813659715237, 
    0.00014049658187586194, 0.00011185666908468435, 7.6766987918561576e-05, 
    3.4712103212062488e-05, -1.4686678016382054e-05, -7.1639137985197185e-05, 
    -0.00013615943952037182, -0.00020804581649628835, 
    -0.00028687298803965506, -0.00037199913068540003, 
    -0.00046257760924084586, -0.00055758606473812458, 
    -0.00065584287144988232, -0.00075604027868038143, 
    -0.00085676930777668246, -0.00095655319960461535, -0.0010538812351570466, 
    -0.0011472487245905206, -0.0012351965459225195, -0.0013163551845566104, 
    -0.0013894850066647005, -0.0014535122700563587, -0.0015075499571341733, 
    -0.0015509127938780286, -0.001583111706588378, -0.001603845192071209, 
    -0.0016129841537240663, -0.0016105537518610494, -0.0015967271754359945, 
    -0.0015718118954438887, -0.0015362447075035568, -0.0014905846505828583, 
    -0.0014355029268440635, -0.0013717704387844274, -0.0013002464001472434, 
    -0.0012218569183170653, -0.0011375801976793258, -0.0010484295507726736, 
    -0.00095543600063633337, -0.00085963112589124786, 
    -0.00076202769412918802, -0.00066359898814843227, 
    -0.00056525578848799177, -0.00046783008237645171, 
    -0.00037205232216058217, -0.00027853573411425702, 
    -0.00018777201660971903, -0.00010011808484755385, 
    -1.5796327280903058e-05, 6.510282765248332e-05, 0.00014260902470123919, 
    0.00021686172142004116, 0.00028808550570601378, 0.00035657709057875555, 
    0.00042268848067595873, 0.0004868192510334296, 0.00054941001326394025, 
    0.00061094194253048155, 0.00067192749923975306, 0.00073289124598391287, 
    0.00079435264349113051, 0.00085679575879528663, 0.00092064569791160578, 
    0.00098624433450753132, 0.0010538284653790124, 0.0011235093154129629, 
    0.0011952658853338085, 0.0012689348881822025, 0.0013442119987872084, 
    0.0014206524186839958, 0.0014976825461541627, 0.0015746121840331578, 
    0.001650653462871837, 0.0017249431493106509, 0.0017965606660794602, 
    0.0018645528606844272, 0.0019279583224841783, 0.0019858379610780525, 
    0.0020372974138494876, 0.0020815186615927802, 0.0021177861337980238, 
    0.0021455134904723575, 0.0021642598455508763, 0.0021737390053259528, 
    0.0021738188566162589, 0.0021645208456599059, 0.0021460072048282838, 
    0.0021185689692301479, 0.0020826146568670447, 0.0020386582335524535, 
    0.001987304675291316, 0.0019292456693185524, 0.0018652473682273045, 
    0.0017961412340633722, 0.0017228154399366062, 0.0016461985015095888, 
    0.0015672422321852428, 0.0014869014040318901, 0.0014061215792033825, 
    0.0013258185975831148, 0.0012468672740436379, 0.0011700889712295869, 
    0.0010962444997117344, 0.0010260267742867599, 0.00096006598845792615, 
    0.00089893401197822624, 0.00084315745182698401, 0.00079322759410818656, 
    0.00074960786985327416, 0.00071274010921517663, 0.00068304593952617319, 
    0.00066092231402651517, 0.00064674351245196289, 0.00064084996559334538, 
    0.00064354684444317386, 0.00065509756152980453, 0.00067571593603359278, 
    0.00070556184194274485, 0.00074473029862053616, 0.00079324649268314737, 
    0.00085105541519932661, 0.0009180145729506846, 0.00099389198157760479, 
    0.0010783584141007432, 0.0011709885965988293, 0.0012712579924997968, 
    0.0013785459872043204, 0.0014921359105648914, 0.0016112189813876972, 
    0.0017349025020793277, 0.0018622203309571683, 0.0019921440010120021, 
    0.0021235999157361999, 0.0022554842535067936, 0.0023866809092869708, 
    0.0025160848256251095, 0.0026426202131141635, 0.0027652629411922471, 
    0.0028830631046442927, 0.0029951641715125622, 0.0031008239039739833, 
    0.0031994253863355279, 0.0032904948134362265, 0.0033737065829284991, 
    0.0034488860828045032, 0.0035160119986345092, 0.0035752152466056262, 
    0.0036267714210415601, 0.0036710939340626183, 0.0037087196049100332, 
    0.003740293850133059, 0.0037665540800721964, 0.0037883082387185157, 
    0.0038064073147489413, 0.0038217197745646077, 0.0038351036083085067, 
    0.0038473774198263507, 0.0038592873766080272, 0.0038714852602574489, 
    0.0038845066890772256, 0.0038987641235108681, 0.0039145375199520398, 
    0.0039319844087187146, 0.0039511533104153703, 0.0039720009901239462, 
    0.0039944146566754882, 0.0040182316786204555, 0.004043260058332181, 
    0.0040692941856774554, 0.0040961241912835485, 0.0041235382219113872, 
    0.0041513229279804059, 0.0041792537057028841, 0.0042070914180156339, 
    0.0042345766578043677, 0.0042614272649513143, 0.0042873427388229286, 
    0.0043120080471370156, 0.0043351060659493797, 0.0043563304213088249, 
    0.0043753984149773033, 0.0043920677074444359, 0.0044061461308475668, 
    0.0044175075835797255, 0.0044261058622767678, 0.0044319854197497005, 
    0.0044352859532973445, 0.0044362337905977092, 0.0044351236458019284, 
    0.0044322915335169742, 0.004428079022653162, 0.0044228030755854063, 
    0.004416725293578159, 0.0044100362557221284, 0.0044028480354044389, 
    0.0043951975167229613, 0.0043870551744021984, 0.0043783394977855508, 
    0.0043689347455997058, 0.0043587029608686684, 0.0043475024926911332, 
    0.0043351913469514012, 0.0043216348079668579, 0.0043067038076031999, 
    0.0042902745697969841, 0.0042722253991052846, 0.0042524328654674612, 
    0.0042307660384820235, 0.0042070807317921202, 0.0041812138766870403, 
    0.0041529804481904228, 0.0041221681774252514, 0.0040885358203738799, 
    0.0040518132133832959, 0.004011702659048497, 0.0039678824545374015, 
    0.0039200170517905523, 0.0038677698458319159, 0.003810814691830605, 
    0.0037488551211135421, 0.0036816383780388009, 0.0036089730361915083, 
    0.0035307386927891445, 0.003446896839971886, 0.0033574949957835745, 
    0.0032626670145513735, 0.0031626334213755531, 0.0030576987243710594, 
    0.0029482480367928076, 0.0028347433895939394, 0.0027177187408178225, 
    0.0025977704450880165, 0.0024755507589891857, 0.0023517559778900975, 
    0.0022271168250032583, 0.0021023918966821412, 0.0019783614561291905, 
    0.0018558188183975866, 0.0017355647203986422, 0.001618393950130318, 
    0.0015050868116977252, 0.0013963905411275401, 0.0012930002613390679, 
    0.0011955419877883887, 0.0011045519719018377, 0.0010204612839572222, 
    0.00094358795984462876, 0.00087413572790022496, 0.00081220020583736355, 
    0.00075778156087618156, 0.00071080156296295344, 0.0006711231764829715, 
    0.00063856695371458465, 0.00061293511671754839, 0.00059402498697732958, 
    0.00058164340512212157, 0.00057561915206014343, 0.00057581018042167104, 
    0.00058210838974528402, 0.00059444003270288565, 0.00061276234447565654, 
    0.00063705438872508897, 0.00066730410195476307, 0.00070349563591952618, 
    0.00074558764029818017, 0.0007934974904023459, 0.00084708057104391317, 
    0.00090611897017274317, 0.00097030510291256874, 0.0010392403464075861, 
    0.0011124267474697217, 0.0011892716233760843, 0.0012690925127385403, 
    0.0013511227219396833, 0.0014345274058233019, 0.0015184150000850912, 
    0.0016018501223589473, 0.0016838759850566305, 0.0017635328717583538, 
    0.001839887738109973, 0.00191206052086548, 0.001979249014425677, 
    0.0020407491476900482, 0.0020959744175967788, 0.0021444671600693672, 
    0.0021859077544533929, 0.0022201115835805943, 0.0022470247832903443, 
    0.0022667108043793729, 0.0022793397500491279, 0.002285170296038014, 
    0.0022845332609208553, 0.0022778137757567441, 0.0022654395687964832, 
    0.002247861606804923, 0.0022255403478722946, 0.0021989424242270933, 
    0.0021685191319965541, 0.0021347067336671653, 0.0020979086018887878, 
    0.0020584887275695938, 0.0020167543007053781, 0.0019729523408618908, 
    0.0019272625571068157, 0.0018797965384809744, 0.0018306042227657941, 
    0.0017796796798652918, 0.0017269711281708096, 0.0016723926659623647, 
    0.0016158435850166806, 0.0015572257628034059, 0.0014964573294929729, 
    0.0014334978592742318, 0.0013683557298959314, 0.0013010969719054804, 
    0.0012318531410766469, 0.0011608183510161561, 0.0010882499717549889, 
    0.0010144584048152341, 0.00093979659508146068, 0.0008646474250883962, 
    0.00078941000788019557, 0.00071448207578360748, 0.00064024125368503039, 
    0.00056702434002572704, 0.00049510623542590548, 0.00042467674499268259, 
    0.00035582259392301743, 0.00028851614289732283, 0.00022260295972036429, 
    0.00015780959765604419, 9.3744069374115816e-05, 2.9911767287658952e-05, 
    -3.4262356628820298e-05, -9.9411627981380751e-05, 
    -0.00016619096398510136, -0.00023523972482457443, 
    -0.00030714935373935166, -0.00038242350475322707, 
    -0.00046144667584889531, -0.00054446102503155343, 
    -0.00063154883726752019, -0.00072262657613763432, -0.0008174465474407622, 
    -0.00091560771097480705, -0.0010165711140354178, -0.0011196878632842699, 
    -0.0012242204249815411, -0.0013293759285692027, -0.0014343362903879466, 
    -0.0015382870270831787, -0.0016404477279164534, -0.0017400956450260008, 
    -0.0018365928760251562, -0.0019294053914490779, -0.0020181247063222009, 
    -0.0021024791644149573, -0.0021823454286144248, -0.0022577553126790629, 
    -0.0023288863122063875, -0.0023960643615241976, -0.0024597518777424274, 
    -0.0025205330800725494, -0.0025791026724150522, -0.002636248494302231, 
    -0.0026928407046897104, -0.0027498163775669625, -0.00280816002643297, 
    -0.0028688895922311898, -0.00293303424544962, -0.0030016101667085034, 
    -0.0030755970046835832, -0.0031559105040816129, -0.0032433743828608041, 
    -0.0033386935083224503, -0.0034424268962923825, -0.003554964323464996, 
    -0.0036765080972810016, -0.0038070601681086265, -0.0039464164547224224, 
    -0.0040941651673380066, -0.0042496973809944272, -0.0044122239599520535, 
    -0.0045807934699509641, -0.0047543230138313341, -0.0049316271060794777, 
    -0.0051114547583101548, -0.0052925248313624093, -0.0054735667778631411, 
    -0.0056533494933731663, -0.0058307150771028686, -0.0060046095044933813, 
    -0.006174109255793505, -0.006338444418297143, -0.0064970091313381103, 
    -0.0066493746027247481, -0.0067952906401365608, -0.006934682637202056, 
    -0.0070676382831114902, -0.0071943924410936468, -0.0073152989336263503, 
    -0.0074308069379011325, -0.007541428554891789, -0.0076477135524749733, 
    -0.0077502274320954238, -0.0078495327519744786, -0.0079461787116531773, 
    -0.0080406920586216651, -0.0081335761731791655, -0.0082253017813646127, 
    -0.0083163073727716853, -0.0084069964594387942, -0.0084977352739427792, 
    -0.0085888596177245303, -0.0086806670942448701, -0.0087734220758577761, 
    -0.0088673498063487292, -0.0089626375869989068, -0.0090594297906903751, 
    -0.0091578195531976589, -0.0092578436531201222, -0.0093594737185297983, 
    -0.0094626138040424263, -0.0095670910068868277, -0.0096726668951690326, 
    -0.0097790453530510833, -0.0098858815897839777, -0.0099928010552737083, 
    -0.010099415902589177, -0.010205336376809529, -0.010310191105757796, 
    -0.010413638627339348, -0.010515377844623296, -0.010615159774929448, 
    -0.010712792847825486, -0.010808155960165357, -0.010901202293574584, 
    -0.010991969090228378, -0.01108058175938988, -0.011167259662172635, 
    -0.011252306784935088, -0.01133610949036846, -0.011419112763744398, 
    -0.011501794780337334, -0.011584649378545135, -0.011668154513971518, 
    -0.011752754158101758, -0.011838828999272218, -0.011926681626838976, 
    -0.012016520914477712, -0.012108459299925075, -0.012202509383575038, 
    -0.012298591584279763, -0.012396533246263521, -0.012496088573502344, 
    -0.012596942503193306, -0.01269871748939928, -0.012800984845353906, 
    -0.012903267244037031, -0.013005049815828902, -0.013105793303570411, 
    -0.013204950636920145, -0.013301985976158982, -0.013396395506946318, 
    -0.013487725384131155, -0.013575586888091405, -0.013659662745682052, 
    -0.01373971153983812, -0.013815563339052286, -0.013887115738907673, 
    -0.013954315205353318, -0.014017144697125413, -0.014075597680710591, 
    -0.014129664652856627, -0.014179310552091189, -0.014224458893322038, 
    -0.014264982263268571, -0.014300692381301397, -0.014331335624137017, 
    -0.014356589886156826, -0.014376070296568623, -0.01438933243946041, 
    -0.014395884488708524, -0.01439519872457224, -0.014386732687200842, 
    -0.014369951958030954, -0.014344349835310776, -0.014309471016630751, 
    -0.014264931999118383, -0.014210438339801007, -0.01414580046397536, 
    -0.014070943451061557, -0.013985909540671304, -0.01389086011267115, 
    -0.013786070172149814, -0.013671913928517316, -0.013548851553144276, 
    -0.013417401398769247, -0.013278112658069165, -0.013131536404992013, 
    -0.012978201580146431, -0.012818587032468373, -0.01265311431506244, 
    -0.012482136390182631, -0.012305946088722505, -0.012124781841075957, 
    -0.011938846361760576, -0.011748327790452415, -0.011553419199958491, 
    -0.011354347530040316, -0.011151395772576051, -0.01094492373100228, 
    -0.010735385742443596, -0.010523340013355351, -0.010309450539432495, 
    -0.010094481470896789, -0.0098792871438156613, -0.0096647894056815283, 
    -0.0094519524310212287, -0.0092417530291984962, -0.0090351450641153429, 
    -0.0088330232365272949, -0.0086361926077423296, -0.0084453438104592788, 
    -0.008261029367795018, -0.0080836517413609647, -0.0079134564413867424, 
    -0.0077505317059657257, -0.0075948145866340582, -0.0074461052025322763, 
    -0.0073040799082599618, -0.0071683122726607911, -0.0070382910903525773, 
    -0.0069134462245267663, -0.0067931729191569798, -0.0066768578601048689, 
    -0.0065639051221565584, -0.0064537631788100331, -0.0063459471120006338, 
    -0.0062400629964299587, -0.0061358259245234293, -0.0060330626435866298, 
    -0.0059317207796500534, -0.0058318588411418607, -0.0057336255654363245, 
    -0.0056372359355673423, -0.005542942324948957, -0.0054510017557847486, 
    -0.0053616346271334941, -0.0052750017275404112, -0.00519117506274803, 
    -0.0051101239428768654, -0.0050317136400260592, -0.0049557068957110885, 
    -0.0048817711963436107, -0.004809492150540844, -0.0047383785314277747, 
    -0.0046678793070574383, -0.004597387735333444, -0.0045262611915941296, 
    -0.0044538405039085804, -0.0043794824554768737, -0.0043025871900856218, 
    -0.0042226253961048128, -0.0041391637419685235, -0.0040518809865891592, 
    -0.0039605802502645608, -0.0038651955156519461, -0.0037657945701610844, 
    -0.0036625817849854094, -0.0035559013605079783, -0.0034462297957871747, 
    -0.0033341734444799044, -0.0032204635840368152, -0.0031059414315191339, 
    -0.0029915473053564391, -0.0028783057161096549, -0.0027672957636561309, 
    -0.002659631202961546, -0.0025564263363462561, -0.0024587602013701917, 
    -0.0023676435186349531, -0.0022839846621977634, -0.0022085654464436963, 
    -0.002142027014486726, -0.0020848659921528642, -0.0020374415298237939, 
    -0.0019999858610397383, -0.0019726146848557486, -0.0019553343310242874, 
    -0.0019480353872234611, -0.0019504810041605816, -0.0019622915214984847, 
    -0.0019829330362296591, -0.0020117186315314842, -0.0020478225307928315, 
    -0.0020903021238824287, -0.0021381243064199141, -0.0021901974315606271, 
    -0.0022453993982864359, -0.0023026041797497253, -0.0023606941463740873, 
    -0.0024185757216552937, -0.002475194278057874, -0.0025295411801190089, 
    -0.0025806646147345986, -0.0026276826271975852, -0.0026697972389791926, 
    -0.0027063084485202311, -0.0027366289384274487, -0.0027602922638063697, 
    -0.0027769628843267763, -0.0027864413863587911, -0.0027886660941724953, 
    -0.0027837148333909557, -0.0027718027833198359, -0.0027532768697559103, 
    -0.0027286001176197719, -0.0026983411552447124, -0.0026631521123665403, 
    -0.0026237513928672029, -0.0025808986724418863, -0.0025353733041462694, 
    -0.0024879480787573282, -0.002439366167436566, -0.0023903176255872832, 
    -0.0023414239715648082, -0.0022932257150918432, -0.0022461728635588532, 
    -0.0022006214936748001, -0.0021568365430434579, -0.0021149947949182946, 
    -0.0020751906566428965, -0.0020374377670498581, -0.0020016825911496113, 
    -0.0019678142068862048, -0.0019356747156321619, -0.0019050707061260145, 
    -0.0018757828037054356, -0.0018475786407653137, -0.0018202167727622443, 
    -0.0017934575289322819, -0.001767065577123235, -0.0017408240548284245, 
    -0.0017145475647727941, -0.0016881030992084902, -0.0016614262437533991, 
    -0.0016345417199002594, -0.0016075849956484454, -0.0015808129220877798, 
    -0.0015546063722774739, -0.0015294647140066348, -0.001505995239250816, 
    -0.0014848915270689962, -0.0014669054285674432, -0.001452817565945811, 
    -0.0014434020748756819, -0.001439397528620314, -0.001441473306272833, 
    -0.0014502025414122441, -0.0014660343659355873, -0.0014892779744886198, 
    -0.0015200891275654695, -0.0015584633463113866, -0.0016042379065928001, 
    -0.0016571052907118, -0.0017166263963710822, -0.0017822502030690344, 
    -0.0018533356769392293, -0.0019291732281210335, -0.0020090071934039883, 
    -0.0020920539067559247, -0.0021775207343244728, -0.0022646267856239162, 
    -0.0023526179374240837, -0.0024407910865138875, -0.0025285157506765238, 
    -0.0026152546990833715, -0.0027005785602307285, -0.0027841836929858163, 
    -0.0028658964493730671, -0.002945671249763472, -0.0030235810135946107, 
    -0.0030997998219955084, -0.0031745852444445919, -0.0032482547781891411, 
    -0.0033211694539832205, -0.0033937147897760097, -0.0034662803757140002, 
    -0.0035392544908131708, -0.0036130134489423768, -0.0036879173169960533, 
    -0.0037643205551878283, -0.0038425767063354549, -0.003923049009880164, 
    -0.0040061218040386348, -0.0040922038590701483, -0.0041817347440401779, 
    -0.0042751793679685788, -0.0043730180177392851, -0.0044757283172552238, 
    -0.0045837624246037323, -0.0046975200516200305, -0.004817316828135753, 
    -0.0049433641617833684, -0.005075745511824401, -0.0052144071803744843, 
    -0.0053591601597571988, -0.0055096836810025474, -0.0056655322714298136, 
    -0.005826153190083872, -0.0059908924288860198, -0.0061590064378660627, 
    -0.0063296577221631286, -0.0065019257918316267, -0.0066747981713155182, 
    -0.0068471769512421024, -0.007017885311539681, -0.0071856732882019797, 
    -0.0073492412977771322, -0.0075072531865052507, -0.0076583644482396693, 
    -0.007801255874999441, -0.0079346551735916711, -0.008057366048353911, 
    -0.0081682929602393938, -0.0082664634713743718, -0.0083510438660883753, 
    -0.0084213503620715648, -0.0084768649483256235, -0.0085172274821542493, 
    -0.0085422361583761732, -0.0085518403778876897, -0.0085461375277234627, 
    -0.0085253640245810877, -0.0084898913479976943, -0.0084402119452838594, 
    -0.0083769334370209347, -0.0083007753962396902, -0.008212562870970953, 
    -0.0081132250101041917, -0.0080037865567597483, -0.0078853588938932583, 
    -0.0077591320183603117, -0.0076263595762961376, -0.0074883316520926602, 
    -0.0073463457860346382, -0.007201680537685295, -0.0070555755380986782, 
    -0.0069092112821159766, -0.0067637099193534203, -0.0066201401635363581, 
    -0.0064795293306365385, -0.0063428787902803669, -0.0062111707042083013, 
    -0.0060853682450308141, -0.0059663920015945778, -0.0058550901361333861, 
    -0.0057521974840728587, -0.0056582946207635668, -0.0055737725285611326, 
    -0.005498818342765931, -0.0054334167743696222, -0.0053773653481693738, 
    -0.0053303041960433067, -0.0052917496181894754, -0.0052611275193489553, 
    -0.0052378067671923403, -0.0052211240658585891, -0.0052104110343537307, 
    -0.0052050114491924253, -0.0052043040422034559, -0.0052077171834156305, 
    -0.0052147491372858774, -0.0052249797942154289, -0.0052380838762361047, 
    -0.0052538392950986544, -0.0052721216833978152, -0.0052928951308297365, 
    -0.0053161900303655609, -0.0053420774336281028, -0.0053706413413365708, 
    -0.0054019469708628939, -0.0054360245222204485, -0.0054728478297399758, 
    -0.0055123206106661542, -0.0055542697760107215, -0.0055984423519902429, 
    -0.0056445033536158783, -0.0056920362861938153, -0.0057405465809709996, 
    -0.0057894603075327473, -0.0058381238135035195, -0.0058858049620944194, 
    -0.0059316910086256299, -0.0059748866747456235, -0.0060144229361625097, 
    -0.0060492514975842666, -0.0060782574629199195, -0.0061002706059289482, 
    -0.0061140859718215208, -0.0061184899937027099, -0.0061122911568369659, 
    -0.0060943506571573486, -0.006063614379039327, -0.0060191457187965449, 
    -0.0059601447172440937, -0.0058859662199789459, -0.0057961143691296554, 
    -0.0056902306084066837, -0.0055680639968431304, -0.0054294470590560435, 
    -0.0052742711143392608, -0.0051024812989818348, -0.0049140875500130066, 
    -0.00470918591037333, -0.0044879826093798961, -0.0042508084331004618, 
    -0.0039981283672725441, -0.003730551411379875, -0.0034488264344704417, 
    -0.0031538318007368485, -0.0028465607177169984, -0.0025281194942064372, 
    -0.002199702380417343, -0.0018625812738491919, -0.0015180933441593294, 
    -0.0011676271606144459, -0.00081260961210442666, -0.00045448688430818314, 
    -9.4720274148621733e-05, 0.00026523215439748071, 0.00062391947482141137, 
    0.00097990738575910708, 0.001331787344287651, 0.0016781828010880946, 
    0.0020177671239739957, 0.0023492762867795359, 0.0026715341667796423, 
    0.0029834708190954115, 0.0032841367167237095, 0.0035727255427608707, 
    0.0038485757978185655, 0.0041111787893991295, 0.0043601695152405166, 
    0.0045953278645709328, 0.0048165750733625157, 0.0050239709151322148, 
    0.005217708890179272, 0.0053981229768719045, 0.005565680286953408, 
    0.0057209847119074151, 0.0058647788977806321, 0.0059979376491199011, 
    0.0061214648758691724, 0.0062364825538477053, 0.0063442156828246313, 
    0.0064459708745118246, 0.0065431040382301934, 0.0066369914342676436, 
    0.006728991376916179, 0.0068204097823824882, 0.006912479143308314, 
    0.0070063347877970493, 0.0071029942671921812, 0.0072033570843454582, 
    0.0073082013978229016, 0.0074181829842782255, 0.0075338388575428754, 
    0.0076555991359459914, 0.0077837902430893061, 0.0079186399293081113, 
    0.0080602835642252547, 0.0082087623657478952, 0.0083640246104881751, 
    0.0085259238407402078, 0.0086942244473135755, 0.008868611441593446, 
    0.009048711797168275, 0.0092341105431677211, 0.0094243700611716386, 
    0.0096190497981732577, 0.0098177164687862552, 0.010019951380130872, 
    0.010225343848487027, 0.010433489028806604, 0.010643972995373136, 
    0.010856348538136067, 0.011070106861283473, 0.011284641775724247, 
    0.011499220782850761, 0.011712950954129752, 0.01192477040669367, 
    0.01213344770407465, 0.012337614204343927, 0.01253581263927364, 
    0.012726540036804847, 0.012908300595501234, 0.013079646505704963, 
    0.013239204974931128, 0.013385703546762304, 0.013517978488844342, 
    0.013634989181201648, 0.013735836559986319, 0.013819776931222607, 
    0.013886236056858436, 0.013934823744706872, 0.013965338065051482, 
    0.013977757649510082, 0.013972237415686668, 0.013949091985196786, 
    0.01390877455396175, 0.013851858539506287, 0.013779009427991758, 
    0.013690957988838848, 0.013588476934319081, 0.013472358979289032, 
    0.013343408073845256, 0.013202417841198617, 0.013050169646030362, 
    0.012887428120454488, 0.012714937332844864, 0.012533423216644152, 
    0.012343588824740645, 0.012146127285331676, 0.011941713180810342, 
    0.011731006101705212, 0.011514646634196751, 0.011293258885269214, 
    0.011067429246243822, 0.010837702613702822, 0.010604558932566682, 
    0.01036840172202768, 0.01012953896829287, 0.0098881837911196889, 
    0.0096444509654288069, 0.0093983595147484143, 0.0091498545962831, 
    0.0088988133639786304, 0.0086450613576709162, 0.0083883885996520798, 
    0.0081285616049313839, 0.0078653256096807723, 0.0075983839824078116, 
    0.007327391276234778, 0.0070519193296741493, 0.0067714654906220976, 
    0.0064854602684479689, 0.0061932917162547249, 0.0058943396659838828, 
    0.005588014973355742, 0.0052737899020579059, 0.0049512316648722661, 
    0.0046200158188174894, 0.0042799553269639787, 0.0039309976085721019, 
    0.0035732467997881931, 0.0032069525797088832, 0.002832508579668892, 
    0.002450448735965143, 0.0020614315934091463, 0.0016662319505576283, 
    0.0012657408158606252, 0.00086095619059932274, 0.00045297447504153988, 
    4.2993993860948089e-05, -0.00036769350277814392, -0.00077770735029595521, 
    -0.0011855988358881893, -0.0015898685303297432, -0.0019889939301657444, 
    -0.002381457286489262, -0.0027657809662859014, -0.0031405496717233855, 
    -0.003504437673702484, -0.0038562376639846305, -0.0041948832869830111, 
    -0.0045194707747213915, -0.0048292753076737797, -0.0051237473606153472, 
    -0.0054025128117845623, -0.0056653652611188309, -0.0059122637555132406, 
    -0.0061433344764935368, -0.0063588702484164619, -0.0065593337922562412, 
    -0.0067453438732234016, -0.0069176710345700545, -0.007077214089415201, 
    -0.0072249719629577684, -0.0073620069448369395, -0.0074894102759473745, 
    -0.0076082513845851345, -0.007719535448131018, -0.0078241549698523059, 
    -0.0079228476126401246, -0.0080161514348205554, -0.0081043759968604141, 
    -0.0081875842025611306, -0.0082655841101290598, -0.0083379499848032328, 
    -0.0084040536321185744, -0.0084631194508879969, -0.0085142773748313177, 
    -0.0085566231007005878, -0.0085892640811623608, -0.0086113589159267888, 
    -0.008622142331649367, -0.0086209328570482913, -0.0086071453791392808, 
    -0.0085802867743866636, -0.0085399635438732184, -0.0084858775509903759, 
    -0.0084178362352971443, -0.0083357473071223962, -0.0082396315828845972, 
    -0.00812962954792921, -0.0080060079725694754, -0.0078691722166078625, 
    -0.0077196780992950798, -0.0075582582092791929, -0.0073858331057360237, 
    -0.0072035277107627858, -0.0070126741739437674, -0.0068147921773962098, 
    -0.0066115683935395048, -0.0064048094861649495, -0.006196380074153407, 
    -0.0059881293161464181, -0.0057818235844960897, -0.0055790703589742637, 
    -0.0053812597317851665, -0.0051895126130876955, -0.0050046464184065479, 
    -0.0048271625657028156, -0.0046572530961569584, -0.0044948186592586046, 
    -0.0043394947816950804, -0.0041906856196188644, -0.0040476090130707196, 
    -0.0039093295819903669, -0.0037748037768332078, -0.0036429201121087199, 
    -0.003512530969350018, -0.0033824919925411301, -0.0032516975916001053, 
    -0.003119097074855747, -0.0029837177917361388, -0.0028446739482659612, 
    -0.0027011546739994551, -0.0025524236056721954, -0.0023978094958478032, 
    -0.0022366975913444848, -0.0020685236424678793, -0.0018927785054009781, 
    -0.0017090104019599275, -0.0015168370668123957, -0.0013159547385741515, 
    -0.0011061508185004022, -0.00088731239700559953, -0.0006594287681847659, 
    -0.00042259841815946273, -0.00017701486855250018, 7.7030956752506281e-05, 
    0.00033916150061490472, 0.0006089258672571686, 0.00088578905765111272, 
    0.0011691445962562692, 0.0014582935704905216, 0.0017524525494566241, 
    0.0020507632196591755, 0.002352301222068416, 0.0026561026099793084, 
    0.002961183464317146, 0.0032665537132123535, 0.0035712375042860388, 
    0.0038742873423962812, 0.0041747953547329984, 0.0044718871345096082, 
    0.0047647328559635585, 0.0050525420445553379, 0.0053345701194592995, 
    0.0056101159340020221, 0.0058785093843762588, 0.0061391087847574265, 
    0.0063912888722382826, 0.006634452659635112, 0.0068680510623198646, 
    0.007091615453219938, 0.0073047836824423392, 0.0075073371771053809, 
    0.0076992083953212592, 0.007880468517519593, 0.0080512994926188308, 
    0.0082119598137698098, 0.0083627423632540304, 0.0085039289155245112, 
    0.0086357540938029869, 0.0087583852083078506, 0.0088718932667114937, 
    0.0089762621350653153, 0.0090713904262857865, 0.009157092815821952, 
    0.0092331042889563578, 0.0092990818717480824, 0.009354579611333274, 
    0.0093990378810438115, 0.0094317532439024149, 0.0094518650333221994, 
    0.0094583809097806698, 0.0094502504178852597, 0.0094265066448059008, 
    0.0093863919791976232, 0.0093294621559445439, 0.0092556301018635219, 
    0.0091651547663469841, 0.0090586092416365081, 0.0089368237663534755, 
    0.0088008341558064376, 0.0086518349197255498, 0.0084911516756948479, 
    0.0083202144942064477, 0.0081405343442151733, 0.0079536942533374351, 
    0.0077613361612508761, 0.0075651586883477111, 0.0073668865828278793, 
    0.0071682501735083953, 0.0069709627551404127, 0.0067766699069470972, 
    0.0065869344419271321, 0.0064031812196341494, 0.0062266773443550704, 
    0.0060585043755417029, 0.0058995312458963254, 0.0057504006202007312, 
    0.0056115284484414395, 0.0054831069755097049, 0.0053651070545993676, 
    0.0052573105166435537, 0.0051593258377972415, 0.0050706295488354815, 
    0.0049905867054433331, 0.0049185062373137455, 0.0048536790240254852, 
    0.0047954276332995097, 0.0047431288237215234, 0.0046962307668785607, 
    0.0046542577491954897, 0.0046168148092982347, 0.0045835620695883102, 
    0.0045542055751700344, 0.0045284885985354909, 0.0045061841572699686, 
    0.0044870748785739208, 0.0044709663931169763, 0.0044576893607520852, 
    0.0044471274819564473, 0.0044392404867797559, 0.0044340963142921533, 
    0.004431900303232152, 0.0044330202202149758, 0.0044379830709136425, 
    0.0044474553025463381, 0.0044622248192269171, 0.0044831516378553166, 
    0.004511121975153163, 0.0045469975317603039, 0.0045915769074054095, 
    0.0046455519332279467, 0.0047094767224915282, 0.0047837392130333205, 
    0.0048685397559486603, 0.0049638676670386832, 0.0050694863852819884, 
    0.0051849161343379101, 0.0053094221490733937, 0.0054420092093354841, 
    0.0055814477819313875, 0.0057263043356074843, 0.0058749769862497282, 
    0.0060257562617147533, 0.0061768691553704975, 0.0063265433688499354, 
    0.0064730522265731751, 0.006614773424652119, 0.0067502175269155392, 
    0.0068780863350087051, 0.0069972994063851558, 0.0071070116948744365, 
    0.0072066432983600255, 0.0072958741992854093, 0.0073746320791400564, 
    0.0074430569053595772, 0.0075014486181765568, 0.0075502381883509858, 
    0.0075899457062995404, 0.0076211440133297625, 0.0076444361393299895, 
    0.0076604215575122791, 0.0076696690433855344, 0.0076727079845640622, 
    0.0076700126126152514, 0.0076620087226502162, 0.0076490619240109298, 
    0.0076314803024959237, 0.0076095231160721536, 0.0075834075421542498, 
    0.0075533184326567948, 0.0075193967972384552, 0.00748174290714079, 
    0.0074404100995591688, 0.0073954086083135324, 0.0073466967058069066, 
    0.0072941913465559161, 0.0072377787244531254, 0.0071773092609926075, 
    0.0071126145495426533, 0.0070434995318224749, 0.0069697759643625838, 
    0.0068912509349603199, 0.00680774196695533, 0.006719081922430036, 
    0.0066251212369785014, 0.0065257439684558369, 0.0064208829764101898, 
    0.0063105276058360782, 0.0061947659873086008, 0.0060737907851738764, 
    0.0059479355515736519, 0.0058177086207560373, 0.0056838052614161224, 
    0.0055471420651869051, 0.0054088753905521371, 0.0052704024598024327, 
    0.0051333556248532915, 0.0049995705437322424, 0.0048710511538407296, 
    0.0047499026916228123, 0.0046382516986680873, 0.0045381630615778448, 
    0.0044515534981882663, 0.0043800997463941428, 0.0043251510895567355, 
    0.0042876715943489466, 0.0042681948380550753, 0.0042667924194863252, 
    0.0042830906661122971, 0.0043162962221615572, 0.0043652627187762685, 
    0.0044285531006082448, 0.0045045200411466769, 0.0045913772053596813, 
    0.0046872705191862013, 0.0047903561147374426, 0.0048988327724743671, 
    0.0050109965634118105, 0.0051252894070580668, 0.0052403385004121585, 
    0.0053549535450216363, 0.0054681407576491238, 0.0055790860569140902, 
    0.0056871625719082499, 0.005791901575316288, 0.0058929928317239012, 
    0.0059902693650348863, 0.0060836954414593275, 0.0061733468622281731, 
    0.0062594097338777481, 0.006342165828065475, 0.0064219844198396651, 
    0.0064992983639996383, 0.00657459323971522, 0.0066483899256680207, 
    0.006721246354493832, 0.0067937415376574497, 0.0068664830619639804, 
    0.0069401232847500641, 0.0070153645642003631, 0.0070929796668346649, 
    0.0071738162328313431, 0.0072587990518104325, 0.0073488990497390314, 
    0.0074451061416674503, 0.0075483786081626822, 0.00765960530018003, 
    0.0077795626182019942, 0.0079088824227803358, 0.0080480150205218051, 
    0.0081972143679085833, 0.0083565400159897538, 0.0085258796776710652, 
    0.0087049658434131417, 0.0088933996332591705, 0.0090906769318595433, 
    0.0092962072239989712, 0.0095093095628058597, 0.0097292028238543365, 
    0.0099549929708954484, 0.010185628217310436, 0.010419870904229014, 
    0.010656273122219357, 0.010893155540906491, 0.011128619990772505, 
    0.011360574117675272, 0.011586772541247885, 0.011804871008841252, 
    0.012012487914238401, 0.012207295081868342, 0.012387063055928486, 
    0.012549734119056848, 0.01269345925253266, 0.01281663833927164, 
    0.012917959313785969, 0.012996418994706558, 0.013051340270266313, 
    0.013082361667569828, 0.013089415320656758, 0.013072695271521587, 
    0.013032663366327024, 0.012970050323789076, 0.012885887528399802, 
    0.012781530078130853, 0.012658671793777764, 0.012519355217361168, 
    0.012365925302252986, 0.012200984683674197, 0.012027362262732384, 
    0.011848025898193427, 0.011666025566774714, 0.011484402704759039, 
    0.011306093249593297, 0.011133809778067157, 0.010969954304093095, 
    0.010816530615623866, 0.010675136159435432, 0.010546946516366021, 
    0.010432756129232508, 0.010332974631711272, 0.01024766901511982, 
    0.010176582949463574, 0.010119191999610882, 0.010074765427383326, 
    0.01004241543383072, 0.010021129037323268, 0.010009808691988337, 
    0.010007283703832855, 0.010012301519238227, 0.01002348897468998, 
    0.010039334358942704, 0.010058157998972646, 0.010078088707359253, 
    0.010097049957431584, 0.010112756206398394, 0.010122744929037123, 
    0.010124375611281041, 0.010114885362552525, 0.010091453903059782, 
    0.010051240551656907, 0.0099914506307837644, 0.0099093681407829877, 
    0.0098023841620624962, 0.009668023281447639, 0.0095039608290364824, 
    0.0093080445043442414, 0.0090782805028679445, 0.0088128649442811118, 
    0.0085101687997211333, 0.0081687331090264693, 0.0077872743325936265, 
    0.0073646911197340426, 0.0069000991276906287, 0.0063928392636464406, 
    0.0058425132672248956, 0.0052490251917267821, 0.0046126040213695582, 
    0.0039338079505795067, 0.0032135519003120717, 0.0024531293691758263, 
    0.0016542741853807989, 0.00081922340854987427, -4.9210333176877199e-05, 
    -0.00094759935494678456, -0.0018719370085914884, -0.0028176942879609293, 
    -0.0037799223658502136, -0.0047533861141832254, -0.0057326262417477089, 
    -0.0067120666655018854, -0.0076860279926545417, -0.0086488338270431769, 
    -0.0095948454079084547, -0.010518550238398178, -0.011414656595435115, 
    -0.012278173251959056, -0.013104504351015574, -0.013889540501412345, 
    -0.014629757476344787, -0.015322232359876417, -0.015964680365706231, 
    -0.016555505724649835, -0.017093804518183871, -0.017579331381128164, 
    -0.018012525672011746, -0.018394460096043237, -0.018726809844630255, 
    -0.01901181670196184, -0.019252196254688991, -0.019451150100572301, 
    -0.019612300406386455, -0.01973965530695777, -0.019837591529485762, 
    -0.019910788261126286, -0.019964181142952498, -0.020002848881431983, 
    -0.020031909649045759, -0.020056375255542953, -0.020081008035746896, 
    -0.020110143306267265, -0.020147581529782722, -0.020196468836204774, 
    -0.020259237581644399, -0.020337547986590643, -0.020432318272517808, 
    -0.020543747764751444, -0.020671403435982956, -0.020814225005555784, 
    -0.020970571640080003, -0.02113820718060333, -0.021314274747467585, 
    -0.021495357150707294, -0.021677501021861847, -0.021856363012634657, 
    -0.022027374595801397, -0.022185929291270688, -0.022327596574863558, 
    -0.022448300453677746, -0.022544431466659281, -0.022612923421508401, 
    -0.02265130409117018, -0.022657736507666754, -0.022630979373771672, 
    -0.022570432575202068, -0.022476069204549122, -0.022348366485798955, 
    -0.022188293525194223, -0.021997073987424804, -0.021776106523704371, 
    -0.021526790119887094, -0.021250431145185173, -0.020948062515270188, 
    -0.020620481529042941, -0.020268202355307127, -0.019891490842336199, 
    -0.019490423675398136, -0.019065045574178464, -0.018615507952546909, 
    -0.018142135638797612, -0.01764570800168961, -0.017127581426946863, 
    -0.01658980146507328, -0.016035188334431686, -0.015467113117892881, 
    -0.014889560051068498, -0.014306799468696851, -0.013723140940174348, 
    -0.013142653435514367, -0.012568907200759672, -0.01200483385081047, 
    -0.011452752568822002, -0.010914384322090227, -0.010391032102215172, 
    -0.0098837707756510313, -0.0093934831720388738, -0.0089208748698496217, 
    -0.0084664393788260548, -0.0080303441678876569, -0.007612484832932245, 
    -0.0072126970149904643, -0.0068307130823590714, -0.0064661014694550288, 
    -0.0061180883973944913, -0.0057854278270354732, -0.0054660302101407678, 
    -0.0051572472691003863, -0.0048556141267997845, -0.0045573130600854526, 
    -0.0042582034586958212, -0.003954294103057478, -0.0036418710840130132, 
    -0.0033178685749254487, -0.0029798218143694175, -0.0026261222892088702, 
    -0.0022562379221817658, -0.0018708581099617114, -0.001471642309669646, 
    -0.0010614967676505173, -0.00064280115033850155,
  // Fqt-F(3, 0-1999)
    1, 0.99823067080000405, 0.99295429850473882, 0.98426504801492232, 
    0.97231595183133446, 0.95731275191775378, 0.93950594196421144, 
    0.91918156677484786, 0.89665136846823745, 0.87224285159782022, 
    0.84628976115175503, 0.81912337509324173, 0.79106490360065052, 
    0.76241915137945437, 0.73346953316893426, 0.70447442173469388, 
    0.67566474206366378, 0.64724271278940337, 0.61938157037956276, 
    0.59222610532835918, 0.56589387039426353, 0.54047688551296735, 
    0.51604369664723793, 0.49264165356156542, 0.47029928397650905, 
    0.44902868282350794, 0.4288278420189407, 0.40968288380029882, 
    0.39157014688315539, 0.37445812683687102, 0.35830924809491632, 
    0.34308143670285135, 0.32872952061556515, 0.31520641820971312, 
    0.30246415369345969, 0.29045470279074614, 0.27913068263973789, 
    0.26844591600955048, 0.25835587832756668, 0.24881805254826697, 
    0.23979219842466079, 0.23124056380432015, 0.22312801006596442, 
    0.21542209753980091, 0.20809308719809866, 0.20111389890871725, 
    0.19446002023149886, 0.18810937046881479, 0.18204214131884622, 
    0.1762406169181403, 0.17068898626310275, 0.16537314278128687, 
    0.16028049052827895, 0.15539975532621156, 0.15072078801895222, 
    0.14623438319606744, 0.14193210185159474, 0.13780610135904237, 
    0.13384898109682003, 0.13005364213382153, 0.1264131744353833, 
    0.1229207663389793, 0.1195696486375261, 0.11635306856527562, 
    0.11326428667854892, 0.11029660202413269, 0.10744339209591484, 
    0.10469815484740774, 0.1020545632225391, 0.099506503742290406, 
    0.097048116472322907, 0.094673810592642363, 0.092378282848023296, 
    0.090156501181396953, 0.088003692790303789, 0.085915309600138393, 
    0.083886994530780343, 0.081914550100116695, 0.079993906291706385, 
    0.078121101433592993, 0.076292272676923706, 0.074503655117679174, 
    0.072751608978765536, 0.071032639429364886, 0.069343434160673262, 
    0.067680900566004343, 0.066042196956380514, 0.064424765973212866, 
    0.062826356289006069, 0.061245041892496702, 0.059679233957786862, 
    0.058127681097306934, 0.056589465069776974, 0.055063990590165701, 
    0.053550972992092827, 0.05205042033277528, 0.05056261156686867, 
    0.049088077238723722, 0.047627564228023639, 0.04618200299062656, 
    0.044752470449557817, 0.04334016313523386, 0.041946364413511149, 
    0.040572421086250872, 0.039219727223294025, 0.037889702838322506, 
    0.036583771106976297, 0.035303337126246483, 0.034049771276337362, 
    0.03282437794512625, 0.031628377010892217, 0.030462876881394825, 
    0.029328863124593367, 0.028227183166082876, 0.027158539984944829, 
    0.026123489867793035, 0.02512244751961875, 0.024155692285049941, 
    0.023223396054927098, 0.022325647680383441, 0.021462491477575323, 
    0.020633964178442946, 0.019840136791165329, 0.01908115629957639, 
    0.018357275199912863, 0.017668883242869523, 0.017016523261036916, 
    0.01640090152901778, 0.015822881817297404, 0.015283469837105129, 
    0.014783778985022693, 0.014324988495310217, 0.013908285620652151, 
    0.01353480035112401, 0.013205540022291887, 0.012921321474769945, 
    0.012682714817270724, 0.012489993686629872, 0.012343098129441198, 
    0.012241613082996755, 0.012184749299904957, 0.012171349825726287, 
    0.012199893992793573, 0.012268520936267853, 0.012375046863771619, 
    0.012517005232599384, 0.012691684927826902, 0.012896179984732701, 
    0.013127439722130093, 0.013382318649439239, 0.013657634907368777, 
    0.01395022092840313, 0.014256968902034933, 0.014574864504740055, 
    0.014901024737304475, 0.015232708426954504, 0.015567333350631112, 
    0.015902471946506295, 0.016235842924165477, 0.016565287561759987, 
    0.016888749121122586, 0.017204242781791747, 0.017509830808016085, 
    0.017803604535347527, 0.018083684750355256, 0.018348228956426998, 
    0.018595465561603342, 0.018823733524642464, 0.019031538605225051, 
    0.019217610420391586, 0.019380964274345613, 0.019520959848001441, 
    0.019637349854251748, 0.019730307713124125, 0.019800427583952403, 
    0.019848700727825141, 0.019876462251556735, 0.019885321600667236, 
    0.01987708914431845, 0.019853692771585219, 0.019817100971068785, 
    0.019769255029584435, 0.019712011942876608, 0.019647097203331094, 
    0.01957608069692272, 0.01950036122747863, 0.019421168355008168, 
    0.019339567376998996, 0.019256475380846676, 0.019172675773091934, 
    0.019088837859370173, 0.019005530887663366, 0.018923237011777668, 
    0.018842356686056178, 0.018763214593009472, 0.018686053828457512, 
    0.01861103424771416, 0.018538227238624957, 0.018467612612224293, 
    0.018399082732751995, 0.018332445214474802, 0.018267429275576071, 
    0.018203696023928288, 0.018140852888612696, 0.018078468319162506, 
    0.018016093464157279, 0.017953287516561917, 0.017889637766095513, 
    0.017824786945566509, 0.017758446310265033, 0.017690408076053859, 
    0.017620546951557597, 0.017548815071121465, 0.017475224714643165, 
    0.01739981719665265, 0.017322632633553915, 0.017243671481832083, 
    0.017162858951622874, 0.017080007191753975, 0.016994788631542957, 
    0.016906714868315086, 0.016815125052876405, 0.016719186956696712, 
    0.016617906039928177, 0.01651014474098832, 0.016394651277307288, 
    0.016270089147796894, 0.016135086217646269, 0.015988271280369195, 
    0.0158283258009786, 0.015654023652152245, 0.015464268794702906, 
    0.015258127983449173, 0.015034857779028736, 0.014793925029268188, 
    0.014535013985610763, 0.014258039620075496, 0.013963148103074667, 
    0.013650712578365407, 0.013321324280576868, 0.012975767265425348, 
    0.012615000282359774, 0.012240125464376217, 0.011852358008880643, 
    0.011452994029455628, 0.011043384449183551, 0.010624911210307097, 
    0.010198966088342575, 0.0097669320078688573, 0.0093301763273854425, 
    0.008890038631667558, 0.0084478385023535277, 0.0080048845274059942, 
    0.0075624790352707381, 0.0071219245900892049, 0.0066845252854706412, 
    0.0062515864932119894, 0.005824408430153743, 0.0054042778157187719, 
    0.0049924616348032812, 0.0045901964426501912, 0.0041986722293414951, 
    0.00381902364462637, 0.0034523017525231181, 0.0030994475653511712, 
    0.0027612608369619873, 0.0024383619698509712, 0.0021311564690992633, 
    0.0018398055397232456, 0.0015642014337074771, 0.0013039487223300531, 
    0.0010583538783839018, 0.00082642842752742951, 0.00060689844140861802, 
    0.00039822384851181069, 0.00019862742525122046, 6.1318985234767994e-06, 
    -0.00018139442042096224, -0.00036617663648445863, -0.0005504651970776297, 
    -0.0007364605688643162, -0.00092623403076071988, -0.0011216481670729395, 
    -0.0013242881839979877, -0.0015354016063453256, -0.0017558539632486561, 
    -0.0019861028525925322, -0.0022261847073076911, -0.0024757267030426217, 
    -0.0027339607557822767, -0.0029997612186117482, -0.0032716880925025573, 
    -0.0035480364557076778, -0.0038268940770129715, -0.004106196180039462, 
    -0.004383780183940607, -0.0046574413891546781, -0.0049249709437061738, 
    -0.0051842021120870807, -0.0054330433873011064, -0.0056695106496371193, 
    -0.0058917547049550647, -0.0060980896658248121, -0.0062870164629095686, 
    -0.0064572441339999335, -0.0066077055073065528, -0.0067375700377138407, 
    -0.0068462556018692158, -0.0069334358446818739, -0.006999039204081587, 
    -0.007043242357195752, -0.0070664443553590138, -0.0070692393095253721, 
    -0.0070523818382394283, -0.0070167515656494621, -0.0069633212425613475, 
    -0.0068931276405055936, -0.0068072493467817808, -0.0067067873607528777, 
    -0.0065928443777287888, -0.0064665082005351364, -0.0063288395378977144, 
    -0.006180858950941801, -0.0060235385690204446, -0.0058577910306488179, 
    -0.0056844669626832439, -0.0055043518682781059, -0.0053181617260676817, 
    -0.0051265413373460357, -0.0049300660554631908, -0.0047292391116448892, 
    -0.0045244957542931565, -0.0043162086185571788, -0.0041046968227424051, 
    -0.0038902302513382377, -0.0036730342539322042, -0.0034532901130002167, 
    -0.0032311354931373213, -0.0030066624441850132, -0.0027799121947476094, 
    -0.0025508743983592287, -0.002319485230692345, -0.0020856314080996479, 
    -0.0018491472931647982, -0.0016098291202405327, -0.001367437848323178, 
    -0.0011217165917189575, -0.00087240358627556445, -0.00061924597878591987, 
    -0.00036201693091417962, -0.00010053168549325906, 0.0001653410464203186, 
    0.000435666428730888, 0.00071043356440234453, 0.00098954562324551714, 
    0.0012728135735403606, 0.0015599535085744692, 0.001850595398366536, 
    0.0021443010538186136, 0.0024405786136587099, 0.0027388995544846582, 
    0.0030386991220256896, 0.003339364949464684, 0.003640207933287089, 
    0.0039404281943383936, 0.0042390751829679977, 0.004535016588607544, 
    0.0048269124711024921, 0.0051132068524795335, 0.0053921373371593577, 
    0.0056617596709337232, 0.0059199850716749247, 0.0061646314991432929, 
    0.0063934823964029754, 0.0066043496505016012, 0.0067951401319069939, 
    0.0069639161165543336, 0.0071089500146685235, 0.0072287666748473249, 
    0.0073221794017992343, 0.0073883051192238786, 0.0074265592852236191, 
    0.0074366390194507094, 0.0074184986916433771, 0.0073723108427810827, 
    0.0072984336866266375, 0.0071973752330868855, 0.0070697653312260245, 
    0.0069163448675926562, 0.006737953731447162, 0.0065355342751237163, 
    0.0063101275580537183, 0.0060628711597801978, 0.0057949925244754385, 
    0.0055078028543976611, 0.005202692704231477, 0.0048811278423656285, 
    0.0045446458261453318, 0.004194857652575797, 0.0038334465379059597, 
    0.0034621652639137503, 0.0030828319113467956, 0.0026973246559371549, 
    0.0023075756324892659, 0.0019155547761617363, 0.001523263404760087, 
    0.0011327273331447475, 0.00074599070401021534, 0.00036511703047797418, 
    -7.8122683961757804e-06, -0.00037070340199625926, 
    -0.00072145682016659142, -0.0010579906178622524, -0.0013782676783346518, 
    -0.0016803400454344412, -0.0019623919768859415, -0.0022227920394416534, 
    -0.002460137153848926, -0.0026732959026050398, -0.0028614355289683828, 
    -0.0030240449267380171, -0.0031609430455996524, -0.0032722751000768538, 
    -0.0033585036715905172, -0.0034203877481008829, -0.0034589540442413547, 
    -0.0034754628711373466, -0.003471369725678566, -0.0034482874576069675, 
    -0.0034079503949839031, -0.0033521788183999311, -0.0032828509820913691, 
    -0.0032018757871624124, -0.0031111696908009403, -0.003012632020315487, 
    -0.0029081336673228882, -0.0027994956163254698, -0.0026884702092458256, 
    -0.0025767161759996686, -0.0024657694392623448, -0.0023570111697741583, 
    -0.0022516326917585748, -0.0021506010561881655, -0.0020546367470864863, 
    -0.0019642015815628912, -0.0018795040414221419, -0.0018005227181698219, 
    -0.0017270466882275458, -0.001658730127066919, -0.0015951532078040216, 
    -0.0015358826283364334, -0.0014805167891687168, -0.0014287250258360699, 
    -0.0013802686938486541, -0.0013350140750699414, -0.0012929267082464595, 
    -0.0012540619019870934, -0.001218550220869144, -0.0011865752305419382, 
    -0.0011583541954063054, -0.0011341225033979457, -0.0011141267781856136, 
    -0.0010986202575276266, -0.0010878619015455189, -0.0010821246112167416, 
    -0.0010816959632083899, -0.0010868773861035658, -0.0010979835662641804, 
    -0.0011153308293740118, -0.0011392214467271337, -0.0011699200656553764, 
    -0.0012076261003466184, -0.0012524390786915296, -0.0013043259227785865, 
    -0.0013630880954338372, -0.0014283348113465137, -0.0014994698299297577, 
    -0.0015756924374183397, -0.0016560161095417263, -0.0017392994244498779, 
    -0.0018242900891629601, -0.0019096752563172253, -0.0019941271393126223, 
    -0.0020763525562263372, -0.0021551215465720501, -0.0022292991192111636, 
    -0.0022978561892823381, -0.0023598783399226917, -0.0024145685475681316, 
    -0.0024612469139795754, -0.0024993495743095471, -0.0025284373936939886, 
    -0.0025481977751128787, -0.0025584594911453526, -0.0025592084797635018, 
    -0.002550604686570257, -0.0025329972066495091, -0.0025069312918717507, 
    -0.0024731530395859578, -0.0024326001007812193, -0.0023863850519542256, 
    -0.002335775520230616, -0.0022821656094877988, -0.0022270450261149067, 
    -0.0021719626901021095, -0.0021184786956792308, -0.0020681117515890949, 
    -0.002022279361634704, -0.0019822325857155928, -0.0019489991117576568, 
    -0.0019233336051696494, -0.0019056934808959652, -0.0018962260790578896, 
    -0.0018947801628921503, -0.0019009222102625615, -0.00191397464450358, 
    -0.0019330543107975101, -0.0019571217420762902, -0.0019850244005881661, 
    -0.0020155496056171989, -0.0020474680501440701, -0.0020795857827712394, 
    -0.0021107980341036783, -0.0021401444766418801, -0.0021668609139160271, 
    -0.0021904200700952033, -0.0022105573574165384, -0.0022272832189462813, 
    -0.0022408757859079332, -0.0022518644362213881, -0.002260993783393131, 
    -0.0022691737858566339, -0.0022774248698289915, -0.0022868221899402449, 
    -0.0022984429557529979, -0.0023133176178768739, -0.0023323934020907707, 
    -0.0023564902557990613, -0.0023862699528623315, -0.0024222088033458867, 
    -0.002464567635986431, -0.0025133684908300678, -0.0025683716290851549, 
    -0.0026290508571174911, -0.0026945831616790924, -0.0027638471271721346, 
    -0.0028354330335430516, -0.0029076784878881608, -0.0029787160538887374, 
    -0.0030465314244694751, -0.0031090305008260105, -0.0031641062279449093, 
    -0.0032097164919559131, -0.0032439474013525832, -0.0032650825817845458, 
    -0.0032716548559814677, -0.0032624790775980183, -0.0032366730567693494, 
    -0.0031936565514942899, -0.0031331403542814939, -0.0030551108750541309, 
    -0.0029598191956168949, -0.0028477689895785364, -0.0027197075535121862, 
    -0.002576608539227484, -0.0024196533805801845, -0.0022502174526405632, 
    -0.0020698503939428079, -0.0018802537294938387, -0.001683256994637599, 
    -0.0014807881206028667, -0.0012748455982427994, -0.0010674666592134564, 
    -0.00086069141629452101, -0.00065653152774849976, 
    -0.00045693219072976489, -0.00026373910730707439, 
    -7.8660658928327791e-05, 9.6762487251466842e-05, 0.00026118955370010914, 
    0.00041351154037379246, 0.00055287179876370961, 0.00067869545427958334, 
    0.000790702412673396, 0.00088891710631774641, 0.00097366403874080652, 
    0.0010455530009548543, 0.0011054573354739991, 0.0011544716289347277, 
    0.0011938697322498313, 0.0012250469600381371, 0.0012494618503693109, 
    0.0012685734639478314, 0.0012837859025272866, 0.0012963890515877076, 
    0.0013075055804198158, 0.0013180585034455784, 0.001328737197849889, 
    0.0013399907556751489, 0.0013520254295555111, 0.0013648221303016303, 
    0.001378152662196917, 0.0013916078368187933, 0.0014046252893798095, 
    0.0014165170203800249, 0.0014265012167707604, 0.0014337338273888263, 
    0.0014373409083147585, 0.0014364504257648938, 0.0014302178195656902, 
    0.0014178550696409842, 0.0013986576729437461, 0.0013720301308424057, 
    0.0013375013243064988, 0.0012947493566616906, 0.0012436150816740297, 
    0.001184112419873543, 0.0011164380652338678, 0.0010409663088751515, 
    0.0009582422737166136, 0.00086896848206532615, 0.0007739846033763089, 
    0.00067424936022099661, 0.00057082055713662512, 0.00046483554713236267, 
    0.00035748421631244103, 0.00024999385697792537, 0.00014360857557854499, 
    3.9581316007600525e-05, -6.0835474285676782e-05, -0.00015639820348450927, 
    -0.00024588449479212386, -0.00032811429160439103, 
    -0.00040197709870750894, -0.00046645476601373523, -0.0005206419842296783, 
    -0.00056376174177301592, -0.00059516818014298156, 
    -0.00061435248955805195, -0.00062093859640839915, 
    -0.00061468109438458951, -0.00059546249431074159, 
    -0.00056329369577088305, -0.0005183134354295022, -0.00046078745758078093, 
    -0.00039110210667232299, -0.00030976025947548018, 
    -0.00021736142761815042, -0.00011458301582106388, 
    -2.1575990244227568e-06, 0.00011914794670859108, 0.00024854802686909128, 
    0.00038524724930186932, 0.00052844951641596702, 0.00067736195168480943, 
    0.00083118366271330306, 0.00098909765227199681, 0.0011502528620219487, 
    0.0013137447280872738, 0.0014785937864871561, 0.001643726558854175, 
    0.0018079634077559923, 0.001970025985894493, 0.0021285491025250297, 
    0.0022821162571369769, 0.0024292916816835669, 0.0025686605368953948, 
    0.0026988699027420213, 0.0028186612044808577, 0.0029269009417049784, 
    0.003022603764360057, 0.0031049563193161793, 0.0031733279030061001, 
    0.0032272854823842687, 0.0032665919012434862, 0.0032912036906291536, 
    0.0033012596490359855, 0.0032970586755956019, 0.0032790355139917194, 
    0.0032477255896311676, 0.0032037357588098098, 0.0031477121810813144, 
    0.0030803127335155694, 0.003002189904167298, 0.0029139827221473995, 
    0.0028163168940155796, 0.0027098105123163963, 0.0025950798434128076, 
    0.0024727490766506014, 0.0023434535528722737, 0.002207837350982123, 
    0.0020665506565298837, 0.001920229640434402, 0.0017694808306792707, 
    0.0016148624186535184, 0.0014568710685889507, 0.0012959378319417252, 
    0.0011324355915283222, 0.00096668655626901481, 0.00079898826772267556, 
    0.00062963064203314654, 0.00045892327293218192, 0.00028721685953454019, 
    0.00011492423588729817, -5.7466586177342229e-05, -0.00022938573023694212, 
    -0.00040017696695637708, -0.00056911002865532242, 
    -0.00073539642592026382, -0.00089821087885459889, -0.0010567219068195717, 
    -0.0012101246613855621, -0.0013576745834161931, -0.0014987259406647269, 
    -0.0016327658223948629, -0.0017594403113633879, -0.0018785752713053176, 
    -0.0019901846219432984, -0.0020944633588194771, -0.0021917752662106212, 
    -0.0022826296829086983, -0.0023676518841910838, -0.0024475534433051529, 
    -0.0025230978351214357, -0.002595076875744061, -0.0026642874700923266, 
    -0.0027315172405707952, -0.0027975336223142792, -0.0028630675211126395, 
    -0.0029288078550623567, -0.0029953825752703066, -0.0030633489435005685, 
    -0.003133186730075726, -0.0032052877950062035, -0.0032799559684352606, 
    -0.0033574005525524985, -0.0034377347423876414, -0.0035209686614261289, 
    -0.0036070040362282197, -0.0036956332528981597, -0.003786537651447272, 
    -0.0038793015506785886, -0.0039734243649477193, -0.0040683447489651935, 
    -0.0041634634036653772, -0.0042581633712612593, -0.004351826081978016, 
    -0.0044438321773742386, -0.0045335612383636641, -0.0046203741095842688, 
    -0.0047036001924016342, -0.00478252242202825, -0.0048563614881415905, 
    -0.0049242737610986458, -0.0049853551900805697, -0.0050386468798360347, 
    -0.0050831476239227092, -0.0051178294057477357, -0.0051416569841303775, 
    -0.0051536113305731294, -0.0051527235844216349, -0.0051381097883546048, 
    -0.0051090104178053404, -0.0050648327030772822, -0.0050051954262841378, 
    -0.0049299593494977409, -0.0048392597943560031, -0.0047335116123009367, 
    -0.0046134098309802514, -0.0044799060522613008, -0.0043341826827067208, 
    -0.0041776044043812964, -0.0040116758540927376, -0.0038379876775248897, 
    -0.0036581649104845551, -0.0034738165933038932, -0.0032864917073389464, 
    -0.0030976298175432698, -0.0029085276265317537, -0.0027203050893624256, 
    -0.002533878775623099, -0.0023499441568132374, -0.0021689613206639742, 
    -0.0019911609828229884, -0.0018165480526741351, -0.0016449259111959188, 
    -0.0014759273092388072, -0.0013090497870206226, -0.0011437020452940438, 
    -0.00097924408612830869, -0.00081503555589901126, 
    -0.00065046043670431383, -0.00048495360207815994, 
    -0.00031801137410575922, -0.00014919286841286398, 2.1881020424076644e-05, 
    0.00019553414305837735, 0.00037203237514802105, 0.00055158772387455381, 
    0.00073434190230856782, 0.00092035670309226149, 0.0011095907934861693, 
    0.0013018786848781351, 0.0014969062501784772, 0.0016941873623706957, 
    0.0018930502271723155, 0.0020926323417076237, 0.0022918839526774033, 
    0.0024895847557254622, 0.0026843696706085195, 0.0028747652710985803, 
    0.0030592310205545315, 0.0032362046874747528, 0.0034041485821863587, 
    0.0035616014516963094, 0.003707216924320033, 0.0038398092372950582, 
    0.003958389241363755, 0.004062189120399246, 0.0041506866936711958, 
    0.0042236147119330946, 0.0042809640198776186, 0.0043229811596068269, 
    0.004350156841120661, 0.004363216545491681, 0.0043631004643945905, 
    0.0043509532665507444, 0.0043281031597979403, 0.0042960386289242541, 
    0.0042563786423848709, 0.0042108399777436457, 0.0041611850526304655, 
    0.0041091787372535635, 0.0040565293998990719, 0.004004839614687475, 
    0.003955562828572943, 0.0039099586300113381, 0.0038690683508933637, 
    0.0038336946534822912, 0.0038043908651708268, 0.0037814582183546535, 
    0.0037649524207858608, 0.0037546984022177035, 0.0037503047351183571, 
    0.0037511989779291516, 0.0037566578315162869, 0.0037658457933127652, 
    0.0037778634913045771, 0.0037917850857981401, 0.0038067067832418455, 
    0.0038217855248363088, 0.0038362736989459461, 0.0038495478145597613, 
    0.0038611258048683117, 0.0038706748473459856, 0.0038780114134827292, 
    0.0038830892539092909, 0.0038859799885908263, 0.0038868526588044855, 
    0.0038859468304322433, 0.0038835519562366787, 0.0038799863735796223, 
    0.0038755712154914706, 0.0038706163703374585, 0.0038653980536081196, 
    0.0038601446989629546, 0.0038550216097958624, 0.0038501149394228364, 
    0.0038454376214360642, 0.0038409331818644006, 0.0038364880909105628, 
    0.0038319499171720209, 0.0038271576764117984, 0.0038219640894030567, 
    0.0038162606933834281, 0.0038099955848926994, 0.0038031846020382233, 
    0.0037959212086279394, 0.0037883680403522552, 0.0037807558337643486, 
    0.0037733633556379306, 0.0037664931267150535, 0.0037604511745289015, 
    0.0037555161780066931, 0.0037519233799840701, 0.0037498479320199054, 
    0.0037493951146185026, 0.0037506047248170955, 0.0037534558476072597, 
    0.0037578923396701831, 0.0037638342617868246, 0.0037712072338081941, 
    0.0037799617531005547, 0.0037900972607975208, 0.0038016777432467097, 
    0.0038148534153089192, 0.003829877881828544, 0.0038471172033179551, 
    0.0038670571348236671, 0.003890306603087079, 0.0039175951139854941, 
    0.0039497552333105836, 0.0039877065903888755, 0.0040324210127682036, 
    0.0040848844902787416, 0.0041460471330274024, 0.0042167748320154335, 
    0.004297803685111793, 0.0043897011913338517, 0.0044928377931836103, 
    0.0046073793936820895, 0.0047332889162245836, 0.0048703443659522672, 
    0.0050181619913340064, 0.005176231575933189, 0.0053439412183216625, 
    0.0055206129109327453, 0.0057055195401656631, 0.0058979065761274457, 
    0.0060969992261017646, 0.0063020062644765463, 0.0065121168081954759, 
    0.0067264957616972989, 0.006944271169676562, 0.0071645291151262863, 
    0.0073863068053925691, 0.0076085781268499407, 0.0078302419581140099, 
    0.0080501089897463875, 0.0082668787808403282, 0.0084791348174856791, 
    0.0086853298932656284, 0.0088837788723137908, 0.0090726641943809135, 
    0.0092500534064236008, 0.0094139182954834279, 0.0095621675545900821, 
    0.0096926870389801439, 0.0098033888746929046, 0.0098922571233542363, 
    0.0099574008942129137, 0.0099970961350882761, 0.010009832371612501, 
    0.0099943459453897127, 0.0099496482481631343, 0.009875047759916997, 
    0.0097701599199567328, 0.0096349105339842873, 0.0094695337778209921, 
    0.0092745659974492779, 0.0090508377461179443, 0.0087994630251438215, 
    0.0085218302100090459, 0.0082195910088836595, 0.0078946492826010937, 
    0.0075491593624754522, 0.007185510928117418, 0.0068063220743693701, 
    0.0064144271395086758, 0.0060128606602570115, 0.0056048294902726328, 
    0.0051936857326511238, 0.0047828825815696141, 0.0043759255721878415, 
    0.0039763126997210217, 0.0035874676239863439, 0.0032126678740397843, 
    0.002854971136932971, 0.0025171528968249098, 0.0022016452419809447, 
    0.0019104942453571729, 0.0016453339536327855, 0.0014073725646390695, 
    0.0011974072066679082, 0.001015858774533228, 0.00086282557572334032, 
    0.00073813756134947334, 0.00064141547854351297, 0.00057213289753118863, 
    0.00052966536063498164, 0.00051333082714695856, 0.00052242364397913688, 
    0.0005562424569184565, 0.00061411651370831216, 0.00069541893033564766, 
    0.00079957365875357007, 0.00092604618074224, 0.001074314700115076, 
    0.0012438320823161951, 0.0014339716262523436, 0.0016439694036949324, 
    0.0018728784097445735, 0.0021195264448259843, 0.0023824927544667334, 
    0.0026600990026674747, 0.0029504151715376049, 0.0032512846954533105, 
    0.0035603609782233598, 0.0038751552088348881, 0.0041930921682498436, 
    0.0045115720355257379, 0.0048280203391083505, 0.005139938532310517, 
    0.0054449410898314418, 0.0057407973438201683, 0.0060254665971153391, 
    0.0062971193217639197, 0.0065541544479231807, 0.006795198814253227, 
    0.007019091404879144, 0.0072248544698393768, 0.0074116547030255199, 
    0.0075787646175056993, 0.0077255338238403394, 0.0078513735760036927, 
    0.0079557647150580828, 0.0080382782299688871, 0.0080986101890819749, 
    0.008136619097237641, 0.0081523661766411508, 0.0081461505462984782, 
    0.0081185383486008077, 0.008070378999781096, 0.0080028106707810027, 
    0.0079172447791769959, 0.0078153479164107306, 0.0076990058513529188, 
    0.0075702725135599978, 0.0074313209755635032, 0.007284379386404004, 
    0.0071316789641459131, 0.0069753978925299852, 0.0068176136971440007, 
    0.0066602554533329063, 0.00650506859794313, 0.0063535853599568232, 
    0.0062071022140185225, 0.0060666749575389867, 0.0059331157083725343, 
    0.0058070130070205558, 0.0056887610825528305, 0.0055785879005408757, 
    0.0054766009336853485, 0.0053828239784398926, 0.0052972306122089155, 
    0.0052197731334739069, 0.0051503930536388205, 0.0050890286696817152, 
    0.0050356104069031555, 0.0049900562315235274, 0.0049522603853297698, 
    0.0049220711243215471, 0.0048992715641316166, 0.0048835543691130856, 
    0.004874494602858292, 0.0048715310385544514, 0.0048739532981273937, 
    0.0048809095573668932, 0.0048914354586012346, 0.0049044807930491074, 
    0.004918957873483067, 0.0049337748723306939, 0.0049478615805273211, 
    0.0049601862819047609, 0.004969758408862668, 0.004975629441094441, 
    0.004976892593659743, 0.0049726864454669797, 0.0049622035124289501, 
    0.0049447000729098663, 0.0049195099428833737, 0.0048860635009803158, 
    0.0048439052500736544, 0.0047927075067695146, 0.0047322864367688238, 
    0.0046626086608792146, 0.0045837893109049108, 0.0044960810523712183, 
    0.0043998510282687959, 0.0042955586096075507, 0.0041837167871761199, 
    0.0040648572149508868, 0.0039394833559063249, 0.0038080324324547559, 
    0.003670830336648387, 0.0035280422350296393, 0.0033796413687338643, 
    0.003225375939217073, 0.0030647535993660268, 0.002897045481564422, 
    0.0027213078027093556, 0.0025364148139718884, 0.0023410984517493049, 
    0.0021339984203798631, 0.0019137069967767408, 0.0016788195184013022, 
    0.0014279780411389329, 0.0011599188584641212, 0.00087351634798338361, 
    0.00056783112986363014, 0.00024215772512606499, -0.00010392800859460564, 
    -0.00047052113917495905, -0.00085733991246488505, -0.0012636936073332657, 
    -0.001688461798482204, -0.0021300807020578822, -0.0025865536358843648, 
    -0.0030554754331985623, -0.0035340780112895673, -0.00401928574315663, 
    -0.0045077850524318473, -0.0049961050921402987, -0.0054807076102430241, 
    -0.0059580751354775963, -0.0064247899839150963, -0.0068776201143739791, 
    -0.0073135862544816332, -0.0077300283274986505, -0.0081246542125907387, 
    -0.0084955743333456103, -0.0088413219458393401, -0.0091608763042972143, 
    -0.009453659476430008, -0.00971953387673446, -0.0099587789625790318, 
    -0.01017206205761239, -0.010360383421081717, -0.010525009218786985, 
    -0.010667406872372521, -0.010789170237424902, -0.010891953983130613, 
    -0.010977420938721017, -0.011047191094396022, -0.011102805104563105, 
    -0.011145683429298276, -0.011177103596984405, -0.011198174263434158, 
    -0.011209824039381989, -0.01121278852461538, -0.011207611746825915, 
    -0.011194651477919294, -0.011174097239205847, -0.011145995250585751, 
    -0.011110281511238563, -0.011066821926779092, -0.011015460666288049, 
    -0.010956073976712085, -0.010888615390177327, -0.010813154415475069, 
    -0.010729917096809207, -0.010639308473777682, -0.010541930044498807, 
    -0.010438584308715845, -0.010330281876568925, -0.010218234180555515, 
    -0.010103843726582908, -0.0099886865462612794, -0.0098744836899795976, 
    -0.0097630733079446599, -0.0096563665139945843, -0.0095563051921563578, 
    -0.0094648140229758593, -0.0093837492857383777, -0.0093148531873568381, 
    -0.0092597100869598152, -0.0092197065444769456, -0.0091960014564438051, 
    -0.0091894936031391358, -0.0092007929447443081, -0.0092301908967633052, 
    -0.0092776414380945776, -0.0093427396605486844, -0.0094247244065984986, 
    -0.0095224740503150693, -0.00963453312820595, -0.0097591494204627739, 
    -0.0098943130259183058, -0.010037822803073674, -0.010187345099713375, 
    -0.010340487929190388, -0.010494865459839568, -0.010648174777049657, 
    -0.010798247162068493, -0.010943095574601236, -0.011080947261020773, 
    -0.011210271616662888, -0.01132977960015381, -0.011438435726982294, 
    -0.011535441867565841, -0.011620227143578868, -0.011692434411301569, 
    -0.011751889810875944, -0.011798583002433203, -0.011832627809242534, 
    -0.011854218106742359, -0.011863583652221111, -0.011860949715416579, 
    -0.01184649734523697, -0.011820334405537538, -0.011782488304186611, 
    -0.011732903733507258, -0.011671452159773587, -0.011597955891089995, 
    -0.011512212699383425, -0.011414015989049236, -0.011303185729666782, 
    -0.011179579643593415, -0.011043111633892528, -0.010893772683244757, 
    -0.010731637361870586, -0.010556870687609479, -0.010369735292876745, 
    -0.010170592536003397, -0.0099598899191891133, -0.0097381421548292605, 
    -0.009505907454984348, -0.0092637546805394034, -0.0090122225070343766, 
    -0.0087517912777239654, -0.008482853629075332, -0.0082057010706701912, 
    -0.0079205181125020421, -0.0076273944401322128, -0.0073263425744093573, 
    -0.007017318460751867, -0.0067002558769914591, -0.0063750846528263811, 
    -0.0060417601659341199, -0.0057002747450064393, -0.0053506664698431553, 
    -0.0049930290068963146, -0.0046274995927979966, -0.0042542561427441174, 
    -0.0038735047037255182, -0.0034854749635451713, -0.0030904151913372802, 
    -0.0026886050053935889, -0.0022803675790258942, -0.0018660992769022704, 
    -0.0014463086879050496, -0.0010216567826691714, -0.0005930062937177697, 
    -0.0001614644020881292, 0.0002715934011381278, 0.00070450898768598092, 
    0.0011353480659916711, 0.0015619188320608536, 0.0019818157984674476, 
    0.0023924625015308044, 0.0027911662592709045, 0.0031751600203588828, 
    0.0035416370699895652, 0.0038877872708598742, 0.0042108275425335974, 
    0.0045080564092721794, 0.0047768916834057314, 0.0050149405394262934, 
    0.0052200523494143839, 0.0053903822923133853, 0.005524444117426832, 
    0.005621156630228945, 0.0056798658087552061, 0.0057003564232163345, 
    0.0056828328758631646, 0.0056278963296161923, 0.0055365197336151193, 
    0.0054100025809908428, 0.0052499388386137869, 0.005058153633927147, 
    0.0048366524187544663, 0.0045875565921826931, 0.0043130439689203085, 
    0.0040152896582298881, 0.0036964296691110589, 0.0033585370787314042, 
    0.00300362027823106, 0.0026336380242301932, 0.0022505303665788451, 
    0.0018562553307161535, 0.0014528350670751596, 0.0010423922827702643, 
    0.00062717518623668568, 0.00020958488377176634, -0.0002078265905695756, 
    -0.00062235208315347017, -0.0010311488992597296, -0.0014312552758199884, 
    -0.0018196283598794672, -0.002193185813922376, -0.0025488534462297166, 
    -0.0028836197583894697, -0.0031945962804673764, -0.0034790825048805316, 
    -0.0037346313036597605, -0.0039591055254755789, -0.0041507390086151404, 
    -0.0043081857380059003, -0.0044305610779573189, -0.0045174615426330066, 
    -0.0045689785540537712, -0.0045856962379931792, -0.0045686670582135592, 
    -0.0045193725104385966, -0.0044396637941926725, -0.0043316892262449435, 
    -0.0041977966891805106, -0.0040404382398279938, -0.0038620606443757134, 
    -0.0036650309882094788, -0.0034515617642333612, -0.0032236950085808981, 
    -0.0029833158460746477, -0.0027321881813418144, -0.0024720048675367836, 
    -0.0022044459430040175, -0.001931223085439987, -0.0016541165201123013, 
    -0.0013749823100979513, -0.0010957542221384786, -0.00081842733157541344, 
    -0.0005450400974280706, -0.00027763532988026615, -1.8223296640820406e-05, 
    0.00023127109176003074, 0.00046907216314846561, 0.00069362864472539683, 
    0.00090367003283789351, 0.001098275684884697, 0.0012769273194466976, 
    0.0014395389413244305, 0.0015864653324322014, 0.0017184816548460905, 
    0.0018367391164350938, 0.0019426911185349541, 0.0020380156530652406, 
    0.0021245189442094998, 0.0022040523144831372, 0.0022784338138652225, 
    0.0023493736786434913, 0.0024184253351007311, 0.002486934455673385, 
    0.0025560113321646933, 0.0026265164960244409, 0.0026990428502203321, 
    0.0027739171257051597, 0.0028511970447607144, 0.0029306792596249451, 
    0.0030119190131339627, 0.0030942561581251641, 0.0031768593295558628, 
    0.0032587746524037173, 0.0033389914471431054, 0.0034164999835927553, 
    0.0034903536768047406, 0.0035597289367489929, 0.0036239664793929665, 
    0.0036826057939803904, 0.0037354066737884314, 0.0037823565149447168, 
    0.0038236835921920641, 0.0038598633184258003, 0.0038916283550767166, 
    0.0039199683904284433, 0.0039461076299509385, 0.0039714867860975306, 
    0.0039977166811130393, 0.0040265257039755649, 0.0040596999898262895, 
    0.0040990111660806931, 0.0041461387689663764, 0.0042025913588699297, 
    0.004269628359870636, 0.0043481902365093382, 0.004438849097533823, 
    0.0045417685760791712, 0.0046567309703218927, 0.0047831611200583974, 
    0.0049201914551198498, 0.0050667275328859862, 0.0052215241950248183, 
    0.0053832467873825458, 0.005550542757143488, 0.0057220966597653061, 
    0.0058966708067717992, 0.00607314813273042, 0.0062505507951147081, 
    0.0064280487610042063, 0.0066049598231996617, 0.0067807227380739079, 
    0.0069548608122677429, 0.0071269256430736066, 0.0072964570389746856, 
    0.0074629113025631187, 0.007625619204876876, 0.0077837350311569485, 
    0.0079362167494679801, 0.0080818134847722347, 0.0082190848427636659, 
    0.0083464171419940555, 0.0084620594027398771, 0.0085641534572235469, 
    0.0086507788132512663, 0.0087199839644315092, 0.0087698437976204413, 
    0.0087985164258492787, 0.0088043141399537488, 0.008785780413615012, 
    0.0087417588650389455, 0.008671460087909472, 0.0085745003176227984, 
    0.0084509396798297873, 0.0083012913273227355, 0.0081265110601719658, 
    0.0079279668735229656, 0.0077073858546482755, 0.0074667904741046271, 
    0.0072084288672930024, 0.0069346993446347208, 0.0066480809602101187, 
    0.0063510713072434935, 0.0060461216206716987, 0.0057355817884513112, 
    0.0054216460510539792, 0.0051062978303430956, 0.0047912676477841988, 
    0.0044779887299489143, 0.0041675493185065523, 0.0038606791599462985, 
    0.0035577512544194361, 0.0032588008943310797, 0.002963580700030605, 
    0.0026716117833900286, 0.002382255514062404, 0.0020947823119420212, 
    0.0018084211896732475, 0.0015224088065438918, 0.0012360218542802827, 
    0.00094859851866342648, 0.00065956582257203629, 0.0003684593814765974, 
    7.4938922520784271e-05, -0.00022119297142063736, -0.00051999015041246971, 
    -0.00082137247571500299, -0.0011251486978578955, -0.0014310375780651908, 
    -0.0017386976039020358, -0.0020477423807715479, -0.0023577672081372299, 
    -0.002668358336146935, -0.0029791114268779176, -0.0032896252475265223, 
    -0.0035995106844006826, -0.0039083798876514506, -0.0042158342044281419, 
    -0.0045214459862371161, -0.0048247453128659763, -0.0051251894598319482, 
    -0.0054221601642186947, -0.0057149369431622396, -0.0060027118287384329, 
    -0.0062845916850310431, -0.0065596311002496018, -0.0068268548449869184, 
    -0.007085290026450356, -0.0073339854891867349, -0.0075720114456519589, 
    -0.0077984819252537039, -0.0080125566034558067, -0.0082134737808437375, 
    -0.0084005698629026331, -0.0085733280446921561, -0.0087314231839849803, 
    -0.0088747866737709843, -0.0090036425595094987, -0.009118553364065465, 
    -0.0092204231724223751, -0.0093104882709455893, -0.0093902707633260283, 
    -0.0094615180391410883, -0.0095261211672065284, -0.0095860452292712388, 
    -0.0096432454866372166, -0.0096995994173467055, -0.009756851477301022, 
    -0.0098165643643094973, -0.0098801052068350267, -0.0099486423509533069, 
    -0.010023160387143189, -0.010104485983495629, -0.010193336011048574, 
    -0.010290358731735762, -0.010396182456776362, -0.010511432678968903, 
    -0.010636753371475141, -0.010772802299575258, -0.010920240502679672, 
    -0.011079701977734361, -0.011251757455481542, -0.011436877077725919, 
    -0.011635390638687477, -0.0118474546209328, -0.012073015262082726, 
    -0.012311800538519522, -0.012563304537218356, -0.012826797013519124, 
    -0.013101333414035366, -0.01338576422352623, -0.013678760192254009, 
    -0.013978821543974403, -0.014284294034696079, -0.01459337912936704, 
    -0.014904126716195799, -0.015214436151859911, -0.015522053623978255, 
    -0.015824573003405007, -0.016119435313466438, -0.016403954648653588, 
    -0.016675332749103485, -0.016930709732125619, -0.017167215234329722, 
    -0.017382015979624882, -0.017572377015921611, -0.017735718238798756, 
    -0.017869655173025144, -0.017972068722865654, -0.018041152464171199, 
    -0.018075474369338856, -0.018074030727854636, -0.018036285641200803, 
    -0.017962194486061907, -0.017852203859242199, -0.017707225348082823, 
    -0.017528580713368463, -0.017317931398463625, -0.017077200632568616, 
    -0.01680847836476668, -0.016513959738977346, -0.016195872207059304, 
    -0.015856427298342791, -0.015497783695647572, -0.015122033288615694, 
    -0.014731208827310511, -0.014327285950476575, -0.013912212262956499, 
    -0.013487940003507819, -0.013056460986838022, -0.012619844097034712, 
    -0.012180256837215665, -0.011740001233040627, -0.011301512359317525, 
    -0.010867335669158072, -0.010440084287192505, -0.010022381446734752, 
    -0.0096167600262618419, -0.0092255928786151228, -0.0088510020202128593, 
    -0.0084948150160030628, -0.0081585174761739498, -0.0078432312597554125, 
    -0.0075497123470060316, -0.0072783477058048504, -0.0070291734420250872, 
    -0.006801887916469576, -0.0065958821774837551, -0.0064102479723543541, 
    -0.0062438153990755458, -0.0060951762773980168, -0.0059627093426680242, 
    -0.0058445996326832199, -0.0057388643470185127, -0.0056433719878432823, 
    -0.0055558791115091558, -0.0054740567176302978, -0.0053955444074501799, 
    -0.0053180050777442839, -0.0052391841739375033, -0.0051569691489902723, 
    -0.0050694393244149673, -0.0049749088915536201, -0.0048719587964724895, 
    -0.0047594503039148969, -0.0046365416808625826, -0.0045026639168055113, 
    -0.0043575011352474779, -0.0042009542314245443, -0.0040331143199593437, 
    -0.0038542350414264635, -0.0036647371120317367, -0.0034651979406304639, 
    -0.003256366550384822, -0.0030391578908826747, -0.0028146693901310721, 
    -0.0025841725159962401, -0.0023491081502297621, -0.0021110582990681945, 
    -0.0018717050678137069, -0.0016328082050590107, -0.0013961408097568314, 
    -0.0011634351027508922, -0.00093633036058939989, -0.00071631449366863344, 
    -0.00050468794092483498, -0.00030252559154572169, 
    -0.00011067224919445091, 7.0248269632673362e-05, 0.00023977864412929434, 
    0.00039758942534252818, 0.00054340775229878401, 0.00067695902582969275, 
    0.00079790712139560173, 0.00090584818533227492, 0.0010003210862848152, 
    0.0010808658688827703, 0.0011470801479993758, 0.001198701643492723, 
    0.0012356552036507629, 0.0012581342240461616, 0.0012666298563246338, 
    0.0012619597667744922, 0.0012452707966802503, 0.0012180320171310379, 
    0.0011820074825908021, 0.0011391979672987951, 0.00109177993616666, 
    0.0010420128794810292, 0.00099213446299447174, 0.00094423649111394789, 
    0.00090016842548398118, 0.00086144815068151881, 0.00082918097459400045, 
    0.00080404580238422002, 0.00078626680550954718, 0.00077561989956689077, 
    0.000771461385787832, 0.00077277539480237532, 0.00077825743440399224, 
    0.00078640672610024104, 0.00079563830972560908, 0.00080441369716351824, 
    0.00081135484543629478, 0.00081536079531945482, 0.00081566357997564249, 
    0.00081190317015919261, 0.00080413568709213719, 0.00079282699259891577, 
    0.00077880097290530651, 0.00076314870025974576, 0.00074714709237389508, 
    0.00073216155748778299, 0.00071958544568549157, 0.00071076739259947285, 
    0.00070698570349802311, 0.00070940580449787996, 0.00071905528365810581, 
    0.00073678239721567578, 0.00076324705404321315, 0.00079890582737773309, 
    0.00084401217223371069, 0.00089863648389655604, 0.00096268835451121374, 
    0.0010359561123018156, 0.0011181623391998069, 0.0012089926250062487, 
    0.0013081471920077614, 0.0014153788306898001, 0.0015305124254378962, 
    0.0016534539531527738, 0.0017841916286367981, 0.0019227820799619527, 
    0.002069335327610547, 0.0022239808388735851, 0.0023868266867516164, 
    0.0025579058722344618, 0.0027371413591394476, 0.0029243142304536257, 
    0.0031190386063314427, 0.0033207555257444626, 0.0035287371026227468, 
    0.0037421072390422267, 0.0039598472505295423, 0.0041808088630489329, 
    0.0044036987978038344, 0.0046270850078160087, 0.0048493880359095024, 
    0.0050688692708085433, 0.0052836546059749955, 0.0054917398905996451, 
    0.0056910423598670982, 0.0058794500163703214, 0.006054889397717947, 
    0.0062154128721680279, 0.0063592644158937941, 0.0064849566151091841, 
    0.0065913036488791437, 0.0066774416053047457, 0.0067428143030301866, 
    0.0067871421052961662, 0.0068103977382851823, 0.0068127713850271495, 
    0.0067946437350134324, 0.0067565758133247096, 0.0066993171075978158, 
    0.0066237862606792, 0.006531071872305459, 0.0064224256666004578, 
    0.0062992355415116405, 0.0061630328531100172, 0.0060154596674402306, 
    0.0058582559200049608, 0.0056932563040547994, 0.0055223790825093518, 
    0.0053476180842102743, 0.0051710258966375794, 0.0049946892048099451, 
    0.004820712290598027, 0.0046511665266507959, 0.0044880442425391477, 
    0.0043331841988556909, 0.0041881981339420204, 0.0040544053659569146, 
    0.0039327546209551433, 0.0038237591258601894, 0.003727448885218222, 
    0.0036433175819697932, 0.0035703219157033348, 0.0035068843686144741, 
    0.0034509261876862563, 0.0033999135298321452, 0.0033509016600459032, 
    0.0033006133524483092, 0.0032454995295554782, 0.0031818285309868893, 
    0.0031057822549269963, 0.003013568386747034, 0.0029015425508665703, 
    0.0027663149533839549, 0.0026048439501715273, 0.002414513106219705, 
    0.002193167039534265, 0.0019391212352955422, 0.0016511445776624129, 
    0.0013284460182174367, 0.00097062872889265355, 0.00057767049426057037, 
    0.0001499298088343125, -0.00031188414811417306, -0.00080674072228910094, 
    -0.00133330049419275, -0.0018899862314556504, -0.0024750357946783617, 
    -0.0030865540463459913, -0.0037225494466851736, -0.0043809202334848252, 
    -0.0050594009631833746, -0.0057554841975031553, -0.0064663968100351476, 
    -0.007189069034493371, -0.0079201597471028947, -0.008656102047833427, 
    -0.0093931864003268528, -0.010127641143543309, -0.010855712827071746, 
    -0.011573750482727416, -0.012278282329209389, -0.012966084244227388, 
    -0.013634238893375712, -0.014280170434952074, -0.014901680727839145, 
    -0.015496949624065179, -0.016064500871348964, -0.016603191784894066, 
    -0.017112176026320421, -0.017590870407464265, -0.018038939477890557, 
    -0.018456342441524175, -0.018843341359130177, -0.019200588952235975, 
    -0.019529134887476578, -0.019830480510837772, -0.020106555224345315, 
    -0.020359654655314221, -0.020592351733021347, -0.020807372912121896, 
    -0.021007448412038433, -0.021195139648581936, -0.021372731075227545, 
    -0.021542099991248925, -0.021704637423382699, -0.021861244825305381, 
    -0.022012352248473359, -0.022157976376719783, -0.022297834061134628, 
    -0.022431446003413104, -0.022558249856975542, -0.022677676749082692, 
    -0.022789238099124379, -0.022892576585776845, -0.022987489455334725, 
    -0.023073920986487646, -0.023151927937370524, -0.023221672770971244, 
    -0.02328334958860959, -0.023337214031801886, -0.023383620410312059, 
    -0.023423056761310877, -0.023456199408979021, -0.023483964852741124, 
    -0.023507541032852027, -0.023528380809143285, -0.023548179677027988, 
    -0.023568830638250993, -0.023592362671616962, -0.023620863285916307, 
    -0.023656364888250774, -0.02370075950594815, -0.023755659115635569, 
    -0.023822262032876997, -0.023901231376680029, -0.023992565862123887, 
    -0.024095516858680201, -0.02420854710372599, -0.024329368159835864, 
    -0.024454957766419337, -0.024581609119897173, -0.024704985331786212, 
    -0.024820155338639616, -0.02492168064389565, -0.025003729561243741, 
    -0.025060209074011189, -0.025084953341906344, -0.025071904740748479, 
    -0.025015275152662681, -0.024909709999273957, -0.0247504109549961, 
    -0.024533270778608361, -0.024254988930137868, -0.023913154556312825, 
    -0.023506354220562298, -0.023034203113105133, -0.022497349796859613, 
    -0.021897446998693806, -0.021237094404917573, -0.020519753966318485, 
    -0.019749674407531705, -0.018931787851622583, -0.018071640923986668, 
    -0.017175271911394927, -0.01624914733197683, -0.015300062579101601, 
    -0.014335105619692994, -0.013361577463612896, -0.01238692632037173, 
    -0.011418708489546079, -0.010464566925629309, -0.0095321995163303586, 
    -0.008629307774542452, -0.007763561074171841, -0.0069425500644253214, 
    -0.0061736957855176768, -0.0054641872784754577, -0.0048208483401758415, 
    -0.00425002237989721, -0.0037574237458061913, -0.0033479694086043358, 
    -0.0030256748576623907, -0.0027935539347358428, -0.0026535552892419652, 
    -0.0026065402642965309, -0.002652340543690344, -0.002789790445946798, 
    -0.0030167861599453669, -0.0033303722991204895, -0.0037267974134007542, 
    -0.0042016108451188349, -0.004749729763293368, -0.0053655348682615581, 
    -0.006042929344051309, -0.0067754334077201311, -0.0075562455701350621, 
    -0.0083782258491382801, -0.0092338998982851358, -0.01011539313576581, 
    -0.011014404710858346, -0.011922274647492629, -0.01283011752829771, 
    -0.013728958057518783, -0.014609935307727027, -0.015464419419551203, 
    -0.016284129393815353, -0.017061230753987869, -0.017788400024503343, 
    -0.018458865982207039, -0.019066419106528881, -0.019605432310504784, 
    -0.020070781410476343, -0.020457874115411685, -0.020762560013872156, 
    -0.020981218427499834, -0.021110726698816602, -0.021148470639432655, 
    -0.02109238038361156, -0.020941006093656227, -0.020693519940117679, 
    -0.020349817588426505, -0.01991061107373816, -0.01937754721035034, 
    -0.018753325585772702, -0.018041789011902683, -0.017248032599889284, 
    -0.016378366364196213, -0.015440198787819317, -0.014441896242212331, 
    -0.01339252177762418, -0.012301644774928027, -0.011179127474859312, 
    -0.010034926038736226, -0.0088789902411624596, -0.0077210634557266129, 
    -0.0065705259709876009, -0.0054362935320630551, -0.0043266653650865195, 
    -0.0032492292547148319, -0.0022108322567675164, -0.0012175760586420339, 
    -0.00027488839343882106, 0.00061234178480702901, 0.0014397339791355265, 
    0.0022032742793221837, 0.0028992744043615085, 0.003524433656569805, 
    0.004075826062926515, 0.0045510512015471734, 0.0049482729554610524, 
    0.0052662642029593938, 0.0055044955986362819, 0.0056629974912754417, 
    0.0057425286926010644, 0.0057444548822079009, 0.0056707731983014539, 
    0.0055241199038175677, 0.0053077472961486245, 0.0050254551800182779, 
    0.0046815137951358131, 0.0042804497411071665, 0.0038269002519831785, 
    0.0033255014164013485, 0.0027808380442067393, 0.0021974210532397743, 
    0.0015797412633107842, 0.00093238429592396466, 0.00026015814727405918, 
    -0.00043182682480147816, -0.0011379648850962346, -0.0018521665298837082, 
    -0.0025679240872109954, -0.0032784303064660471, -0.0039766472383285009, 
    -0.0046554576855671864, -0.0053078819843478363, -0.0059272241774525926, 
    -0.0065072139680604334, -0.0070423623808023549, -0.0075281758689819461, 
    -0.0079612705960822108, -0.0083395149251009777, -0.0086620325708811757, 
    -0.0089289060870073218, -0.0091410828816153554, -0.0092999619885583574, 
    -0.0094070523713360235, -0.0094637004510197114, -0.0094712155744928559, 
    -0.0094310159441754714, -0.0093449593485701483, -0.0092160696382431549, 
    -0.0090488416246176963, -0.0088492899385292801, -0.0086246040529234982, 
    -0.0083826087640792284, -0.0081311584576423488, -0.0078777451282763967, 
    -0.0076296067369402559, -0.0073937143598172177, -0.0071771003411437856, 
    -0.006986955183590899, -0.0068306041567815804, -0.0067153255519584436, 
    -0.006648388362544856, -0.0066364304381389145, -0.0066855265764143466, 
    -0.0068001653413138873, -0.0069834075995618521, -0.007236393659481667, 
    -0.007558022196920788, -0.0079444814875386013, -0.0083894690787017969, 
    -0.0088836631339748208, -0.0094157722220574065,
  // Fqt-F(4, 0-1999)
    1, 0.99719415632104857, 0.98884452633408215, 0.97515210325167989, 
    0.9564408275378723, 0.93314126002716757, 0.90576979593159157, 
    0.87490512254018016, 0.84116368865939095, 0.8051758260810401, 
    0.76756388553298605, 0.72892339594043143, 0.68980787333073268, 
    0.6507175166983491, 0.61209176173115332, 0.57430538872076331, 
    0.53766772314469047, 0.50242441348383227, 0.4687611878367936, 
    0.43680900951022161, 0.40665015333795046, 0.37832470996445045, 
    0.3518371568361453, 0.32716269747125809, 0.30425314434714235, 
    0.28304224745184386, 0.26345038164518769, 0.24538861695729355, 
    0.22876217307832861, 0.21347331947105957, 0.19942376836603709, 
    0.18651658491047074, 0.17465769459657116, 0.16375700168376806, 
    0.15372920166440654, 0.14449433024381614, 0.13597809518116713, 
    0.12811204853843086, 0.12083362080790436, 0.11408605917465958, 
    0.10781827368764185, 0.1019846290799479, 0.096544656936743412, 
    0.091462727978227257, 0.086707655848307391, 0.082252271332827906, 
    0.078072985526946165, 0.074149336718240283, 0.070463567214134659, 
    0.067000216220641826, 0.063745756529304309, 0.060688259032452202, 
    0.057817097843635833, 0.055122695369743423, 0.0525962878124289, 
    0.050229723126323012, 0.048015284417046319, 0.045945530465301691, 
    0.044013162068097231, 0.042210913549424328, 0.040531471623716016, 
    0.038967425296869952, 0.037511251433715656, 0.036155333587513848, 
    0.034892000033301826, 0.033713579774327811, 0.032612472029984088, 
    0.031581205040291813, 0.03061250600194703, 0.029699352660930298, 
    0.028835038786604213, 0.028013214407725893, 0.027227936057898094, 
    0.026473676211324775, 0.025745335758407626, 0.025038228240073769, 
    0.024348050641047513, 0.023670862219249984, 0.023003058621989779, 
    0.022341358199788934, 0.02168280217319744, 0.021024753929866715, 
    0.020364929790083572, 0.019701409790107271, 0.019032662353807375, 
    0.018357557671769574, 0.01767537239586997, 0.016985788381304358, 
    0.016288878686387419, 0.015585081480512736, 0.014875162935857724, 
    0.014160160523659624, 0.013441309698602775, 0.012719969893190332, 
    0.011997547175824987, 0.011275429381871881, 0.010554938236080417, 
    0.0098373075308812018, 0.0091236781272197951, 0.0084151150362910508, 
    0.0077126344028926735, 0.0070172495845726912, 0.006330014125510347, 
    0.0056520611740501501, 0.0049846417314405268, 0.0043291322380238501, 
    0.0036870197788579184, 0.0030598735342093229, 0.0024492920814533858, 
    0.001856834374301669, 0.0012839560552623109, 0.00073193774916615879, 
    0.00020183751227959186, -0.00030554388276659444, -0.00078967410219805501, 
    -0.0012502777532786072, -0.0016872981727124297, -0.0021008433618809825, 
    -0.0024911136586997064, -0.002858335859370743, -0.0032027011751794799, 
    -0.0035243139917076208, -0.0038231617622576384, -0.0040990915843508152, 
    -0.0043518036811801561, -0.0045808495473599192, -0.0047856357214520195, 
    -0.0049654253657232675, -0.0051193427140146883, -0.0052463832447469634, 
    -0.0053454276266126938, -0.0054152663840098007, -0.0054546414808800577, 
    -0.0054622957781560871, -0.00543703159065598, -0.0053777809055134294, 
    -0.0052836673254279274, -0.0051540675376318497, -0.0049886626405295049, 
    -0.0047874733927070487, -0.0045508920340469085, -0.0042796835103210071, 
    -0.0039749870738880746, -0.0036382879578947354, -0.0032713903290904466, 
    -0.0028763706627721406, -0.0024555296677438963, -0.0020113415081710303, 
    -0.0015464091183541645, -0.0010634328469526764, -0.00056517777367930946, 
    -5.4461164251658721e-05, 0.00046585006554669076, 0.0009928305527135404, 
    0.0015234961683305327, 0.0020547919039332371, 0.0025836011222952148, 
    0.0031067596108754671, 0.0036210967873765766, 0.0041234799967698006, 
    0.0046108803643824543, 0.005080441279639419, 0.0055295422447198686, 
    0.0059558587495942674, 0.0063574124705740864, 0.0067326044678752747, 
    0.0070802507068249958, 0.0073995849924118721, 0.0076902594500907967, 
    0.0079523157889816037, 0.0081861472268423743, 0.00839246459061419, 
    0.0085722609744246486, 0.0087267806695053365, 0.0088574775446921029, 
    0.0089659752235578868, 0.0090539985920669534, 0.0091232966617725564, 
    0.0091755664867794861, 0.0092123687607775437, 0.0092350670543280746, 
    0.0092447788263582548, 0.0092423579747803984, 0.0092283925304582817, 
    0.0092032319744708869, 0.0091670194772981734, 0.0091197316251430682, 
    0.009061216972446183, 0.0089912313364711033, 0.0089094662819689495, 
    0.008815578459198321, 0.0087092119417150685, 0.0085900273378853448, 
    0.008457726318725255, 0.0083120917446515997, 0.0081530171411854872, 
    0.0079805547681681844, 0.0077949571522244595, 0.0075967200605229004, 
    0.0073866222026242878, 0.0071657567790053105, 0.0069355568544313562, 
    0.0066978100862971329, 0.0064546683766818352, 0.0062086479122300912, 
    0.0059626178614756963, 0.0057197778384313397, 0.0054836136073829799, 
    0.0052578382073929751, 0.0050463076145184187, 0.0048529098340406012, 
    0.0046814449257099964, 0.0045354942273955912, 0.0044182772906206508, 
    0.0043325115894532534, 0.0042802822653971815, 0.0042629326705511394, 
    0.0042809718379767624, 0.0043340187529513161, 0.0044207837490942382, 
    0.0045390852399431903, 0.0046859104093325294, 0.0048575083062281149, 
    0.0050495158024392592, 0.0052570993881948889, 0.0054751205880706538, 
    0.0056983081912453486, 0.0059214412741429232, 0.0061395172834756402, 
    0.0063479180177100931, 0.0065425434545539713, 0.0067199247096129452, 
    0.0068772937537021801, 0.0070126233278495018, 0.0071246129699068699, 
    0.0072126417729336855, 0.0072766908814505165, 0.0073172407352413002, 
    0.0073351579642799295, 0.0073315759147042315, 0.0073077947936643689, 
    0.0072651915093348129, 0.0072051559524033519, 0.0071290572654651753, 
    0.0070382201908340807, 0.0069339371328042687, 0.006817481202628867, 
    0.0066901376916376921, 0.0065532287394099486, 0.0064081422478875017, 
    0.0062563461943501873, 0.0060993873580516807, 0.0059388726906766205, 
    0.0057764242649602704, 0.0056136237824107645, 0.0054519396038878289, 
    0.0052926595011539342, 0.0051368198120027376, 0.0049851496755175155, 
    0.004838029960358519, 0.0046954802622110525, 0.0045571571993271174, 
    0.0044223859058423621, 0.0042901884043736044, 0.0041593335682010742, 
    0.0040283879483315492, 0.0038957697138430145, 0.003759804953244743, 
    0.0036187976192534814, 0.0034710933042825733, 0.0033151502806814865, 
    0.0031496046405936622, 0.0029733344264040503, 0.0027855212184235397, 
    0.0025857003901668561, 0.0023738078068415895, 0.0021502119141474174, 
    0.0019157418341781553, 0.0016716945212752782, 0.0014198257609256298, 
    0.0011623219479028684, 0.00090175359183489114, 0.00064099711028769242, 
    0.00038314026258094578, 0.00013137765217095221, -0.00011110808741517379, 
    -0.00034125667814036132, -0.00055622933560575292, 
    -0.00075349084849805404, -0.00093086976550375811, -0.0010866007703068965, 
    -0.0012193523338480676, -0.0013282423504548048, -0.0014128493487218119, 
    -0.0014732111058427184, -0.0015098083759421805, -0.001523536374784648, 
    -0.0015156460361745239, -0.0014876766494575286, -0.0014413705916967517, 
    -0.0013785812513509208, -0.0013011825708993899, -0.0012109957466259192, 
    -0.0011097358763986929, -0.00099897785975640307, -0.00088016088951976411, 
    -0.00075460140627939612, -0.00062352497427057424, 
    -0.00048808958184514361, -0.00034939506252800834, 
    -0.00020848491748884414, -6.6347129669199579e-05, 7.6072719935526911e-05, 
    0.00021784838184787009, 0.00035803745522738586, 0.00049565932791636829, 
    0.00062968822320730571, 0.00075905891508085371, 0.00088269708165202975, 
    0.00099955648704018636, 0.0011086650474864872, 0.0012091666714792821, 
    0.001300354138496349, 0.0013816922869749363, 0.0014528330845344313, 
    0.0015136192185879296, 0.0015640872310987257, 0.0016044771596954769, 
    0.0016352341516375751, 0.0016570043389409093, 0.001670634174746602, 
    0.0016771562502278384, 0.0016777702803986295, 0.0016738179783589218, 
    0.0016667541047004171, 0.0016581143722355141, 0.00164947839673659, 
    0.0016424306744118454, 0.001638516122780815, 0.0016392033258817963, 
    0.0016458437614832067, 0.0016596407215705056, 0.0016816119262112318, 
    0.0017125741798185027, 0.0017531063911171525, 0.0018035310539486183, 
    0.0018638877381180335, 0.0019339163425197241, 0.002013046317942154, 
    0.0021003905209978622, 0.0021947556928997385, 0.002294666345613771, 
    0.0023983976166527185, 0.002504003564244895, 0.0026093605832122899, 
    0.0027121960802348661, 0.0028101273297100097, 0.0029007005828070322, 
    0.0029814498586064522, 0.003049964688364994, 0.0031039771031410269, 
    0.0031414294307966538, 0.0031605404397845758, 0.0031598533075106613, 
    0.0031382680161664966, 0.003095054937897261, 0.0030298603292946251, 
    0.002942695209205808, 0.0028339241075465392, 0.0027042536418692541, 
    0.0025547095048450968, 0.0023866206433807444, 0.0022015933916523546, 
    0.0020014815465184427, 0.001788349191302279, 0.0015644272529655718, 
    0.0013320671967090351, 0.0010936830826696728, 0.00085168829616652768, 
    0.00060843375092830914, 0.00036614769505811571, 0.00012688373541057082, 
    -0.00010751937095083617, -0.00033545529239054832, 
    -0.00055555008436090848, -0.00076663898176855202, -0.0009677458504344272, 
    -0.0011580507361275366, -0.00133686828946315, -0.0015036418179946265, 
    -0.0016579371749545404, -0.0017994443947374488, -0.0019279760846027528, 
    -0.0020434586612940926, -0.002145922263146762, -0.0022354836474124699, 
    -0.0023123284963893938, -0.0023766928588426794, -0.002428848320572699, 
    -0.0024690880184642227, -0.002497719944616499, -0.0025150596478198087, 
    -0.0025214252631474187, -0.0025171341131317395, -0.0025024996846786918, 
    -0.0024778282677559958, -0.0024434175181167524, -0.0023995691880465452, 
    -0.0023466004817070348, -0.002284862074499646, -0.0022147650045415313, 
    -0.0021368045578783056, -0.0020515797771120752, -0.0019597910622779005, 
    -0.0018622362413271802, -0.0017597807611400452, -0.0016533248621284444, 
    -0.001543760241462386, -0.0014319227086344317, -0.0013185392644195276, 
    -0.0012041886546366796, -0.0010892682835676, -0.00097398025886656571, 
    -0.00085834225523695093, -0.00074221254068432578, 
    -0.00062532581194897608, -0.00050734537760440952, 
    -0.00038791730100258244, -0.00026671930191463165, 
    -0.00014350880294158007, -1.815404809678311e-05, 0.00010934334288011918, 
    0.00023884095011068396, 0.00037006183481072053, 0.00050261062807650857, 
    0.00063599317250985976, 0.00076964111060779197, 0.00090294276139816154, 
    0.0010352689862657568, 0.0011660031892938788, 0.0012945630463209348, 
    0.0014204245790275379, 0.001543141073183318, 0.0016623595352527028, 
    0.0017778221975671196, 0.0018893616647361544, 0.0019968730619247701, 
    0.0021002654904829117, 0.002199400188008978, 0.002294023439604958, 
    0.0023837175446454052, 0.0024678806092554573, 0.0025457475535645749, 
    0.0026164302207725134, 0.0026789820435075395, 0.0027324661719586849, 
    0.0027760246631341025, 0.0028089393521996552, 0.0028306834509940503, 
    0.0028409724495279337, 0.0028397794328100527, 0.0028273477321913106, 
    0.0028041814727809019, 0.0027710238007003988, 0.0027288161602417593, 
    0.0026786513543747758, 0.0026217185308467545, 0.0025592402279814939, 
    0.002492406927074641, 0.0024223187202455426, 0.002349926305040332, 
    0.0022759891345397231, 0.0022010528200997921, 0.0021254206365018775, 
    0.0020491558586522018, 0.0019720925565600194, 0.001893860168004185, 
    0.0018139157048555209, 0.0017315853934958272, 0.0016461237486415337, 
    0.0015567713342504231, 0.0014628177197798708, 0.0013636605364205855, 
    0.0012588529332682871, 0.0011481365643999551, 0.0010314584090236711, 
    0.00090896327485588137, 0.00078097466813709343, 0.00064796400746805483, 
    0.00051050598451253461, 0.00036923170734510635, 0.00022478401609457075, 
    7.7783994890442867e-05, -7.1194605069334029e-05, -0.00022163954233285818, 
    -0.00037309984102895123, -0.00052517389772199189, -0.0006774956216837163, 
    -0.0008297141747419098, -0.00098147067042625045, -0.0011323769059034118, 
    -0.0012820031405291967, -0.0014298593647914697, -0.0015753924135509705, 
    -0.0017179794835948869, -0.0018569124665451533, -0.0019914006021064423, 
    -0.0021205622161342879, -0.0022434352930429799, -0.0023590001067018045, 
    -0.0024662139374582457, -0.00256405343762646, -0.0026515605782376104, 
    -0.0027278948072496064, -0.0027923593477906334, -0.0028444447784798251, 
    -0.0028838465520467363, -0.0029104921362486822, -0.0029245561848567424, 
    -0.0029264714058332706, -0.0029169189379910825, -0.0028968122992791183, 
    -0.0028672484978778476, -0.002829440264392621, -0.0027846309075761498, 
    -0.0027340040773869059, -0.0026785959504242226, -0.0026192384394069148, 
    -0.0025565156613947589, -0.0024907649387287951, -0.0024220955958530756, 
    -0.0023504279413305508, -0.0022755552911988665, -0.0021972107804527955, 
    -0.0021151543944873423, -0.0020292556788618979, -0.0019395767536839513, 
    -0.0018464317506871422, -0.0017504230255260106, -0.0016524465759178127, 
    -0.0015536735498382687, -0.00145549551703879, -0.0013594607873198901, 
    -0.0012671883867894323, -0.0011802750677111246, -0.0011001968189798858, 
    -0.0010282021174941359, -0.00096521300674310242, -0.00091173460909218921, 
    -0.00086778247626997332, -0.00083283388483304131, 
    -0.00080581038835174758, -0.00078508692722713681, 
    -0.00076853271589386854, -0.00075358665187332842, 
    -0.00073734825868249825, -0.00071668871118894329, 
    -0.00068837075830674812, -0.0006491764103862365, -0.00059602710552652443, 
    -0.00052608898158005614, -0.00043687190175312646, 
    -0.00032631377752615582, -0.00019285893067914355, 
    -3.5522704958251567e-05, 0.00014605039680709228, 0.00035154073361049794, 
    0.0005799263757350734, 0.00082948362996742285, 0.0010978099798269227, 
    0.0013818736660462902, 0.0016780850738758149, 0.0019823824731015315, 
    0.002290337491242256, 0.0025972538810960497, 0.0028982796234255847, 
    0.0031885072675177598, 0.0034630699332024069, 0.0037172398769172903, 
    0.0039465190007254639, 0.004146726926588724, 0.004314079182554208, 
    0.0044452606132122539, 0.0045374939382588683, 0.0045885972176479967, 
    0.0045970402032163528, 0.0045619809728528211, 0.0044832940419326176, 
    0.004361571251095272, 0.0041981130237193093, 0.0039948845811595655, 
    0.003754452307027627, 0.0034798980598618871, 0.0031747134850093339, 
    0.0028426849425108444, 0.0024877727128407657, 0.0021140040775296867, 
    0.0017253756591798742, 0.0013257755237162715, 0.00091893931312963671, 
    0.00050841939038749357, 9.7565762258870585e-05, -0.00031048342411735865, 
    -0.0007128228895427873, -0.0011068056122757772, -0.0014900749025705084, 
    -0.0018605886705400842, -0.0022166404107348088, -0.0025568681731505862, 
    -0.0028802414796283006, -0.0031860392283780143, -0.0034738170599937545, 
    -0.0037433719734826757, -0.003994715975416817, -0.0042280412893217056, 
    -0.0044437064189712747, -0.0046422090481889906, -0.0048241624616754174, 
    -0.0049902680025560135, -0.0051412822387165947, -0.0052779719262457236, 
    -0.0054010652361508107, -0.0055111997812083632, -0.0056088721853702009, 
    -0.0056943851224277109, -0.0057678247954132053, -0.0058290386543655747, 
    -0.0058776369078176365, -0.0059130136901892096, -0.0059343819593878104, 
    -0.0059408248152142866, -0.0059313472364502396, -0.0059049399888884049, 
    -0.0058606316955622595, -0.0057975409708262973, -0.0057149192427950486, 
    -0.0056121765034101443, -0.005488909269720104, -0.0053449124199774793, 
    -0.0051801958221618519, -0.0049949927404042641, -0.00478977378161222, 
    -0.0045652614407079633, -0.004322444624236749, -0.0040625943072472373, 
    -0.0037872852912846883, -0.0034984087874077871, -0.0031981932856710057, 
    -0.0028892039065605397, -0.0025743346911521019, -0.0022567850975996812, 
    -0.001940005923849744, -0.0016276397294037832, -0.0013234301618336587, 
    -0.0010311279698672574, -0.0007543796944945425, -0.00049661511207761894, 
    -0.00026094475033672216, -5.0059092888541866e-05, 0.00013384787173959238, 
    0.0002891550047802234, 0.00041485855890757895, 0.00051059939071606381, 
    0.00057666813483649431, 0.0006139802795770093, 0.00062403071726616598, 
    0.00060882573303207212, 0.00057080513134777594, 0.00051274674558722891, 
    0.00043765649520480265, 0.00034865656141569467, 0.00024885709467580919, 
    0.00014123580585251669, 2.8526531824199768e-05, -8.687581747111883e-05, 
    -0.00020298089903625691, -0.00031823798290791128, 
    -0.00043155058831572486, -0.00054226788821480512, 
    -0.00065015945293366332, -0.00075537498289587771, 
    -0.00085839675585067153, -0.00095997582310882986, -0.0010610611070570844, 
    -0.0011627144019947173, -0.0012660228556501943, -0.0013720071741523709, 
    -0.0014815340964039068, -0.0015952397777352335, -0.0017134632777737265, 
    -0.0018362043131640601, -0.0019631015169041446, -0.0020934438769261736, 
    -0.0022262224788828335, -0.0023602067785049915, -0.002494053551997168, 
    -0.0026264276663288681, -0.0027561131982411884, -0.0028821107560220724, 
    -0.0030037034053946197, -0.0031204931152081562, -0.0032323989897515629, 
    -0.0033396373208040391, -0.0034426648593240405, -0.0035421051055133414, 
    -0.003638653675030243, -0.0037329824618681203, -0.0038256433859923437, 
    -0.0039169897231335748, -0.0040071143648726234, -0.0040958217941466576, 
    -0.0041826220124790061, -0.0042667640714946177, -0.0043472847604069977, 
    -0.0044230878986860882, -0.0044930274789231651, -0.0045560007865792385, 
    -0.0046110412076476774, -0.0046573949485030925, -0.0046945852988642565, 
    -0.0047224672841842397, -0.0047412454464295841, -0.0047514777844078881, 
    -0.0047540461964299405, -0.0047501050172213677, -0.0047410034573807242, 
    -0.0047281926693457186, -0.0047131358555969607, -0.0046972183537075099, 
    -0.0046816723847687295, -0.0046675277385834716, -0.0046555726436277841, 
    -0.0046463312853719171, -0.0046400584379795882, -0.0046367403799492616, 
    -0.0046361095208513484, -0.0046376670941247842, -0.00464071557580608, 
    -0.0046443972151050577, -0.0046477404659975756, -0.0046497073208816323, 
    -0.0046492435918035245, -0.0046453200138971227, -0.0046369747154279368, 
    -0.0046233506300461438, -0.0046037262207090212, -0.0045775420270850117, 
    -0.0045444135563191762, -0.0045041351192681572, -0.0044566605329761757, 
    -0.0044020637905717126, -0.0043404813076618302, -0.0042720532891186826, 
    -0.0041968610533186321, -0.0041148871917741723, -0.004025991919208916, 
    -0.0039299086515593362, -0.0038262504986137365, -0.0037145278820789212, 
    -0.0035941799428275754, -0.0034646113825755748, -0.0033252312367188378, 
    -0.0031755135262894964, -0.0030150452406954844, -0.0028435849069509728, 
    -0.0026611169171084775, -0.0024678983429621579, -0.0022645060315933264, 
    -0.0020518714568299816, -0.0018313105159935507, -0.0016045390387901559, 
    -0.0013736725889805829, -0.001141209243723725, -0.00090998987295210724, 
    -0.00068314433233024308, -0.00046401585516991038, 
    -0.00025607025169253179, -6.2793777785169285e-05, 0.00011241210016551466, 
    0.00026633983807357569, 0.0003960763137104067, 0.00049908922856620403, 
    0.00057331008364595946, 0.00061718421163323481, 0.00062971698026091682, 
    0.00061049119521951309, 0.00055966733200681995, 0.0004779650455704978, 
    0.00036663053481604437, 0.00022739094397911574, 6.2397930102029093e-05, 
    -0.00012582675274355011, -0.00033445681826066269, 
    -0.00056042504402263019, -0.00080048639799712906, -0.001051287371344, 
    -0.0013094365538849815, -0.0015715801604852546, -0.0018344812690613234, 
    -0.0020950989669695961, -0.0023506730195016006, -0.0025987928707226107, 
    -0.0028374600351071212, -0.0030651304409541119, -0.0032807303423961543, 
    -0.003483647643722429, -0.0036737015700252199, -0.0038510848626277382, 
    -0.0040162969526853533, -0.0041700579059435914, -0.0043132273574395478, 
    -0.0044467260523911771, -0.0045714673301239387, -0.0046883018797445027, 
    -0.0047979865956900404, -0.0049011689420886467, -0.004998393508207721, 
    -0.0050901162479204936, -0.0051767334375135273, -0.0052586073860074111, 
    -0.005336094057428061, -0.0054095629516511985, -0.0054794182725641438, 
    -0.0055461107212154406, -0.0056101492641922115, -0.0056720946621225078, 
    -0.0057325521184501231, -0.0057921603652122018, -0.0058515660219602382, 
    -0.0059113970538985303, -0.0059722354495907902, -0.0060345927823755845, 
    -0.0060988959292196604, -0.0061654813234194999, -0.0062345946224730935, 
    -0.0063063976976528661, -0.0063809773349200027, -0.0064583471150013614, 
    -0.0065384368103003311, -0.0066210771432893062, -0.0067059610938886979, 
    -0.0067926053381226993, -0.0068803109740961177, -0.0069681239331988382, 
    -0.0070548165361902209, -0.0071388871354673041, -0.0072185847925518281, 
    -0.0072919581663756236, -0.0073569358736041536, -0.0074114198440762454, 
    -0.0074533912468551797, -0.0074810234836102107, -0.0074927870751395264, 
    -0.0074875398854582637, -0.0074645958541753373, -0.0074237632732671206, 
    -0.0073653499398189486, -0.0072901376598881705, -0.0071993350723357878, 
    -0.007094499621482891, -0.0069774612496777636, -0.0068502303095879626, 
    -0.0067149113697942539, -0.0065736208808917958, -0.0064284140712619351, 
    -0.0062812316763185194, -0.0061338499667300357, -0.0059878539370665368, 
    -0.0058446218512509997, -0.0057053276154247559, -0.0055709523854957062, 
    -0.0054423154379637665, -0.0053201021455861483, -0.0052049003841743409, 
    -0.0050972282223434506, -0.004997547484043365, -0.0049062537929570917, 
    -0.0048236437900729245, -0.0047498667645407338, -0.004684860479766643, 
    -0.0046282845722289342, -0.004579478039924389, -0.0045374249064546925, 
    -0.0045007523538689535, -0.0044677597569578896, -0.0044364821205009385, 
    -0.0044047726615103209, -0.004370407807966761, -0.0043312102583074252, 
    -0.00428516559308893, -0.0042305431318525001, -0.0041660009401969572, 
    -0.0040906831267200627, -0.0040042788174843294, -0.0039070471955384226, 
    -0.0037998167672802534, -0.0036839313832320621, -0.0035611739554584827, 
    -0.003433659273502484, -0.0033037101970206134, -0.0031737310835850624, 
    -0.0030460872335976081, -0.0029229996050445526, -0.0028064712082193702, 
    -0.0026982393604254085, -0.0025997605002352339, -0.0025122100571289608, 
    -0.0024364974099235254, -0.0023732772676269523, -0.0023229406359800515, 
    -0.0022856000273395434, -0.0022610520026828998, -0.0022487325829318038, 
    -0.0022476711637241359, -0.0022564602200556435, -0.0022732419450312924, 
    -0.0022957275949875948, -0.0023212448104802737, -0.0023468042591390198, 
    -0.00236918885646412, -0.0023850343310257184, -0.0023909253496937196, 
    -0.0023834868326235914, -0.0023594796529836826, -0.0023158845650094479, 
    -0.0022499938997733648, -0.0021594929217959818, -0.0020425365382639145, 
    -0.0018978110846833288, -0.0017245872448999363, -0.0015227404821784082, 
    -0.0012927580671353235, -0.0010357186020610266, -0.00075324850473724927, 
    -0.00044746002782841481, -0.00012087458858099706, 0.00022366106096602807, 
    0.00058306688961684496, 0.00095413000084668858, 0.0013335935472551857, 
    0.0017182442250229764, 0.0021049768780304614, 0.0024908389245485245, 
    0.0028730457471275892, 0.0032489765271682884, 0.0036161554665817873, 
    0.0039722270133569727, 0.0043149291733011862, 0.0046420909157512897, 
    0.004951642375597109, 0.005241630709725378, 0.0055102640014744247, 
    0.0057559499073023407, 0.0059773352700649793, 0.0061733471860454222, 
    0.0063432118952955231, 0.0064864666029329568, 0.0066029471014781788, 
    0.0066927590862050383, 0.0067562254406758511, 0.0067938182150652053, 
    0.0068060929522295753, 0.0067936264055456583, 0.0067569742848475698, 
    0.006696648304292261, 0.0066131230969675827, 0.0065068610914840496, 
    0.006378349598741645, 0.0062281588152154855, 0.0060569993083794344, 
    0.00586577935462916, 0.0056556566246595049, 0.0054280725507257306, 
    0.0051847751750110412, 0.0049278130277774579, 0.0046594987084537468, 
    0.004382334329716602, 0.0040989081711885781, 0.0038117733538745508, 
    0.0035233204110565143, 0.0032356677000092383, 0.0029505675070158983, 
    0.0026693485532940748, 0.0023928919468336365, 0.0021216335697227529, 
    0.0018556033771072286, 0.001594491253773879, 0.0013377363031627635, 
    0.0010846391741192746, 0.00083448292125083354, 0.00058666463576264563, 
    0.00034080597410185496, 9.6861447622707841e-05, -0.00014480530085980508, 
    -0.00038336321240651399, -0.00061747854883587288, 
    -0.00084530342195215978, -0.001064497485252451, -0.0012722727628560995, 
    -0.0014654768346842055, -0.0016407005418773847, -0.0017944126789511314, 
    -0.0019231130952496905, -0.0020234852496188718, -0.0020925397250063024, 
    -0.0021277367511634902, -0.0021270946882953595, -0.0020892684475234866, 
    -0.0020136081461319113, -0.0019001902230148496, -0.001749816754583072, 
    -0.0015639938959407045, -0.0013448653369570241, -0.0010951289753289128, 
    -0.00081792863374353475, -0.00051672643823142956, 
    -0.00019519202703540482, 0.00014291119603286408, 0.00049380687470395668, 
    0.00085374695054527233, 0.0012190400820532323, 0.0015860247623582851, 
    0.0019510415715847671, 0.0023103929190325676, 0.0026603217868523482, 
    0.0029970110712757175, 0.0033166162711496267, 0.003615331239062556, 
    0.0038894970093946027, 0.0041357307428161886, 0.0043510806340477451, 
    0.0045331618265083574, 0.0046802784865677561, 0.0047915189569015266, 
    0.0048667987956131026, 0.0049068620790556575, 0.0049132428532027306, 
    0.0048881808797391971, 0.0048345057219149491, 0.0047554924334103337, 
    0.0046547053817024165, 0.0045358482628077091, 0.0044026274225169018, 
    0.0042586477560694622, 0.0041073423098126434, 0.0039519278818894053, 
    0.0037953832087910229, 0.0036404412429683706, 0.0034895850630191003, 
    0.0033450463260621291, 0.0032088009004482428, 0.0030825640594357834, 
    0.0029677860836942035, 0.0028656516031530946, 0.0027770586229560468, 
    0.0027025985605444872, 0.002642532609744798, 0.0025967761950181564, 
    0.0025648975680807973, 0.0025461487357430358, 0.002539508900924066, 
    0.0025437451149704863, 0.0025574574928566903, 0.002579123858882237, 
    0.0026071201333266094, 0.00263972942041759, 0.0026751698531529353, 
    0.0027116245987044907, 0.0027472939849533503, 0.0027804581377712106, 
    0.0028095549762082589, 0.0028332339971383798, 0.0028504315585955375, 
    0.0028604178268806595, 0.0028628246207250906, 0.0028576518497584989, 
    0.0028452507563149002, 0.002826290353101773, 0.0028017097456867202, 
    0.0027726584211301406, 0.0027404351155151593, 0.0027064336689548809, 
    0.0026720949513727222, 0.0026388571563085144, 0.0026081166756452934, 
    0.0025812003821846967, 0.0025593343809077037, 0.0025436280560331903, 
    0.0025350557803883022, 0.0025344381045377816, 0.0025424236031293735, 
    0.002559469408671819, 0.0025858272188476568, 0.0026215269040983889, 
    0.0026663824045210925, 0.0027200005271456398, 0.0027817935036847344, 
    0.0028510000499737701, 0.0029266767749852327, 0.0030076993565902647, 
    0.0030927363813023157, 0.0031802431129155273, 0.0032684500930544903, 
    0.0033553709131556898, 0.0034388271673194627, 0.0035165076895905902, 
    0.0035860326728018766, 0.0036450426171608604, 0.0036912949394967386, 
    0.0037227715644940853, 0.0037377772222954822, 0.0037350403865345928, 
    0.0037138060893190839, 0.0036739086512463845, 0.003615829996739981, 
    0.0035407263626927917, 0.0034504329043688461, 0.0033474372893390041, 
    0.0032348167415491339, 0.0031161395228959136, 0.0029953322284801999, 
    0.0028765117088513561, 0.0027637939227524201, 0.0026610859878744854, 
    0.0025718853252231851, 0.0024990779319029551, 0.0024447900877862163, 
    0.0024102800791470716, 0.0023958953667294323, 0.0024010930967150027, 
    0.002424510695053591, 0.0024640705031096933, 0.0025171031002870431, 
    0.002580476076829809, 0.0026507377831306938, 0.0027242518857163935, 
    0.0027973243029356392, 0.002866340650228076, 0.0029278821893913964, 
    0.0029788304503356468, 0.0030164629992898164, 0.003038513990706611, 
    0.0030432061121694366, 0.003029251614547986, 0.0029958028099356599, 
    0.0029423871658074367, 0.0028688090954072801, 0.0027750518228945669, 
    0.0026611869171945285, 0.0025273060882538014, 0.0023734896901757992, 
    0.0021997998946332014, 0.0020063087786542947, 0.0017931545177020999, 
    0.0015606150085630348, 0.0013091949626595888, 0.0010397113507323954, 
    0.00075336764124335823, 0.00045182029529173477, 0.0001372069804092046, 
    -0.00018784948973335516, -0.00052026248426787077, 
    -0.00085653667228748976, -0.0011928413486602943, -0.001525113396361548, 
    -0.0018491640055306995, -0.0021608006022343948, -0.0024559460197944591, 
    -0.0027307562732418644, -0.0029817121742988749, -0.0032057029426840215, 
    -0.003400079892836558, -0.0035627065222977247, -0.0036919709999732797, 
    -0.0037868102905233977, -0.003846703867816533, -0.0038716695360420461, 
    -0.0038622453195130122, -0.0038194623234130412, -0.0037448113014458342, 
    -0.003640191190901503, -0.0035078513565161935, -0.0033503330248641412, 
    -0.0031704086202096211, -0.002971019395201628, -0.0027552267188765594, 
    -0.002526151593095694, -0.002286931194889606, -0.0020406698423722116, 
    -0.0017903866642346737, -0.0015389779408114094, -0.0012891896017449653, 
    -0.0010436009086530387, -0.0008046201956323374, -0.00057448509783670403, 
    -0.00035524889601085629, -0.00014876218472820453, 4.3376436806349974e-05, 
    0.00021988160144138682, 0.00037984759050663664, 0.00052280254895706443, 
    0.00064873336918785962, 0.00075808276666578997, 0.00085170174170616736, 
    0.00093078766202822258, 0.00099676893990616254, 0.0010512075242513756, 
    0.0010956902278432372, 0.0011317559462059273, 0.0011608352122656584, 
    0.0011842359320506641, 0.0012031698518837845, 0.0012187912723173916, 
    0.0012322565611820682, 0.0012447851411357587, 0.0012577094240396442, 
    0.0012724994704342274, 0.0012907640085247116, 0.0013142105933739107, 
    0.0013445853165975283, 0.0013835779730844448, 0.0014327194967555495, 
    0.0014932787382963826, 0.0015661670279204761, 0.0016518603400365972, 
    0.0017503446413923937, 0.001861081861274057, 0.0019830040800592852, 
    0.0021145381314861926, 0.0022536518773446671, 0.0023979284685222038, 
    0.0025446546015700814, 0.0026909286544284077, 0.002833777010369444, 
    0.0029702639315450051, 0.0030976151999863076, 0.0032133100198444868, 
    0.0033151654847481137, 0.003401391321434832, 0.0034706323938632926, 
    0.0035219841087292666, 0.0035550045813256478, 0.0035696943109124035, 
    0.0035664779323014819, 0.0035461645858920862, 0.0035098872601323924, 
    0.0034590295452525763, 0.0033951401422263471, 0.0033198500846120891, 
    0.0032347772872754498, 0.0031414447485131509, 0.0030412012725102274, 
    0.0029351443367536005, 0.0028240661369862588, 0.0027083955671095301, 
    0.0025882071396599957, 0.0024632474709181712, 0.0023330467686533247, 
    0.0021970425125862315, 0.0020547423346347375, 0.0019058797730638472, 
    0.0017505403559482445, 0.0015892413216996759, 0.0014229719919917234, 
    0.0012531900512922078, 0.0010817963432875103, 0.00091108415637993173, 
    0.0007436693374328156, 0.0005824134863659609, 0.00043031151668285693, 
    0.00029038682123998022, 0.00016557773589356432, 5.8623041053009731e-05, 
    -2.8053071732167241e-05, -9.2437313247521464e-05, 
    -0.00013301590632579902, -0.000148845823060489, -0.00013962124657094485, 
    -0.00010572245920983708, -4.8258947345988193e-05, 3.0929435331755089e-05, 
    0.00012929207068719319, 0.00024364210734654612, 0.00037026873325057591, 
    0.00050508445926084836, 0.00064381891626105422, 0.00078220162823227691, 
    0.00091614477558351031, 0.0010419108556733404, 0.0011562311190145952, 
    0.0012564026176859967, 0.0013403311330133171, 0.0014065334280832611, 
    0.0014541096373143988, 0.001482679535655822, 0.0014923123034619669, 
    0.0014834419510666003, 0.0014568105222979011, 0.0014134101903264217, 
    0.0013544389521007608, 0.0012812711237642498, 0.0011954243062112422, 
    0.0010985332566739617, 0.00099233131460567023, 0.00087864567060306456, 
    0.00075940315552557014, 0.00063663971551149862, 0.00051252204742467254, 
    0.00038935727634040434, 0.00026958458713982852, 0.00015577305476877719, 
    5.0588759063739555e-05, -4.3244425848316254e-05, -0.00012300273171855986, 
    -0.00018603547434669135, -0.00022983997981128248, 
    -0.00025215604539827478, -0.00025105419216197168, 
    -0.00022501360690920056, -0.00017298743190261501, -9.444813280655006e-05, 
    1.0583595007538889e-05, 0.00014154236894969928, 0.00029735000006901889, 
    0.0004764732794226333, 0.00067699891208438203, 0.00089672875401382605, 
    0.0011332639474640163, 0.001384105535694331, 0.0016467072690597771, 
    0.0019185372019427036, 0.0021971089119374003, 0.002480009958900015, 
    0.0027649368265315476, 0.0030497352283532582, 0.0033324478556054286, 
    0.0036113669387496136, 0.0038850687388165043, 0.0041524368722304248, 
    0.0044126580453529964, 0.0046652024232348753, 0.0049097671131449203, 
    0.0051462075775571521, 0.0053744589765362854, 0.0055944424654676052, 
    0.0058059921308692523, 0.0060087758017157225, 0.0062022610206999155, 
    0.0063856855933306445, 0.0065580534333700763, 0.0067181540123700725, 
    0.0068645904906313353, 0.006995815527385923, 0.0071101753970506673, 
    0.0072059689021740352, 0.0072815180960833139, 0.0073352470193353341, 
    0.0073657764107136914, 0.0073720086651511176, 0.0073531943307282811, 
    0.0073089835049697698, 0.0072394452337854204, 0.0071450539600785533, 
    0.0070266641822143315, 0.0068854780320852012, 0.0067230069395146589, 
    0.006541033170492417, 0.0063415798411443425, 0.0061268786874625484, 
    0.0058993187015429563, 0.005661403231305622, 0.005415692046752749, 
    0.0051647488204494265, 0.0049110945006729982, 0.0046571769155609186, 
    0.0044053480652267935, 0.0041578634891461814, 0.0039168682282895353, 
    0.0036843857806119137, 0.0034622875644574414, 0.0032522580139775475, 
    0.0030557580273641717, 0.0028739735798852997, 0.0027077809720597273, 
    0.002557716694892841, 0.0024239540816444801, 0.0023063134364364273, 
    0.0022042688801500445, 0.002116976652169662, 0.0020433224384297502, 
    0.0019819715129431917, 0.0019314269842036274, 0.0018901035183564148, 
    0.0018563919273844156, 0.0018287387443080099, 0.0018057086969529002, 
    0.0017860547065472689, 0.0017687562568663069, 0.0017530713192164457, 
    0.0017385512195824307, 0.0017250551574109979, 0.0017127550717916467, 
    0.0017021180595913077, 0.0016938647999620723, 0.0016889281442764937, 
    0.0016883801604615398, 0.0016933648061130875, 0.0017050057279775622, 
    0.0017243451171891316, 0.0017522394399968211, 0.0017892998502675021, 
    0.0018358367084538661, 0.0018918044588551804, 0.001956783837877952, 
    0.0020299526056894932, 0.0021100798358082763, 0.0021955219741939787, 
    0.0022842401797041204, 0.002373854096187037, 0.002461721863063079, 
    0.0025450343461861985, 0.0026209636053088591, 0.002686804141426362, 
    0.0027401345398094584, 0.0027789441367843679, 0.002801750779841604, 
    0.0028076641878143141, 0.0027963846511152206, 0.0027681841508787053, 
    0.0027238231843089542, 0.002664473360155642, 0.0025916333989097571, 
    0.0025070573516636418, 0.0024127247188923395, 0.0023108171413796369, 
    0.0022037045263246517, 0.0020939123808572432, 0.0019840758363101549, 
    0.001876860597187689, 0.0017748545045252594, 0.0016804493421126282, 
    0.0015957206763198104, 0.0015223097826539693, 0.0014613403186150499, 
    0.0014133630236635509, 0.0013783457422100018, 0.0013556912878840909, 
    0.0013443095761901773, 0.0013427208084325569, 0.0013491635892289786, 
    0.0013617373774670459, 0.0013785271185658423, 0.0013977134249758506, 
    0.0014176675818117039, 0.0014370373479615881, 0.0014548181559616985, 
    0.001470412807366706, 0.0014836651898758782, 0.0014948976141081077, 
    0.0015049002532029326, 0.0015148952672138802, 0.0015264391557016077, 
    0.0015412801084402014, 0.0015612059989758063, 0.0015878636568949945, 
    0.00162261156893676, 0.0016663896847560738, 0.0017196312361059118, 
    0.0017822030669495301, 0.0018533731047806821, 0.0019317913031297795, 
    0.002015467974152238, 0.0021017835661192082, 0.0021875320117779704, 
    0.0022690515625204519, 0.0023423975982166884, 0.0024035650410399018, 
    0.0024487355897814442, 0.0024744858182002274, 0.002477964323443816, 
    0.0024570298979800721, 0.002410350732938459, 0.0023374907659688233, 
    0.0022389482357967061, 0.0021161603043753975, 0.0019714750996477938, 
    0.0018080560271159717, 0.0016297447971775447, 0.0014409127689718737, 
    0.0012462635767726655, 0.0010506337802844983, 0.00085880542796804211, 
    0.00067532242281016818, 0.00050435122511356505, 0.00034956760639036951, 
    0.00021409046975328434, 0.00010045550689437717, 1.0617365551405671e-05, 
    -5.4010934560855657e-05, -9.2517435214107261e-05, 
    -0.00010445150062788231, -8.9772654278405089e-05, 
    -4.8798003874182024e-05, 1.78462921747099e-05, 0.00010929047868393744, 
    0.00022448593313934522, 0.00036224356701633552, 0.00052127848853983014, 
    0.00070024016608044581, 0.00089773297466534294, 0.0011123420077263307, 
    0.0013426626875799319, 0.0015873348010190676, 0.0018450737136310453, 
    0.002114691198850853, 0.0023951026256845173, 0.0026853042317821004, 
    0.0029843403971170773, 0.0032912581704011849, 0.0036050455881711419, 
    0.003924553409996874, 0.0042484453239556678, 0.0045751260681326815, 
    0.0049026990778206587, 0.0052289260729305436, 0.0055512097827157851, 
    0.0058666124334660766, 0.0061719147247228873, 0.0064636982705840243, 
    0.0067384771604104112, 0.0069928321947158242, 0.0072235878369092156, 
    0.007427965040382979, 0.0076037359961166453, 0.0077493271902541695, 
    0.0078638994777761977, 0.0079473863040992673, 0.0080004767102348114, 
    0.008024566341091624, 0.0080216863186862806, 0.0079944086503205627, 
    0.0079457198663561192, 0.0078788716094556656, 0.0077972086510753923, 
    0.0077039964204141656, 0.007602246477347252, 0.007494559315937053, 
    0.0073830036856124097, 0.0072690338453117341, 0.007153441085779126, 
    0.0070363485246956103, 0.0069172404836720458, 0.0067950235016405666, 
    0.0066681255363048716, 0.0065346860319860619, 0.0063927789899982292, 
    0.0062406489914777078, 0.0060769604654300488, 0.0059009798511435538, 
    0.0057127265491967163, 0.0055130495323830412, 0.005303652225717455, 
    0.0050870674727834155, 0.0048666040643350027, 0.00464623173904053, 
    0.0044304351075816744, 0.0042240188623367285, 0.0040318902953096576, 
    0.003858809761530131, 0.0037091510648307748, 0.003586669088969846, 
    0.0034942962197911324, 0.0034339801808001896, 0.0034065632994454255, 
    0.0034116700010183945, 0.0034477098500540629, 0.0035118896925861827, 
    0.0036003571228213366, 0.0037083908356266393, 0.003830638264285726, 
    0.0039613504477660306, 0.0040945942732061617, 0.0042244058954374678, 
    0.0043449189194500653, 0.0044504898161778069, 0.0045358332389614951, 
    0.0045962382559181156, 0.0046277884210393794, 0.0046275554423489684, 
    0.0045937200179927955, 0.0045256137602972986, 0.0044236652668826499, 
    0.004289258820169675, 0.0041245718262517212, 0.003932355429525366, 
    0.0037157445960090806, 0.0034780639452539051, 0.0032226698684603579, 
    0.0029528417044171911, 0.0026716976132254043, 0.0023821594011196674, 
    0.0020869413556051427, 0.0017885574759996994, 0.0014893440141859396, 
    0.0011914746343824625, 0.00089698695727551386, 0.00060781781233250755, 
    0.0003258435341143712, 5.2900675470942754e-05, -0.00020919214008242499, 
    -0.00045864903167317671, -0.00069374927010623481, 
    -0.00091285731296710719, -0.0011144444149429216, -0.0012970751829461491, 
    -0.0014593736768988108, -0.0015999963469282867, -0.0017176469704296691, 
    -0.0018111108326285842, -0.0018793682638308222, -0.0019217155771575304, 
    -0.0019378856026779803, -0.0019281143027092154, -0.0018931873749638895, 
    -0.0018344397576568249, -0.0017536739776883501, -0.0016530957684231114, 
    -0.0015351959201651663, -0.001402692490567135, -0.001258450504992196, 
    -0.0011054397003453478, -0.00094670622134541027, -0.00078531848858137861, 
    -0.00062433510539732927, -0.00046675787653669809, 
    -0.00031546607079717799, -0.00017314739692556367, 
    -4.2219399255742694e-05, 7.5246254549653495e-05, 0.00017757994771800355, 
    0.00026355054603417787, 0.0003323903291532356, 0.0003837905598758325, 
    0.00041785925320232068, 0.00043507485016651209, 0.00043621173243537151, 
    0.00042226139244648151, 0.00039434279638245987, 0.00035363326630549741, 
    0.00030127744264994054, 0.0002382880004459578, 0.00016546002189122555, 
    8.3273525900006838e-05, -8.1825329146416391e-06, -0.00010923001824497431, 
    -0.00022055561708011394, -0.00034312127459908397, 
    -0.00047806193371075146, -0.0006265235607344139, -0.00078954165607591912, 
    -0.00096792872111402543, -0.0011622124351174296, -0.0013726011897526309, 
    -0.0015989818100610974, -0.001840939813424649, -0.0020977761331807754, 
    -0.0023685091514292229, -0.0026518427967453817, -0.0029461571575887888, 
    -0.0032494971637875049, -0.0035595599719227423, -0.0038737364665109237, 
    -0.0041891399195051471, -0.0045026602781548008, -0.0048110653285823816, 
    -0.0051110940012397636, -0.0053995199707939714, -0.0056732543576224715, 
    -0.0059293846614934765, -0.0061651799220781159, -0.0063780763875336171, 
    -0.0065656496366404658, -0.0067255657414221296, -0.0068555313529270988, 
    -0.0069532752139289285, -0.0070165355709613259, -0.0070431060767179102, 
    -0.0070308886660750223, -0.0069779928133666888, -0.0068828511714269253, 
    -0.0067443174252137823, -0.0065618136551076735, -0.0063353983738339567, 
    -0.006065841835115774, -0.0057545893840888884, -0.0054036956257699081, 
    -0.0050157091720297959, -0.0045935315020811272, -0.004140276919098876, 
    -0.0036591774501806389, -0.0031534780432782451, -0.0026263822943084557, 
    -0.0020809943113970419, -0.0015202855273892784, -0.00094708449430521043, 
    -0.00036407353481555113, 0.00022615517530570118, 0.00082106747730307248, 
    0.0014181151503046363, 0.0020146640574129839, 0.0026079402572326683, 
    0.0031950103498073713, 0.0037727987024982436, 0.0043381593891015065, 
    0.0048879390086566483, 0.0054191007936901688, 0.0059288148929373518, 
    0.0064145541018833024, 0.0068741371816879024, 0.0073057434488270276, 
    0.0077078685576111305, 0.0080792757947742242, 0.0084189319814081051, 
    0.0087259683025294778, 0.008999660172592204, 0.0092394205569628976, 
    0.0094448559382563999, 0.0096157824469627652, 0.0097522861168303516, 
    0.0098547653399533117, 0.0099239561209793787, 0.009960938720087166, 
    0.0099671386948382758, 0.0099443262481627506, 0.0098945534118569916, 
    0.0098201173633381735, 0.0097234744454903176, 0.0096071205462579263, 
    0.0094734761037413191, 0.0093247702761443986, 0.0091629116703759294, 
    0.0089894059671884637, 0.0088053049372043782, 0.0086111865730775349, 
    0.0084071740233216449, 0.0081929778152352046, 0.0079679652819159355, 
    0.0077312523068602413, 0.0074817925840038289, 0.0072184612061365408, 
    0.0069400997762382073, 0.006645520893516897, 0.0063335365768681113, 
    0.0060029421746480164, 0.0056525429960335178, 0.0052811864080464068, 
    0.0048877786137313988, 0.0044713899503613739, 0.0040313206728879464, 
    0.0035671747019549362, 0.003078946201261324, 0.0025670804068946987, 
    0.0020325293934469134, 0.0014767657764675657, 0.00090177511507327692, 
    0.00031001201348110395, -0.00029565431743747215, -0.00091197396159060007, 
    -0.0015353735798851874, -0.002162015758219402, -0.0027878410461557846, 
    -0.0034086573521936213, -0.0040202267718720975, -0.0046184147048521597, 
    -0.0051993500986816914, -0.0057596052022483918, -0.0062963621096583915, 
    -0.0068075448089743133, -0.007291920784682107, -0.0077491302613855676, 
    -0.0081796992219613038, -0.0085850139230827602, -0.0089672397603819433, 
    -0.0093292285463587553, -0.0096743587787622674, -0.010006352289632241, 
    -0.010329088011458104, -0.010646396804528294, -0.010961911345396511, 
    -0.01127900658545292, -0.011600750605445498, -0.011929971021720564, 
    -0.012269314639539359, -0.012621338078507027, -0.012988518932696197, 
    -0.013373233487197338, -0.013777650312720317, -0.014203624982891886, 
    -0.014652530375735754, -0.015125058386146882, -0.015621079860696939, 
    -0.016139487889632768, -0.016678092989301167, -0.017233605357172669, 
    -0.017801665442496305, -0.018376973576054823, -0.018953453976878455, 
    -0.019524509742974153, -0.020083283840765593, -0.020622970794344508, 
    -0.021137139364888403, -0.021620010561696341, -0.02206672374611799, 
    -0.022473540979718942, -0.022837973829427739, -0.023158846819917249, 
    -0.023436276976775628, -0.023671547370630024, -0.023866987432083164, 
    -0.02402576518170749, -0.024151682165669135, -0.024249026018750633, 
    -0.024322344818084218, -0.024376325916325704, -0.024415606482008592, 
    -0.024444592530227134, -0.024467300752297652, -0.024487177464581372, 
    -0.024507019752345639, -0.024528932153289947, -0.024554366834161435, 
    -0.024584232196630487, -0.024619001321132639, -0.024658782542427215, 
    -0.024703253198403875, -0.02475160784362956, -0.024802347001266115, 
    -0.02485314959423128, -0.024900734468153534, -0.024940791405931882, 
    -0.02496793167687791, -0.02497574188199269, -0.02495691890449412, 
    -0.024903505256577783, -0.024807202334469376, -0.024659712253126038, 
    -0.024453094149834667, -0.024180166291513396, -0.023834761487701941, 
    -0.023412042699395976, -0.022908740549125822, -0.022323371609692461, 
    -0.021656454997482713, -0.02091067055367668, -0.020090917014428701, 
    -0.019204299511267425, -0.01826001177954012, -0.017269147527288104, 
    -0.01624442299066357, -0.015199860608865958, -0.014150406896710965, 
    -0.013111578129793031, -0.012099081656986406, -0.011128381107548149, 
    -0.010214343162761043, -0.0093707484514890804, -0.0086099169137204973, 
    -0.0079422906963504212, -0.0073760424523650276, -0.0069167845041079746, 
    -0.0065673719155255657, -0.0063278325847755095, -0.0061955010470532762, 
    -0.0061651926383401567, -0.0062296022405173039, -0.006379746331348044, 
    -0.0066054250555666839, -0.0068957543404068473, -0.0072396235568571426, 
    -0.0076260788914406328, -0.0080445710669822812, -0.0084850241580308652, 
    -0.0089377869849114628, -0.0093934626663648314, -0.0098427791996464117, 
    -0.010276655128097513, -0.010686399653681688, -0.011064025476808455, 
    -0.011402612825070154, -0.01169658569750506, -0.011941978765573832, 
    -0.012136530228537215, -0.012279769696326846, -0.012372968037484035, 
    -0.012419047049421778, -0.012422408495113042, -0.012388751034753608, 
    -0.012324845732574845, -0.012238309849429332, -0.012137352295518227, 
    -0.012030535023282475, -0.011926574146882082, -0.011834122958005389, 
    -0.011761527034531242, -0.01171658593020047, -0.011706365332239088, 
    -0.011736935740599537, -0.011813248336846072, -0.01193903068275428, 
    -0.012116727695572715, -0.012347506908778496, -0.012631223797782353, 
    -0.012966386840806698, -0.013350022162268898, -0.013777614046840905, 
    -0.014243086657966437, -0.014738950041405331, -0.015256700192914583, 
    -0.015787322936673242, -0.016322029469690465, -0.016852976340229111, 
    -0.017373959263897523, -0.017881031199985402, -0.018372912971038158, 
    -0.018851084310705264, -0.019319670658316364, -0.019784979882519895, 
    -0.020254742504540589, -0.020737269458307322, -0.021240560907926663, 
    -0.021771557074419755, -0.022335526227752391, -0.022935843973421605, 
    -0.023574053444889852, -0.024250146264580826, -0.024962986952643526, 
    -0.025710718198500716, -0.026491235770646639, -0.027302301772076661, 
    -0.028141749364136683, -0.029007333762473404, -0.0298965941296854, 
    -0.030806473999087328, -0.031732935417339132, -0.03267057656313993, 
    -0.033612310704672417, -0.034549309760696423, -0.035470944914427635, 
    -0.036365116559304918, -0.037218584599157681, -0.038017447309277572, 
    -0.038747637307104281, -0.039395565572362561, -0.039948747779180047, 
    -0.040396634784236607, -0.040731235477133185, -0.040947873037564801, 
    -0.041045512086777862, -0.041026979114168513, -0.04089859965887304, 
    -0.040669620856378194, -0.040351217855009287, -0.039955907699081132, 
    -0.039496658163272823, -0.038986482943774499, -0.038437930435558001, 
    -0.037863118641817399, -0.037273854736691703, -0.036681926518108678, 
    -0.036099456914739897, -0.035539190092670377, -0.035014587773638639, 
    -0.034539495918925446, -0.034127922461276654, -0.033793398151334475, 
    -0.033548556286081568, -0.033404700433248655, -0.033371466097782444, 
    -0.033456103195043878, -0.033663156492815788, -0.033993841454254506, 
    -0.034445654126239941, -0.03501260097651842, -0.035685618106505716, 
    -0.036453369630920898, -0.037302276907407485, -0.038216951023044773, 
    -0.039180369971948556, -0.040173541521585809, -0.041175589241897959, 
    -0.042163916343148547, -0.043114835282750986, -0.044004599514642355, 
    -0.044811044206886197, -0.04551647017275242, -0.04610920728324093, 
    -0.046585224026482477, -0.04694951483712647, -0.047215370699370061, 
    -0.047402093239950878,
  // Fqt-F(5, 0-1999)
    1, 0.99603270247494524, 0.98425448944376104, 0.96502982135976823, 
    0.93894127502175539, 0.90675371487132428, 0.86936942167115616, 
    0.8277784589729027, 0.78300858589192235, 0.73607854907868475, 
    0.68795770751977536, 0.63953391868648102, 0.59159056551464417, 
    0.54479264054641896, 0.49968114138112124, 0.45667449777142149, 
    0.41607549120684945, 0.37808212644648814, 0.34280092382298394, 
    0.31026131906865617, 0.28043014526293747, 0.25322537608088785, 
    0.22852859736221895, 0.20619590978991578, 0.186067135859148, 
    0.16797340280960135, 0.15174318647256785, 0.13720702575123775, 
    0.12420106160101109, 0.11256958402697927, 0.10216677662200602, 
    0.092857765879710147, 0.084519158142604411, 0.077039129893241742, 
    0.070317227874026375, 0.064263938178633295, 0.058800111022257982, 
    0.053856290258615179, 0.049371986363974052, 0.045294932755715958, 
    0.04158032995884569, 0.038190102306960148, 0.035092137711836044, 
    0.032259555181368089, 0.029669947869924791, 0.027304661940199332, 
    0.0251481120874378, 0.023187134876719181, 0.021410418922418406, 
    0.019807999688447431, 0.018370843288563841, 0.017090506660577345, 
    0.015958866039470287, 0.014967931029058084, 0.014109692100127564, 
    0.013376021946548409, 0.012758599114011775, 0.012248844011646977, 
    0.011837869193416008, 0.011516435532144955, 0.011274921689368255, 
    0.011103326747767154, 0.010991309730799152, 0.010928275404622424, 
    0.010903503339259201, 0.0109063095588398, 0.010926230432115413, 
    0.010953194633941522, 0.010977693557803954, 0.01099091957228567, 
    0.010984894745263544, 0.01095255522838017, 0.010887832301354825, 
    0.010785683590419983, 0.010642124360743807, 0.010454226968960641, 
    0.010220124873514829, 0.0099390139932634854, 0.0096111480277774625, 
    0.0092378325387935702, 0.0088213968141886666, 0.0083651345643799609, 
    0.0078732315032588995, 0.0073506365597981738, 0.0068029159831732742, 
    0.0062360703207497148, 0.0056563369150723422, 0.005069971342545939, 
    0.0044830329506949391, 0.003901167496565475, 0.0033294043756894121, 
    0.0027719691348852965, 0.0022321311358334947, 0.0017121043574182917, 
    0.0012130130371618636, 0.00073493385496750468, 0.00027701516075007615, 
    -0.0001623255219525161, -0.00058515341563763817, -0.00099372719379572558, 
    -0.0013902068524236752, -0.0017763674975958799, -0.0021533614585050737, 
    -0.0025215527097058239, -0.0028804246281000511, -0.003228590228962189, 
    -0.0035638942836967876, -0.0038835844308335293, -0.0041845548265274542, 
    -0.0044636194640232376, -0.0047177915521437143, -0.0049445451690176088, 
    -0.0051420328704544563, -0.0053092491851253433, -0.0054461211980128066, 
    -0.0055535290776042084, -0.0056332497549007581, -0.0056878417845186054, 
    -0.0057204798080473414, -0.0057347621085885331, -0.0057345090385250083, 
    -0.005723558987883166, -0.0057055877509544243, -0.0056839393380918399, 
    -0.0056614881946899856, -0.0056405252260450876, -0.0056226700229590016, 
    -0.0056088126031292977, -0.0055990800610743047, -0.0055928344417541581, 
    -0.0055887077335092499, -0.005584667115802135, -0.0055781014831644739, 
    -0.0055659380579182807, -0.0055447593400147228, -0.0055109267817085566, 
    -0.0054606964670485076, -0.0053903324872653135, -0.0052962204178164133, 
    -0.0051749849873111119, -0.0050236086217948219, -0.0048395480836638501, 
    -0.0046208561906953523, -0.0043662857785353292, -0.004075381060157833, 
    -0.0037485492723474114, -0.0033871191611555759, -0.0029933588642004592, 
    -0.0025704721057479341, -0.0021225604370986501, -0.0016545420285383463, 
    -0.0011720258998296029, -0.00068115526685429465, -0.00018841664848659261, 
    0.00029958547814824138, 0.00077636760731256008, 0.0012358185771455183, 
    0.00167244252609043, 0.002081594088341009, 0.0024596651856807869, 
    0.0028042278068999621, 0.0031141080731302427, 0.0033893793797737724, 
    0.0036312726382280937, 0.0038420068307857677, 0.0040245631781111154, 
    0.0041824286532738788, 0.0043193118307581716, 0.0044388717301946596, 
    0.0045444665495611497, 0.0046389393290849944, 0.0047244652472150771, 
    0.0048024608939430868, 0.0048735595970011633, 0.0049376533798809619, 
    0.0049939817457843698, 0.0050412528356081994, 0.0050777811134038505, 
    0.0051016356803787605, 0.0051107709821358645, 0.0051031542907500338, 
    0.0050768728575733913, 0.0050302283373985235, 0.0049618063067667232, 
    0.0048705457071361487, 0.0047557714547762598, 0.0046172204941521645, 
    0.0044550357257546825, 0.0042697485777625256, 0.0040622460572457319, 
    0.003833728568577562, 0.0035856643933739061, 0.0033197440449799979, 
    0.0030378435014179915, 0.0027419914022600396, 0.0024343386961951452, 
    0.0021171371556681388, 0.0017927295562994512, 0.0014635489578161899, 
    0.0011321193496198958, 0.00080106493016026195, 0.00047310313654103499, 
    0.00015103205084028082, -0.00016230413093859446, -0.00046404828540712393, 
    -0.00075137701906377878, -0.0010215489153759651, -0.0012719481490496118, 
    -0.0015001357046395595, -0.0017039017358550469, -0.0018813294824378873, 
    -0.0020308677870431112, -0.002151402357834219, -0.0022423348003074491, 
    -0.0023036490310634227, -0.002335960669905835, -0.0023405429929993517, 
    -0.00231932106396688, -0.0022748346493922521, -0.0022101677865236755, 
    -0.0021288395132166905, -0.0020346703732765084, -0.0019316297007413851, 
    -0.001823673698719175, -0.0017145950555061279, -0.0016078914126090595, 
    -0.0015066569840238809, -0.0014135080479475844, -0.0013305428036716111, 
    -0.001259329346561253, -0.0012009283540280549, -0.0011559251824090446, 
    -0.0011244798768196215, -0.0011063775429870828, -0.0011010825924573748, 
    -0.0011077991995061317, -0.0011255351783648914, -0.001153167719629524, 
    -0.001189512927681853, -0.0012333924805849293, -0.0012836848685298316, 
    -0.0013393695052573537, -0.001399555192928688, -0.001463484348934862, 
    -0.0015305525198726576, -0.0016003031500934932, -0.0016724357402081789, 
    -0.0017468070768532054, -0.0018234323379594801, -0.0019024709466470828, 
    -0.001984209432451505, -0.0020690303640214553, -0.0021573738827268454, 
    -0.0022496869090085497, -0.0023463731448061039, -0.0024477302674663598, 
    -0.002553898652900588, -0.0026648074669785326, -0.0027801405361561398, 
    -0.0028993154348504468, -0.0030214846253187335, -0.0031455612089274889, 
    -0.0032702629777553302, -0.0033941722508237342, -0.0035158136838345901, 
    -0.0036337294866641647, -0.0037465664866722474, -0.0038531515590031059, 
    -0.0039525611175640508, -0.0040441771274799011, -0.0041277210602777923, 
    -0.0042032617671986586, -0.0042711946566157928, -0.0043321817671141058, 
    -0.0043870593976308627, -0.0044367202087289472, -0.0044819770055752354, 
    -0.0045234225061574563, -0.0045613079381427064, -0.0045954439557000046, 
    -0.0046251402627147126, -0.0046491912111798362, -0.0046659152690240579, 
    -0.004673241616743669, -0.0046688300462252924, -0.0046502316820436831, 
    -0.0046150615495125624, -0.0045611837487733436, -0.0044868875153284945, 
    -0.0043910513815237379, -0.0042732772117760574, -0.0041339807191120813, 
    -0.0039744335532869548, -0.0037967518195286191, -0.0036038217842218724, 
    -0.003399169162865845, -0.0031867796250810904, -0.0029708790468764303, 
    -0.0027556941593644751, -0.002545202560469445, -0.0023429062388617026, 
    -0.0021516315944193846, -0.0019733787354382177, -0.0018092235610943958, 
    -0.0016592712519067285, -0.0015226664765023016, -0.001397640738112337, 
    -0.0012815936610778924, -0.0011711970680981214, -0.0010625337468015265, 
    -0.00095127165564960921, -0.00083287126477731769, 
    -0.00070283047927910782, -0.00055692630689111193, 
    -0.00039144662209885913, -0.00020337904815891442, 9.4679251659193341e-06, 
    0.00024838195693492539, 0.00051372114925101083, 0.00080492283511470494, 
    0.0011205323783521008, 0.0014582583852716141, 0.0018150367192979744, 
    0.0021871085845753995, 0.0025701211930839693, 0.0029592398439192728, 
    0.0033492831780936923, 0.0037348839466556541, 0.0041106661583585353, 
    0.0044714319481448765, 0.0048123735278790478, 0.0051292602427974307, 
    0.0054186202662190059, 0.0056778751634734368, 0.0059054288110822655, 
    0.0061006954617415475, 0.0062640622004196903, 0.0063967952340770236, 
    0.0065008990355861314, 0.0065789470904599225, 0.006633895998473441, 
    0.0066688956188364181, 0.0066871042677495848, 0.0066915343357054347, 
    0.0066848942212968301, 0.0066694658238813116, 0.0066470157977491159, 
    0.0066187344737023259, 0.0065852131797276654, 0.0065464630981149213, 
    0.0065019634966602584, 0.0064507493454486128, 0.0063915159934919853, 
    0.0063227260492913296, 0.0062427356290265801, 0.0061499011003441004, 
    0.0060426848967732264, 0.0059197333030210405, 0.0057799540542633121, 
    0.0056225568752426222, 0.0054470960609030563, 0.0052534817410844247, 
    0.0050419906470056883, 0.0048132635034784724, 0.0045683049697937718, 
    0.0043084713092828427, 0.0040354626733406247, 0.0037513156366356217, 
    0.0034583933017866175, 0.0031593794232237038, 0.0028572610813354191, 
    0.0025553109085459172, 0.0022570542083696211, 0.0019662193677143494, 
    0.0016866622543038159, 0.0014222682252383444, 0.0011768275912507513, 
    0.00095389529397855977, 0.00075665109234166546, 0.00058777172300894564, 
    0.00044932555647198924, 0.00034270784144202178, 0.00026860859811858107, 
    0.00022700886644354875, 0.00021720443274061952, 0.00023784694658322912, 
    0.00028698916264997029, 0.00036214565079849183, 0.00046034985632269036, 
    0.0005782188714307814, 0.00071202975309063628, 0.00085781569580107133, 
    0.0010114773845596855, 0.0011689207564085729, 0.0013262002719342538, 
    0.0014796557654671778, 0.0016260380115696066, 0.001762595110237871, 
    0.0018871345696861788, 0.0019980429897754086, 0.0020942826203930887, 
    0.0021753490240250259, 0.0022412145448552708, 0.0022922463086921746, 
    0.0023291141126429047, 0.0023526828301827854, 0.0023639125271163355, 
    0.0023637506425060527, 0.0023530374055300519, 0.002332436575950096, 
    0.0023023880213198285, 0.0022630875785779356, 0.0022145088534514228, 
    0.002156445105618513, 0.0020885797552161718, 0.0020105674076252708, 
    0.0019221236446778206, 0.0018230973495580204, 0.0017135268639707213, 
    0.0015936641269909094, 0.0014639764461055057, 0.00132511186497215, 
    0.0011778545326736429, 0.0010230656142839363, 0.00086162234224481033, 
    0.00069436436136167934, 0.00052205025865598663, 0.0003453314926577959, 
    0.00016474603426418181, -1.9264411870804806e-05, -0.00020632484155957943, 
    -0.00039607744569133789, -0.00058812478109963244, 
    -0.00078197636976220272, -0.00097698864603384386, -0.0011723351669852139, 
    -0.0013669877771134826, -0.0015597301895586405, -0.0017491848089171182, 
    -0.0019338613400790923, -0.0021122057389029499, -0.0022826380946395506, 
    -0.0024435822713591532, -0.0025934861803375646, -0.002730853054399505, 
    -0.0028542979899631987, -0.002962632346939444, -0.0030549769043681494, 
    -0.0031308765384065666, -0.0031903814524670646, -0.003234076641491473, 
    -0.0032630393783472816, -0.0032787538880718918, -0.0032829952921683632, 
    -0.0032777149850890717, -0.0032649323364883956, -0.0032466399628821307, 
    -0.0032247111088986617, -0.0032008187585218211, -0.0031763534891884201, 
    -0.0031523587136517042, -0.0031294708326893893, -0.0031078861177380743, 
    -0.0030873333126832949, -0.003067080563221775, -0.0030459672731114793, 
    -0.0030224606042206729, -0.0029947425427068524, -0.0029608154053132811, 
    -0.0029186233676554416, -0.0028661865331715609, -0.0028017202458119027, 
    -0.0027237450107650807, -0.0026311749978090086, -0.0025233675460281961, 
    -0.0024001430173223991, -0.0022617731194840892, -0.0021089490210206016, 
    -0.0019427401470031467, -0.0017645484607105666, -0.0015760624556870641, 
    -0.0013792288006500338, -0.0011762349257722633, -0.00096949277706926621, 
    -0.00076163043389546709, -0.00055547068969548363, 
    -0.00035401030670888315, -0.00016037045753563949, 2.2267705021029481e-05, 
    0.00019075588517980909, 0.00034208261936654303, 0.00047348946144170506, 
    0.00058259568706194509, 0.00066750500516617184, 0.00072690283066701345, 
    0.00076013455007208444, 0.00076725235097697009, 0.00074904025731626614, 
    0.00070700947585751418, 0.00064337336507784158, 0.0005609894107185409, 
    0.00046326438934990324, 0.00035402112986247032, 0.00023732685774115463, 
    0.00011730273430422459, -2.067295936079047e-06, -0.00011712790040008226, 
    -0.00022470215315913849, -0.00032220477106809694, 
    -0.00040772213211418961, -0.00048004688364945063, 
    -0.00053867191475036379, -0.00058374369880125206, 
    -0.00061598660315634866, -0.00063658998038775493, 
    -0.00064710512689698677, -0.00064933073147137429, 
    -0.00064521967968853759, -0.00063680180874621311, 
    -0.00062613003840847857, -0.00061523071585293566, 
    -0.00060607082880649837, -0.00060051061944951887, 
    -0.00060024914267149784, -0.00060675687178930629, 
    -0.00062120090211096788, -0.00064436799774818579, 
    -0.00067660554485354015, -0.00071778185262064099, 
    -0.00076728022359685171, -0.00082402039584813483, 
    -0.00088651309023234982, -0.00095293678099262077, -0.0010212232657445443, 
    -0.0010891672979406587, -0.0011545371493822476, -0.0012151984484229531, 
    -0.0012692401369703008, -0.0013150870547182923, -0.0013515855774836529, 
    -0.0013780529508303026, -0.0013942854573738017, -0.0014005331094331898, 
    -0.0013974368322323255, -0.0013859441913141284, -0.0013672122635471364, 
    -0.0013424951325661087, -0.0013130453618837186, -0.0012800193119919892, 
    -0.0012443990056862607, -0.0012069369079065434, -0.0011681268533456231, 
    -0.001128182905890339, -0.0010870344555913886, -0.0010443371487130575, 
    -0.00099948268926143319, -0.00095162239241550922, 
    -0.00089970284888114935, -0.00084252023454459873, 
    -0.00077878884277937167, -0.00070721991155178114, 
    -0.00062662321039852096, -0.00053600758163650005, 
    -0.00043468044080994931, -0.00032232705603229661, 
    -0.00019905422124931812, -6.54007610365006e-05, 7.7703430868272414e-05, 
    0.00022901821199801967, 0.00038710025830940038, 0.00055040411258083484, 
    0.00071736645074038478, 0.00088645675445971658, 0.0010561765398849447, 
    0.001225025830645385, 0.0013914345428380347, 0.0015536782669873972, 
    0.0017097880692402371, 0.0018574945795409201, 0.0019941882486030106, 
    0.0021169239958430484, 0.002222468380853878, 0.0023073942523718668, 
    0.0023682144291483202, 0.0024015454183321152, 0.0024042920284093792, 
    0.0023738350768099581, 0.00230819712729643, 0.0022061813540425581, 
    0.0020674679136213122, 0.001892665479512042, 0.0016833056090603078, 
    0.0014417885377030865, 0.0011712862428597129, 0.00087560054559443392, 
    0.00055900186839653821, 0.00022605084873415006, -0.00011857781960116406, 
    -0.00047026382793801264, -0.00082457011989381965, -0.0011773528018646394, 
    -0.0015248342444179992, -0.001863644486338507, -0.002190828770489546, 
    -0.002503835254501683, -0.0028004840076591153, -0.0030789219296755402, 
    -0.0033375765613259875, -0.0035751096934169514, -0.0037903845861940806, 
    -0.0039824536964739865, -0.0041505719360829686, -0.0042942275077437258, 
    -0.0044131919023200697, -0.0045075660799311608, -0.0045778262949954284, 
    -0.0046248475223740456, -0.0046498939307582868, -0.0046545890572479718, 
    -0.0046408537601284666, -0.0046108246610183515, -0.0045667651214501932, 
    -0.0045109733215542161, -0.0044456928256850553, -0.0043730338498368798, 
    -0.0042949154179087812, -0.004213020602319646, -0.0041287621362621268, 
    -0.004043247792360565, -0.0039572363390192392, -0.0038710759554711474, 
    -0.0037846376249930269, -0.0036972561581930089, -0.0036077016064087726, 
    -0.0035142096937752706, -0.0034145590577800465, -0.003306211581108223, 
    -0.0031864904702509785, -0.0030527768029868503, -0.0029027157709192323, 
    -0.0027343985607287415, -0.0025465185282985254, -0.0023384835483255973, 
    -0.0021104734784477518, -0.0018634436949416262, -0.0015990723944326298, 
    -0.0013196668159408294, -0.0010280320559875847, -0.00072731697713166539, 
    -0.00042086275352202639, -0.00011205694538827038, 0.0001957909181283885, 
    0.00049954069763760093, 0.00079628794877842205, 0.001083392897557701, 
    0.0013584814378498099, 0.0016194332265452333, 0.0018643489109840894, 
    0.0020915290420790056, 0.0022994499163420468, 0.002486779943051051, 
    0.0026524031305998307, 0.0027954773801903217, 0.002915497346871384, 
    0.0030123577775875089, 0.003086403716984625, 0.0031384578342746848, 
    0.0031698207691348334, 0.0031822322171741811, 0.0031778052358017463, 
    0.0031589414509945947, 0.0031282344476141685, 0.0030883837881719328, 
    0.0030421020715927028, 0.0029920456530132711, 0.0029407498476482974, 
    0.0028905665286527919, 0.0028435958296128966, 0.0028016429845479094, 
    0.0027661659011094871, 0.0027382404145287207, 0.002718547863311856, 
    0.0027073869517803572, 0.0027047000357823129, 0.002710129610564849, 
    0.0027230830461884006, 0.0027428248914746246, 0.0027685569727699194, 
    0.0027995191919513575, 0.0028350583699581545, 0.0028746607115203559, 
    0.002917951825683282, 0.0029646374923673648, 0.0030144173987511026, 
    0.0030668812312201572, 0.0031214224024121782, 0.0031771681155343362, 
    0.0032329538471993729, 0.003287338596204233, 0.0033386551370177646, 
    0.0033850905302274872, 0.0034247886028495934, 0.0034559668302276067, 
    0.0034770434562218294, 0.0034867624965301269, 0.0034843034894025066, 
    0.0034693688524078813, 0.00344222958554544, 0.0034037137923756413, 
    0.0033551541922539649, 0.0032982759103328731, 0.0032350441115398553, 
    0.0031674830591402799, 0.0030974945925548595, 0.0030266857539803767, 
    0.0029562321640131668, 0.0028867916983744669, 0.0028184772606947061, 
    0.0027508818897121648, 0.0026831600993306361, 0.0026141600410623401, 
    0.0025425838100558863, 0.0024671687042623468, 0.0023868797030996724, 
    0.0023010829497150708, 0.0022096913712171028, 0.0021132601826270095, 
    0.0020130110239184431, 0.0019107991991521413, 0.0018090125141367428, 
    0.0017104193172168838, 0.0016179849200642952, 0.0015346679673821947, 
    0.0014632219744513026, 0.0014060183784409949, 0.0013648975517166692, 
    0.0013410673433694096, 0.0013350450276140794, 0.0013466485081705234, 
    0.0013750302027752601, 0.0014187436026453684, 0.0014758285968353082, 
    0.0015439146475362715, 0.0016203207467212059, 0.0017021543786437147, 
    0.0017864121961532347, 0.0018700731736181531, 0.0019501952695403506, 
    0.002024017790134332, 0.0020890710914552033, 0.0021432846216993327, 
    0.0021850935825096156, 0.0022135290291830068, 0.0022282700977312607, 
    0.0022296465877511434, 0.0022185737153622119, 0.0021964400901236477, 
    0.0021649639856170092, 0.0021260219126687384, 0.0020814738631594349, 
    0.0020330192104939778, 0.0019820897927367697, 0.0019297764237877584, 
    0.0018768217559834615, 0.0018236518523249551, 0.0017704499056252299, 
    0.0017172615630608623, 0.0016641001379942265, 0.001611055970081509, 
    0.0015583693174210708, 0.0015064631795728986, 0.0014559388820937092, 
    0.0014075183721038256, 0.0013619516539651183, 0.0013198939786029395, 
    0.0012817753609845872, 0.0012476866734716689, 0.0012172860608510431, 
    0.0011897456305224189, 0.0011637610066564774, 0.0011376127190565366, 
    0.0011092842660711173, 0.0010766458013049705, 0.0010376536761126658, 
    0.00099057962220349175, 0.00093422235441816557, 0.00086808149770481208, 
    0.00079247083307049549, 0.00070855740673014269, 0.00061832385747760514, 
    0.00052445409971416091, 0.00043016248956749098, 0.00033897071767052638, 
    0.00025446341866532259, 0.00018002178568498725, 0.00011856982084390842, 
    7.2354367232238439e-05, 4.2763827773892783e-05, 3.0202520734189391e-05, 
    3.4035691064756223e-05, 5.2592533875122212e-05, 8.3243035975189328e-05, 
    0.00012252686968810557, 0.00016635032724765801, 0.00021021665489396555, 
    0.00024948944359318821, 0.00027964688022470924, 0.00029652929643368448, 
    0.00029654931344965307, 0.00027686662538639736, 0.00023551790646570217, 
    0.00017150175970387171, 8.4799935949740466e-05, -2.3658896131942709e-05, 
    -0.00015209663374037084, -0.00029803677964060501, 
    -0.00045849439612598216, -0.00063020002519777402, 
    -0.00080981391624552156, -0.00099413378076606954, -0.0011802598147567366, 
    -0.0013657113281723772, -0.0015484860608749149, -0.0017270602844892762, 
    -0.0019003438013299959, -0.0020675933117056461, -0.0022283239129453456, 
    -0.0023822150387719466, -0.0025290270372596204, -0.0026685420166848166, 
    -0.0028005192600557239, -0.002924670782971235, -0.0030406393101721158, 
    -0.0031479943540973954, -0.003246230260796062, -0.0033347629218310609, 
    -0.0034129315403883254, -0.0034799872475610606, -0.0035350822209157177, 
    -0.0035772528416133111, -0.0036054048581905499, -0.0036183316899331928, 
    -0.0036147489799261334, -0.0035933813197194715, -0.0035530656336879452, 
    -0.0034928773487457143, -0.0034122636493664205, -0.0033111536321653451, 
    -0.0031900403770311983, -0.003050017151574744, -0.0028927711303270718, 
    -0.0027205289383308742, -0.002535968782895436, -0.0023421090383590856, 
    -0.0021421779367307922, -0.0019394835236798682, -0.0017372811145090782, 
    -0.0015386419787464553, -0.0013463357255313771, -0.0011627230687152876, 
    -0.0009896735047021034, -0.00082850710426480016, -0.00067996670099028302, 
    -0.00054423559160701577, -0.00042097891605724256, 
    -0.00030943724888462452, -0.00020853266038153715, 
    -0.00011701768440295203, -3.3615205954794339e-05, 4.2844415444000272e-05, 
    0.00011331262275758841, 0.00017844680008434157, 0.00023857778174881454, 
    0.00029371341338383804, 0.00034358046928510688, 0.00038767959847902663, 
    0.00042534566761082609, 0.00045581551206993191, 0.00047828228071178228, 
    0.00049194495921156642, 0.00049605191374796202, 0.00048993183541947588, 
    0.00047302181733034361, 0.00044487872903629304, 0.00040517371507634687, 
    0.00035369240787122254, 0.00029032321477825756, 0.00021505584833205718, 
    0.00012797696328717282, 2.9285680232746854e-05, -8.0702140884164131e-05, 
    -0.00020153664605502132, -0.00033261297655350747, 
    -0.00047314704770077751, -0.00062215022558162383, 
    -0.00077839980548678788, -0.00094040950052868525, -0.0011064115692373897, 
    -0.0012743503576576171, -0.0014418989199200445, -0.0016065002982846557, 
    -0.0017654330588399302, -0.0019159131051156332, -0.0020552160878248619, 
    -0.0021808006075077439, -0.0022904335560744431, -0.0023822883790975743, 
    -0.0024550235964933284, -0.002507820121321001, -0.0025403799655022751, 
    -0.0025528913948947422, -0.0025459748697144028, -0.0025206069455639777, 
    -0.0024780462113955797, -0.0024197869084877986, -0.0023475399522381629, 
    -0.002263257865523225, -0.0021691899716973673, -0.0020679352642458139, 
    -0.0019624940019439293, -0.0018562685703478604, -0.0017530230011183999, 
    -0.0016567805323862575, -0.0015716687813483669, -0.0015017156761407359, 
    -0.001450624433506716, -0.0014215429508924505, -0.0014168590159915947, 
    -0.0014380528189017728, -0.001485603317498667, -0.0015589696350860626, 
    -0.001656638798058661, -0.0017762113114532544, -0.0019145319447583958, 
    -0.0020678279323373054, -0.0022318551038792316, -0.0024020516094575895, 
    -0.0025736947953065945, -0.0027420508015436273, -0.0029025136411649668, 
    -0.0030507395261373535, -0.003182752482665455, -0.0032950321563951228, 
    -0.0033846072127696708, -0.00344913416587153, -0.0034870050787195821, 
    -0.003497435509274247, -0.0034805653614643633, -0.0034375071529261433, 
    -0.0033703573853059794, -0.0032821576502157813, -0.0031768135705806809, 
    -0.0030589660175032356, -0.0029338460472826994, -0.0028070995902666272, 
    -0.0026846011040393214, -0.002572261527270977, -0.0024758225566896088, 
    -0.0024006679085263804, -0.0023516314388103148, -0.00233281302989932, 
    -0.0023474232932550409, -0.0023976388432846774, -0.0024845115142406028, 
    -0.0026079241454528088, -0.0027666136857133709, -0.0029582438753867411, 
    -0.0031795211681925973, -0.0034263369294174548, -0.0036939123545926627, 
    -0.0039769401061014314, -0.0042697023447230455, -0.0045661806273464131, 
    -0.0048601637770212909, -0.0051453644738361781, -0.0054155502212650669, 
    -0.0056647078834377983, -0.0058872326962592456, -0.0060781247971909303, 
    -0.0062331815811782557, -0.0063491676012283529, -0.0064239418947782392, 
    -0.0064565374016534822, -0.0064471889104039176, -0.0063973153997386144, 
    -0.0063094759339067568, -0.0061872863549691315, -0.0060352968662893258, 
    -0.0058588290780820142, -0.0056637631740843958, -0.0054562841856902319, 
    -0.0052426003590800262, -0.0050286589036389944, -0.0048198907168977888, 
    -0.0046209931748528218, -0.0044357725673465857, -0.0042670397178384851, 
    -0.0041165537328629988, -0.0039850061127098971, -0.0038720331152618361, 
    -0.0037762611046914013, -0.0036953637877576761, -0.0036261446671706568, 
    -0.0035646410590027162, -0.0035062452251396776, -0.0034458553866422658, 
    -0.003378047920983218, -0.0032972711439413342, -0.0031980637018877733, 
    -0.0030752823688807332, -0.0029243322699667763, -0.0027413895146361274, 
    -0.0025235947787003751, -0.002269201101010396, -0.0019776796014406074, 
    -0.0016497661196520253, -0.0012874686232243544, -0.00089403105357115131, 
    -0.00047384812064181524, -3.2361998867955319e-05, 0.00042408345751057582, 
    0.00088843149949645382, 0.0013531208271774788, 0.0018103347207967292, 
    0.0022522499450078337, 0.0026712934565424574, 0.003060391213981059, 
    0.003413186158841583, 0.0037242138677009012, 0.0039890344597085471, 
    0.0042043087466707907, 0.0043678242785709902, 0.0044784730117614678, 
    0.0045361981711277144, 0.0045419138348441641, 0.0044974086016765077, 
    0.0044052418556154395, 0.004268638942972732, 0.004091375783695346, 
    0.0038776682440348894, 0.0036320494529418035, 0.0033592413447894862, 
    0.0030640367913606615, 0.002751198737838665, 0.0024253846122642159, 
    0.0020910968998774436, 0.0017526716356265648, 0.001414275087189897, 
    0.0010799115436265633, 0.00075340594369651553, 0.00043838697426864235, 
    0.00013823066995989156, -0.00014400358418093379, -0.00040567679407889346, 
    -0.00064466935896935723, -0.0008594837267078679, -0.0010493292551536171, 
    -0.0012141813725389233, -0.0013548018149970669, -0.0014727251972752084, 
    -0.001570190782268779, -0.0016500498955809618, -0.0017156162165744618, 
    -0.0017704962468405769, -0.0018183718612421436, -0.0018627866006207447, 
    -0.0019069014281742364, -0.001953287474972669, -0.0020037348704116291, 
    -0.002059127799623155, -0.0021193785249118704, -0.002183445055200032, 
    -0.0022494062097123966, -0.002314598725964883, -0.0023757822330217754, 
    -0.0024293270850864724, -0.0024714002205559714, -0.0024981407097790093, 
    -0.002505815140352077, -0.002490953462747469, -0.0024504516246190299, 
    -0.0023816476587479301, -0.002282368178375131, -0.0021509685121862097, 
    -0.0019863649721775182, -0.0017880669103034091, -0.0015562189148981879, 
    -0.0012916271312407679, -0.00099577334180504101, -0.00067078768804427157, 
    -0.00031938486873418271, 5.5241131806362084e-05, 0.00044954675325460018, 
    0.00085975769673549802, 0.0012819617970793549, 0.0017121511243615578, 
    0.002146226361077524, 0.002579961980709279, 0.0030089745916854539, 
    0.003428698121596325, 0.0038343814490075729, 0.0042211272024563779, 
    0.0045839558191763351, 0.0049179110209424167, 0.0052181827202011834, 
    0.0054802450540447304, 0.0056999837460834464, 0.0058738309465606632, 
    0.0059988757234486403, 0.0060729542874227854, 0.0060947230305167218, 
    0.0060636963876816259, 0.005980265156309659, 0.0058456944989116986, 
    0.0056621024228682929, 0.0054324028936732867, 0.0051602252520121837, 
    0.0048498224472958784, 0.0045059628953265252, 0.0041338184488800564, 
    0.0037388534276892125, 0.0033267137489131986, 0.0029031308395130254, 
    0.0024738171151515265, 0.0020443765659032154, 0.001620209767665474, 
    0.0012064184096809494, 0.00080770359614606242, 0.00042825816758199612, 
    7.1661878228555705e-05, -0.00025920760820621381, -0.00056222162025696201, 
    -0.00083601328078722239, -0.0010799478138872828, -0.001294048854536759, 
    -0.0014789269850016234, -0.0016357057299336768, -0.0017659560536301177, 
    -0.0018716404979226486, -0.0019550765643854568, -0.0020189028165245454, 
    -0.0020660514282084728, -0.0020997028629041749, -0.0021232347006001342, 
    -0.002140155134901556, -0.0021540167908896354, -0.0021682982442798814, 
    -0.0021862820344341464, -0.0022109397865570858, -0.0022448063045393215, 
    -0.0022898783874337578, -0.0023475470588306467, -0.0024185449632349448, 
    -0.0025029375878921692, -0.0026001400506635722, -0.002708982190846909, 
    -0.002827775353115456, -0.0029543991024589028, -0.0030863950933233126, 
    -0.0032210536289326648, -0.0033554997613613993, -0.0034867753710273413, 
    -0.003611909785344944, -0.003727998238513692, -0.0038322644883173889, 
    -0.0039221329209734122, -0.0039952953553714782, -0.0040497629523728648, 
    -0.0040839124686523438, -0.004096528885356927, -0.0040868211983272271, 
    -0.0040544487435414415, -0.0039995148484721172, -0.0039225676983450017, 
    -0.0038245771855597382, -0.0037068718735334249, -0.0035710650256777754, 
    -0.0034189464006851534, -0.0032523597515845032, -0.0030730703612509148, 
    -0.0028826588567812577, -0.0026824358863268716, -0.0024734028309140342, 
    -0.0022562595969639982, -0.0020314615424792356, -0.0017993003320578829, 
    -0.0015600196189175619, -0.0013139170390171241, -0.0010614449344864669, 
    -0.00080327438226540789, -0.00054031347519104878, 
    -0.00027369186343452403, -4.7089629121817354e-06, 0.00026523722040473313, 
    0.00053471164985085422, 0.00080227157185868716, 0.0010664754430607716, 
    0.001325845532874944, 0.0015788102388773089, 0.0018236416022922295, 
    0.0020583968437110486, 0.0022808713469291931, 0.002488593311838381, 
    0.0026788433983640269, 0.0028487285066913547, 0.0029953097660925586, 
    0.0031157654345043886, 0.0032075975639417327, 0.0032688458390905967, 
    0.0032983116740617612, 0.0032957500048470816, 0.0032620051131645568, 
    0.003199090594546491, 0.0031101752253169111, 0.002999480881295054, 
    0.0028720959789365536, 0.0027337089783803807, 0.0025902841679198061, 
    0.002447726040372444, 0.0023115515551726381, 0.0021865963852265424, 
    0.0020767731579797184, 0.001984920294464856, 0.0019127068886591726, 
    0.0018606373103012546, 0.001828110019924099, 0.001813537807121754, 
    0.0018145136305979038, 0.0018280041405645854, 0.0018505707754087766, 
    0.0018785824302740054, 0.0019084556966251713, 0.0019368771888769749, 
    0.0019610315565253712, 0.0019788074050617671, 0.0019889729441077506, 
    0.0019913078995525296, 0.0019866682375525436, 0.0019769824282639971, 
    0.0019651548787101023, 0.0019548881016937568, 0.0019504106397889647, 
    0.0019561503428296204, 0.001976373127935427, 0.0020148149402132217, 
    0.0020743552047849732, 0.0021567524063849882, 0.0022624470735923717, 
    0.0023904574173565256, 0.0025383460452195012, 0.0027022690024464291, 
    0.0028771224477612111, 0.0030567679094699583, 0.0032343673730131591, 
    0.003402776105290291, 0.0035549667309604707, 0.0036844339183172165, 
    0.0037855376825226749, 0.0038537473326205329, 0.0038858122646080297, 
    0.0038798242958329255, 0.0038352107169066698, 0.0037526650277310185, 
    0.0036340188472917135, 0.0034820718207197151, 0.0033003729233681981, 
    0.0030929787713153164, 0.0028642123898726759, 0.002618424559993485, 
    0.002359815230379429, 0.0020922965815390565, 0.001819407287987566, 
    0.0015442642848349437, 0.0012695741786356214, 0.00099764472806979435, 
    0.00073044577950941332, 0.00046965993600141601, 0.00021675611039649449, 
    -2.6946181123171931e-05, -0.00026021813360435088, 
    -0.00048188393288953104, -0.00069079526397043775, 
    -0.00088582144562608742, -0.0010658733441071303, -0.0012299375969632401, 
    -0.0013771378098708512, -0.0015068035149251925, -0.001618536120257922, 
    -0.0017123016331942603, -0.0017884923070935429, -0.0018479895566655502, 
    -0.0018922145539423678, -0.0019231612691922527, -0.0019434209138699168, 
    -0.0019561933406878769, -0.0019652808505363295, -0.0019750266754457384, 
    -0.00199022875836561, -0.0020159920740599677, -0.0020575275573416324, 
    -0.0021199020410733712, -0.0022077443490476864, -0.0023249569890318013, 
    -0.0024744318393432594, -0.002657830652945831, -0.0028754639692740096, 
    -0.0031263138399694849, -0.0034081897642889735, -0.0037180104837162106, 
    -0.0040521392234204373, -0.004406721371641705, -0.0047779332844172743, 
    -0.0051621372699497134, -0.0055559071646327073, -0.0059559935964395121, 
    -0.0063592560396720614, -0.0067625943469939312, -0.0071629066791053762, 
    -0.0075570505912005096, -0.007941826704561868, -0.0083139542331882536, 
    -0.0086700809392874657, -0.0090067905272548758, -0.0093206339069325534, 
    -0.0096081929796124361, -0.0098661486982943528, -0.010091390932839471, 
    -0.010281117999806088, -0.010432944147194034, -0.01054500999145958, 
    -0.010616071860911923, -0.01064556924490625, -0.010633642137615392, 
    -0.01058111886490321, -0.010489456272580945, -0.010360641356160617, 
    -0.010197060712216549, -0.010001358906422576, -0.0097762956435845337, 
    -0.0095246067560869584, -0.0092489099471495268, -0.0089516355500550981, 
    -0.0086349993120745441, -0.0083010281133232503, -0.0079515903102328929, 
    -0.0075884541510860886, -0.0072133461178480488, -0.0068280190286219055, 
    -0.0064343024179287127, -0.0060341644279387563, -0.0056297506463522436, 
    -0.0052234194886848599, -0.0048177510405928011, -0.0044155287595865744, 
    -0.0040196838738831408, -0.0036332229993191849, -0.0032591312928175169, 
    -0.0029002602303283796, -0.002559222288267536, -0.0022382902606200086, 
    -0.0019393234501858152, -0.0016637243924273806, -0.0014124175781096951, 
    -0.0011858596593599684, -0.00098405532870068555, -0.00080659086774934963, 
    -0.00065265676215738456, -0.00052108275965353937, 
    -0.00041035418227122544, -0.00031864425324091487, 
    -0.00024383824756687121, -0.00018355913565888519, 
    -0.00013521078709269443, -9.6003058128239739e-05, 
    -6.2998337968385356e-05, -3.3164095433179178e-05, 
    -3.4554906544564902e-06, 2.9080263746196012e-05, 6.7175629483250728e-05, 
    0.00011321963873177636, 0.00016913756718224256, 0.00023629335349128686, 
    0.00031543486783820827, 0.00040668418798566223, 0.0005095720007961017, 
    0.0006231129289648652, 0.00074593935439958231, 0.00087642550594314514, 
    0.001012816418373257, 0.0011533278968047507, 0.0012962061859860922, 
    0.001439737017302893, 0.001582214896376903, 0.0017218832341066052, 
    0.0018568597883501878, 0.0019850682489060746, 0.0021042077006029444, 
    0.0022117634885818883, 0.0023050718608696448, 0.0023814508132458463, 
    0.002438355094316791, 0.0024735420446674312, 0.0024852206676393837, 
    0.0024721601545298596, 0.0024337489018309453, 0.0023699964262225708, 
    0.0022815344320011293, 0.0021695811405474802, 0.0020359243283879095, 
    0.0018828821080588956, 0.0017132633947908168, 0.0015303249727025231, 
    0.001337700040289532, 0.0011392932447975676, 0.00093916889499160913, 
    0.00074140589138718183, 0.00054996724261366934, 0.00036860204336604371, 
    0.00020077801748406436, 4.9654633585750484e-05, -8.1939520185730946e-05, 
    -0.00019153483860148671, -0.00027707785906404259, 
    -0.00033702186835101372, -0.00037042708282364686, 
    -0.00037705581226761385, -0.00035743724111451225, 
    -0.00031287870459988939, -0.00024538724118108391, 
    -0.00015755818908322114, -5.241986763462944e-05, 6.6722361128493296e-05, 
    0.00019641250411030399, 0.00033312287320039441, 0.00047328035241625473, 
    0.00061326246249273741, 0.0007494069018197237, 0.00087802616244579289, 
    0.00099548329866524284, 0.0010982766886681939, 0.0011831490175053141, 
    0.0012471876908695374, 0.0012878729775142226, 0.0013030959349394366, 
    0.0012911332414022615, 0.0012506357619565891, 0.0011806359955876945, 
    0.0010805825533798941, 0.00095039815993296702, 0.00079053748627410834, 
    0.00060204617322943445, 0.00038658497675035452, 0.00014644774116367911, 
    -0.00011545494252780469, -0.00039562325513382152, 
    -0.00068999569052976021, -0.00099399418616750827, -0.0013025633127844547, 
    -0.0016102551481754228, -0.0019113205229327516, -0.0021998573216676252, 
    -0.0024699758822153885, -0.0027159603852859931, -0.0029324334327979402, 
    -0.0031144911874906186, -0.003257831554362245, -0.0033589058751199298, 
    -0.0034150860247035078, -0.0034248478152063659, -0.0033879299177662515, 
    -0.003305443650205716, -0.0031798891449044474, -0.0030150323897615776, 
    -0.002815669011002068, -0.0025873223779017017, -0.0023359476988666218, 
    -0.0020676648343316904, -0.001788542564611036, -0.0015044088638816191, 
    -0.0012207118240433997, -0.00094239268279135689, -0.00067379134220662889, 
    -0.00041855904017580126, -0.0001795910314117508, 4.0998356561540699e-05, 
    0.00024185678986146631, 0.00042231075479199097, 0.00058222709672460233, 
    0.00072182454337770333, 0.00084149259566558608, 0.00094160299030422419, 
    0.0010223603826502636, 0.001083686984536544, 0.001125162108823351, 
    0.0011460154834274968, 0.0011451661122034245, 0.0011213241754781059, 
    0.0010730733504631647, 0.00099899516514021652, 0.00089774880565940494, 
    0.00076819959097877526, 0.00060957431148642735, 0.00042169585484937958, 
    0.00020522960293724692, -3.8068135920247539e-05, -0.00030516750960453204, 
    -0.00059172035916692256, -0.00089212284924934139, -0.0011997372731042566, 
    -0.0015072055254743981, -0.0018068249922771548, -0.0020909554704953131, 
    -0.002352364995060364, -0.002584552444126796, -0.002781995661419913, 
    -0.0029403139116080455, -0.0030563435760817457, -0.003128156047007071, 
    -0.0031549901224872923, -0.0031371446749271946, -0.0030758327550346526, 
    -0.0029730287989425024, -0.0028313149530332041, -0.0026537426465658397, 
    -0.0024437052848966636, -0.0022048341833231016, -0.001940931259031132, 
    -0.0016558970145300999, -0.0013536907622367274, -0.0010382962121266981, 
    -0.00071368599532936681, -0.00038378488773507932, 
    -5.2400096407263073e-05, 0.00027685497976312831, 0.00060063394159732978, 
    0.00091592010680890317, 0.0012200835412615597, 0.0015109022747825586, 
    0.0017865568890269689, 0.0020455967213318087, 0.0022869160632658465, 
    0.0025097337941343916, 0.0027135731939913988, 0.0028982813839838737, 
    0.0030640466453930445, 0.0032114071316341024, 0.0033412245844910214, 
    0.0034546368262710651, 0.0035529803980772841, 0.0036376922755940069, 
    0.0037102119995920473, 0.0037719057795962577, 0.0038240000907058848, 
    0.0038675465030787036, 0.0039034173285549317, 0.0039323305993999086, 
    0.0039549446589931068, 0.0039720151923370479, 0.0039845332509095572, 
    0.0039938586359421326, 0.0040017585004397116, 0.004010404404624063, 
    0.0040222746782957244, 0.0040400167964467822, 0.0040662644822285904, 
    0.0041034581826770462, 0.0041536368514735441, 0.0042182837768709579, 
    0.0042981556745522488, 0.0043931912983414846, 0.0045024556622054396, 
    0.00462415980530732, 0.0047557568928676989, 0.0048940710413767786, 
    0.0050354849513096003, 0.0051761298262345858, 0.0053120956906679007, 
    0.0054396308886577429, 0.0055553480107604627, 0.0056564020104146176, 
    0.0057406573930338005, 0.0058068529639158312, 0.0058547186777793327, 
    0.0058850444584285884, 0.0058997062339356272, 0.0059015855407849455, 
    0.0058944065454844662, 0.005882489408023734, 0.0058704625518815967, 
    0.0058629158884994162, 0.0058641191557917633, 0.005877733851417339, 
    0.0059066290691889168, 0.0059527302299731289, 0.0060169318397036171, 
    0.006099051524461419, 0.0061978258155664665, 0.0063109683838268324, 
    0.0064352463133547757, 0.0065666073057076002, 0.0067003769055141663, 
    0.0068314744426823384, 0.0069546724805220946, 0.0070648771210770544, 
    0.0071573752978835682, 0.0072280200760249796, 0.0072734062628158069, 
    0.0072909111745539839, 0.0072787528272130753, 0.0072359418894898751, 
    0.007162195066189361, 0.0070578191426883524, 0.0069235971341525659, 
    0.0067607084815357078, 0.0065706460242547487, 0.0063551667534909378, 
    0.0061162041931868529, 0.0058557509853981431, 0.0055757776368769206, 
    0.0052781701459423932, 0.0049647300271372695, 0.0046372326912826958, 
    0.0042975108930280491, 0.0039475381545026429, 0.0035894628680512323, 
    0.0032256370309735527, 0.0028585364773737686, 0.0024906303757171642, 
    0.0021242280418480607, 0.0017613185056993079, 0.0014034281353938229, 
    0.0010515432536771048, 0.00070606202805282539, 0.0003668447198124172, 
    3.3297154054868691e-05, -0.00029551409412684903, -0.00062076212738657326, 
    -0.00094373398700203434, -0.0012657211567649194, -0.0015878988489614429, 
    -0.0019111862609785138, -0.0022360798703139769, -0.0025624795071759136, 
    -0.002889524332021917, -0.0032154738490844737, -0.003537665071433499, 
    -0.0038525948941354198, -0.0041560911247466078, -0.0044435639899253554, 
    -0.0047102586883212422, -0.0049515614410446619, -0.0051632453109293755, 
    -0.0053417386432191329, -0.0054843543477456616, -0.0055894760500792571, 
    -0.0056566263719487744, -0.0056864579452735988, -0.0056806423621320783, 
    -0.0056417019654985906, -0.0055727919094717502, -0.0054775316349016077, 
    -0.0053598438465271379, -0.0052238787642497845, -0.0050739689365026045, 
    -0.0049146156334332336, -0.0047504662864990199, -0.004586238933686094, 
    -0.0044266223087018964, -0.0042761431574152575, -0.0041389785907565476, 
    -0.0040187623333803801, -0.0039183845386167445, -0.0038398362313689402, 
    -0.0037840571567965523, -0.0037508810464070069, -0.0037390316154381725, 
    -0.003746191862642685, -0.003769184318304101, -0.0038041955523696325, 
    -0.0038470777115039369, -0.0038936948679038851, -0.0039403128258356903, 
    -0.0039839135811598142, -0.0040225037168163114, -0.0040553092244231797, 
    -0.0040828994348490067, -0.0041072027158346857, -0.0041314024286534037, 
    -0.0041597615613072781, -0.0041973371284180268, -0.0042496792801396763, 
    -0.0043225040479110289, -0.0044212961667206745, -0.0045509167650714987, 
    -0.0047152045429884075, -0.0049165304133744619, -0.0051554321871183197, 
    -0.0054303508091966771, -0.0057375592933361502, -0.0060712277508696783, 
    -0.0064236415922821121, -0.0067855307906108699, -0.0071464209894138006, 
    -0.0074950676478153623, -0.0078198894283424813, -0.0081094590131290094, 
    -0.0083529952567100892, -0.0085408351705162072, -0.0086648713188960235, 
    -0.0087189077242687731, -0.0086989086985083518, -0.0086030605938730888, 
    -0.0084317395518972334, -0.0081873179147387148, -0.0078739531914674976, 
    -0.007497324026799152, -0.0070643874050081738, -0.0065831810271338468, 
    -0.0060626645681951998, -0.0055125918108750154, -0.004943353908537197, 
    -0.0043658394184781192, -0.0037912019117518213, -0.0032306405519646666, 
    -0.0026951615004360916, -0.0021953448214431385, -0.0017411901961599421, 
    -0.0013419873366067989, -0.0010062550495264981, -0.00074166116994085448, 
    -0.00055489729966985203, -0.00045153475379267126, -0.000435808561787454, 
    -0.00051037336202222204, -0.00067604073054084953, 
    -0.00093154688305107291, -0.0012734013534601316, -0.0016958256632871749, 
    -0.0021907466759381162, -0.0027479137069342466, -0.0033551539823837347, 
    -0.0039986830554147382, -0.0046635170631469571, -0.0053339216374958132, 
    -0.0059939375854260657, -0.0066278830982016311, -0.007220865952789729, 
    -0.0077592293958841912, -0.0082309399853876721, -0.0086259171541440867, 
    -0.0089362860807766266, -0.0091566041398165997, -0.0092839605569856164, 
    -0.0093180528475703822, -0.0092611495373680526, -0.0091179658909780869, 
    -0.0088954254183781275, -0.0086023333996348948, -0.0082490087193407072, 
    -0.0078468619515473324, -0.0074079923142256962, -0.0069447838119927824, 
    -0.0064695385342859943, -0.0059941076830351079, -0.0055295105761241602, 
    -0.0050855455464118276, -0.0046703781377242523, -0.0042900960490505104, 
    -0.0039483434781801162, -0.0036460441694337415, -0.0033812738315427749, 
    -0.0031493344359800513, -0.0029430486013741412, -0.0027532517784045873, 
    -0.0025694258972383038, -0.0023805165426712066, -0.0021757397433226841, 
    -0.0019454389305177144, -0.001681787543981228, -0.001379425848935401, 
    -0.0010357989171725047, -0.00065133885969742436, -0.00022939582802789581, 
    0.00022400970152354789, 0.00070061488491456676, 0.0011904692675301608, 
    0.0016825967088132856, 0.0021656706232433625, 0.0026286994243692346, 
    0.0030616045357502652, 0.0034557542842594867, 0.0038043556388458444, 
    0.0041026507850320405, 0.0043479354537225273, 0.0045394984021911609, 
    0.0046783532281087807, 0.0047669363884511404, 0.0048087399361776756, 
    0.0048080011284705919, 0.004769427258441125, 0.0046979676973027389, 
    0.0045986348643702523, 0.004476328089050143, 0.0043355960814100659, 
    0.0041804175718711256, 0.0040140181514415419, 0.0038388125367891002, 
    0.0036564168792318384, 0.003467808403206281, 0.0032734936402220903, 
    0.0030735930248939917, 0.0028678787205086631, 0.0026557731681180782, 
    0.0024362960101026922, 0.0022080801230000718, 0.0019694469395287332, 
    0.001718552239612159, 0.0014535745852172492, 0.0011729554330885987, 
    0.00087559653706436626, 0.00056099661881218099, 0.0002292844859618187, 
    -0.00011878577100438181, -0.00048190308033275249, 
    -0.00085830027098596803, -0.0012458937709385017, -0.0016424577554907012, 
    -0.0020458065008774227, -0.0024539874654898384, -0.002865405545498567, 
    -0.0032787866968061259, -0.0036930666566128089, -0.0041071635408730014, 
    -0.0045196459896476981, -0.0049283721320432482, -0.0053301792989888129, 
    -0.0057206582302892425, -0.0060940694163632673, -0.0064433595513082968, 
    -0.0067602924695976648, -0.0070357000280052038, -0.0072598866574406871, 
    -0.0074231419827773312, -0.0075162693235761831, -0.0075312016997711295, 
    -0.0074615012458712198, -0.0073028352671378428, -0.0070533014483204074, 
    -0.0067135142166575863, -0.0062866459123608999, -0.0057782005965857407, 
    -0.0051957374401644524, -0.0045484604350968672, -0.0038468591322241047, 
    -0.0031023328809768949, -0.0023269073256419236, -0.0015330868804501112, 
    -0.00073371331679423254, 5.8069176532051132e-05, 0.00082892817285087341, 
    0.001565350792140163, 0.0022537694477746044, 0.0028807179504243587, 
    0.0034330609816665297, 0.0038983677428624589, 0.0042652929324903267, 
    0.004524059921059892, 0.0046669062842866257, 0.0046884768512136001, 
    0.0045860846544168547, 0.0043598618657735549, 0.0040127107492448928, 
    0.0035501338899773935, 0.0029799068595946234, 0.0023116226876017214, 
    0.0015563259306174816, 0.00072602912398902868, -0.00016662078896159053, 
    -0.001108626980726272, -0.0020867643405582978, -0.003087609909991264, 
    -0.0040973629631083433, -0.0051016393967588123, -0.0060853318186417102, 
    -0.0070327664259342863, -0.0079281751981204636, -0.0087566261920434488, 
    -0.0095050884065880081, -0.010163372415065514, -0.010724848716899616, 
    -0.011186679214811897, -0.01154972269876668, -0.011818048117805357, 
    -0.011998161847640807, -0.012098116843464032, -0.012126593663577349, 
    -0.012092035698829565, -0.012002107074582409, -0.011863410386713395, 
    -0.011681456539949616, -0.01146095070137999, -0.011206226569227491, 
    -0.010921733376633653, -0.010612616473962555, -0.010285079453769086, 
    -0.0099466873302535667, -0.0096064251043711732, -0.0092745973062107103, 
    -0.0089624396186667472, -0.0086817166846242192, -0.0084441480051300911, 
    -0.0082608844878178083, -0.0081420247589419417, -0.0080961977647318172, 
    -0.0081303879294991176, -0.0082497683831827661, -0.0084576316950586497, 
    -0.0087553554960053924, -0.0091423012070975754, -0.0096155944205803222, 
    -0.01017006374291171, -0.010797889884065652, -0.011488449751289686, 
    -0.012228084148457947, -0.012999976095634603, -0.013784246737066722, 
    -0.014558198720703932, -0.015296821883146315, -0.015973577674097468, 
    -0.016561381534726374, -0.01703360477755788, -0.017364960307063006, 
    -0.017532371267580418, -0.017515551719095451, -0.017297523871045221, 
    -0.016865201949754244, -0.016209738480418925, -0.015327002366205799, 
    -0.014217960991238739, -0.01288889490663757, -0.011351325841083207, 
    -0.0096217292593745781, -0.0077209108392324761, -0.0056732959497117902, 
    -0.0035062231108659555, -0.0012492253387137789, 0.0010665540212746153, 
    0.0034089530925620589, 0.00574527707295781, 0.0080430460186122401, 
    0.010270749126575924, 0.012399065044424278, 0.014402045757949938, 
    0.016258435643023511, 0.017952681286184411, 0.019475588877595387, 
    0.020824219318199326, 0.022001021294438448, 0.023012500054898605, 
    0.023867433517888136, 0.024575272688657009, 0.025144843228803049, 
    0.02558313069806321, 0.025894651858578855, 0.026081044314827384, 
    0.026141196172186576, 0.026071764140431587, 0.025867648661968997, 
    0.02552293251764615, 0.025031615166392924, 0.024388446541727685, 
    0.023589518596748467, 0.022633072396166746, 0.021519976656139802, 
    0.020254168841835687, 0.018842545265206269, 0.017294688540078811, 
    0.015622025770935868, 0.013837678419216176, 0.011956370636851744, 
    0.0099950940460827222, 0.0079736897646247775, 0.0059143374115948498, 
    0.0038405856442491606, 0.0017754625617100942, -0.00025981100115550146, 
    -0.0022468387958390862, -0.0041710235944088913, -0.0060207565368462614, 
    -0.0077864131728670885, -0.0094591604694364128, -0.011028994655843484, 
    -0.012482944931472513, -0.013804374420575883, -0.014972593642751299, 
    -0.01596379775960851, -0.016752982514562115, -0.017315865942172631, 
    -0.017633912914645184, -0.017693714317613095,
  // Fqt-F(6, 0-1999)
    0.99999999999999989, 0.99451963138113297, 0.97829897628159479, 
    0.95198395040629702, 0.91659592926405864, 0.87345432023942238, 
    0.82408183826449855, 0.77010316978952975, 0.71314730676179983, 
    0.65476203995077731, 0.59634641256102827, 0.53910398607755583, 
    0.48401704736364753, 0.43183969573030478, 0.38310638753850706, 
    0.33815179752309615, 0.29713779716178929, 0.26008385266803624, 
    0.22689775115934183, 0.19740441199093833, 0.17137141833004851, 
    0.14853051644669699, 0.12859495381584182, 0.11127291199075344, 
    0.096277510868012714, 0.083334012368418559, 0.072184737268829013, 
    0.062592229635505425, 0.054341051753393391, 0.047238505194227821, 
    0.041114557708494232, 0.035821097348283079, 0.031230708899714011, 
    0.027235057039517268, 0.023743034206188739, 0.020678772648531595, 
    0.01797964139781856, 0.015594308175210984, 0.013480938996750697, 
    0.01160560343314756, 0.0099408870466127664, 0.0084647270555270725, 
    0.0071594205349556897, 0.0060107929965863673, 0.0050074397643898117, 
    0.0041400498350081067, 0.0034007685456612959, 0.0027826036745564296, 
    0.0022788960216579834, 0.0018828672077929323, 0.0015872679268456339, 
    0.0013841531503606462, 0.0012647750593775002, 0.0012196272187868834, 
    0.0012385844600828338, 0.0013111433220060081, 0.0014267214395968716, 
    0.0015749636788465887, 0.0017460449259444838, 0.0019309270427938664, 
    0.0021215601265441725, 0.0023110307353478906, 0.0024936457553760578, 
    0.0026649645040939919, 0.0028217704201931172, 0.0029619991270223474, 
    0.0030846207245216737, 0.0031894802640119978, 0.0032771104627251288, 
    0.0033485141606070445, 0.0034049427232506701, 0.0034476671784460879, 
    0.0034777817069364531, 0.0034960210510920318, 0.0035026383115448309, 
    0.0034973189659514487, 0.0034791773589140985, 0.0034468217128864557, 
    0.003398487730920152, 0.0033322412365086873, 0.0032462147153231049, 
    0.003138843828239733, 0.0030091006865111277, 0.0028566531126653222, 
    0.0026819707907460642, 0.0024863348884944592, 0.0022717649554641968, 
    0.0020408557560919324, 0.0017965583761603058, 0.0015419135046526654, 
    0.0012797859590798029, 0.0010126179095196353, 0.00074224539369581542, 
    0.00046980816954721242, 0.00019576254852627365, -8.0000378616568754e-05, 
    -0.00035794022750972043, -0.000638593234088478, -0.00092228007968606464, 
    -0.0012088349093187058, -0.0014974098818328454, -0.0017863550987714551, 
    -0.0020732193741297253, -0.0023548578575115853, -0.0026276359905061885, 
    -0.0028877150878600898, -0.0031313797426417525, -0.0033553751987338469, 
    -0.0035572124496568232, -0.003735405102696346, -0.0038896041382344283, 
    -0.0040206208750143586, -0.0041303331463452336, -0.0042214917161321197, 
    -0.0042974477862450979, -0.0043618288261855452, -0.0044182106661842567, 
    -0.0044698202853785552, -0.0045192949102522964, -0.0045685153748505928, 
    -0.0046185029982174879, -0.0046693745883932053, -0.004720348241199007, 
    -0.0047697823966956297, -0.0048152473838926364, -0.0048536218646637128, 
    -0.0048812070974687469, -0.0048938610203825414, -0.0048871479202114961, 
    -0.0048565135494524833, -0.0047974869097545982, -0.0047059193762221934, 
    -0.004578241696861377, -0.0044117232856818152, -0.004204717398968787, 
    -0.0039568511067019285, -0.0036691500834444076, -0.0033440695441015241, 
    -0.0029854284549500716, -0.0025982610140986772, -0.0021885751642785503, 
    -0.0017630480825229933, -0.001328699577926277, -0.00089254327716380784, 
    -0.00046126849683035922, -4.0972493785711647e-05, 0.00036304116590760101, 
    0.0007463931894419074, 0.0011056756381423666, 0.0014384300185141361, 
    0.0017430673748800988, 0.0020187606262452545, 0.0022653122596095541, 
    0.0024830216775437934, 0.0026725746047619845, 0.0028349632613500625, 
    0.0029714196919129396, 0.0030833776574208855, 0.003172440163430467, 
    0.0032403336715571282, 0.003288860608390965, 0.00331983944428452, 
    0.0033350193624632398, 0.0033359951499883234, 0.0033240983075974954, 
    0.0033003142175047537, 0.0032652113675421695, 0.0032189191342337454, 
    0.0031611451167202543, 0.0030912434592188631, 0.0030083266317586484, 
    0.0029114209668279784, 0.0027996355013683179, 0.0026723738685334964, 
    0.0025295483527604636, 0.0023717843999976822, 0.002200564943105672, 
    0.0020182885916580277, 0.0018282112996622704, 0.0016342859650468617, 
    0.0014409142694970936, 0.0012526579750178929, 0.0010739484299178907, 
    0.00090882509693789037, 0.00076071901895409565, 0.00063229237738105426, 
    0.00052532857685417991, 0.00044066062746368523, 0.00037814600770026544, 
    0.00033667832039073887, 0.0003142306088585766, 0.00030792344752003691, 
    0.00031413350767719024, 0.00032863300333771942, 0.00034677669736114222, 
    0.00036372133523667377, 0.00037469573457063769, 0.0003752998130829476, 
    0.00036182182752504764, 0.00033153495286913768, 0.00028293234506793257, 
    0.00021586679356959675, 0.00013157253187948928, 3.2551456679917319e-05, 
    -7.7647922521162838e-05, -0.00019473944457824822, 
    -0.00031405748163752258, -0.0004309196404678948, -0.00054097398793434765, 
    -0.00064049021158869195, -0.00072657799584963589, 
    -0.00079733187337388534, -0.00085188576777470919, 
    -0.00089039800392937346, -0.00091397139091362338, 
    -0.00092451137455009541, -0.00092454353966274017, 
    -0.00091700106449154684, -0.00090499669209214133, 
    -0.00089159585415103768, -0.00087958011865709894, 
    -0.00087122837677883365, -0.0008681195774597393, -0.0008709874839460262, 
    -0.00087963761132697164, -0.00089295872388080394, 
    -0.00090901820810849435, -0.00092525588822066937, 
    -0.00093874197472273752, -0.00094648332626158884, 
    -0.00094573128758766787, -0.00093426109158012394, 
    -0.00091058668372344766, -0.00087409167661931203, 
    -0.00082505210533812955, -0.0007645725270974753, -0.00069443073832993647, 
    -0.00061686441054541327, -0.00053433608948656784, 
    -0.00044929979295407963, -0.00036399862397105558, 
    -0.00028031389120458005, -0.00019966528349313112, 
    -0.00012295359866793231, -5.0555679102774753e-05, 1.7671380966387832e-05, 
    8.2352255566757617e-05, 0.0001445528325838732, 0.00020572887293751648, 
    0.00026767050217407849, 0.00033243921536915802, 0.00040229462198065186, 
    0.00047960693379914656, 0.00056675626639584393, 0.00066602551849050898, 
    0.00077947510564581053, 0.00090881799380045786, 0.0010552948940264594, 
    0.0012195459136466762, 0.0014014971139072574, 0.0016002605998006582, 
    0.0018140730733795843, 0.002040275115127829, 0.0022753576940390268, 
    0.0025150638438570573, 0.0027545689047222097, 0.0029886935514807224, 
    0.0032121575811417009, 0.0034198369110800919, 0.003607015784414943, 
    0.0037696073583974861, 0.0039043430150531352, 0.0040089060432265513, 
    0.0040820205156580835, 0.0041234863781732288, 0.0041341683877605525, 
    0.0041159384321615682, 0.0040715888063897736, 0.0040047017558967083, 
    0.0039195028688840073, 0.0038206833122153105, 0.00371320347499154, 
    0.0036020724268753094, 0.0034921187180431369, 0.0033877570091016959, 
    0.003292765169192908, 0.0032100761225888532, 0.0031415939179251459, 
    0.0030880458714871448, 0.003048865668340426, 0.0030221260606298518, 
    0.0030045194178341538, 0.0029914105977617757, 0.0029769690417539244, 
    0.0029544056385184163, 0.0029163060852057361, 0.0028550589814088307, 
    0.0027633553336272494, 0.002634719405928194, 0.0024640219438301458, 
    0.0022479281549420134, 0.0019852242091090381, 0.0016770110374068584, 
    0.0013267399273775224, 0.00094008686774386333, 0.00052470073544729032, 
    8.983179540423907e-05, -0.0003541027137898597, -0.00079598894134672677, 
    -0.0012245042001867092, -0.0016286047458775417, -0.001997997673654489, 
    -0.0023235596597581355, -0.0025976600714966323, -0.0028143690495935868, 
    -0.0029695500959365365, -0.0030608585158021099, -0.0030876916203973542, 
    -0.0030511099285034952, -0.0029537555454308079, -0.0027997633120852919, 
    -0.0025946566503987608, -0.002345221449102315, -0.0020593390607285995, 
    -0.0017457883893069747, -0.0014140078008001477, -0.0010738272372865041, 
    -0.00073516509524728497, -0.00040771452001564658, 
    -0.00010061580884351162, 0.00017787726096783903, 0.00042070054033499, 
    0.00062226719623779719, 0.00077868261140370256, 0.00088790774275023323, 
    0.00094982539137632507, 0.00096621979239515778, 0.00094065878585948841, 
    0.00087828794352000947, 0.00078553666479930901, 0.00066975869151544853, 
    0.00053881461464512612, 0.0004006290343521973, 0.00026275776043161695, 
    0.00013198666443628288, 1.4000674713401972e-05, -8.6837516642266358e-05, 
    -0.00016761360144556514, -0.00022686915127095265, 
    -0.00026451158212813448, -0.00028166292772387446, 
    -0.00028044819854471494, -0.00026376458036955422, 
    -0.00023505609036503163, -0.00019807959222759746, 
    -0.00015669167282636792, -0.0001146356282948167, -7.5338941138753047e-05, 
    -4.1718013500989575e-05, -1.6029990887159276e-05, 2.4497592244972525e-07, 
    6.4564087328780357e-06, 2.8000592612258639e-06, -9.7282366899108745e-06, 
    -2.9405752637433002e-05, -5.3911747304961151e-05, -8.048789838998948e-05, 
    -0.00010615386410843407, -0.00012795111119545455, 
    -0.00014321133489690764, -0.00014982210159821923, 
    -0.00014646834625411665, -0.00013281637587595846, -0.0001096215324895078, 
    -7.8743738367891055e-05, -4.3074249299300971e-05, 
    -6.3741850277004538e-06, 2.6966880329768134e-05, 5.2232805086643928e-05, 
    6.471728237506365e-05, 6.0064735167836872e-05, 3.4591707708806537e-05, 
    -1.4454294845480612e-05, -8.8714456624881181e-05, 
    -0.00018862914333050252, -0.00031342640656002285, 
    -0.00046120110585129182, -0.00062904031736745088, 
    -0.00081318220084155841, -0.0010091898197748641, -0.0012121210755342521, 
    -0.0014166965154076465, -0.0016174631544118613, -0.0018089506503007372, 
    -0.001985817947830819, -0.0021429792695214158, -0.0022757036512726383, 
    -0.0023797065697564929, -0.0024512359610164049, -0.0024871678422009485, 
    -0.002485104966631852, -0.0024435026101185921, -0.0023617932105146787, 
    -0.0022405118614178344, -0.0020813937497443126, -0.0018874324984653359, 
    -0.0016628615005139366, -0.0014130752182376859, -0.0011444431896700377, 
    -0.00086403817217173544, -0.00057928979463117865, -0.000297593843871862, 
    -2.5915989792811458e-05, 0.00022957133797149067, 0.00046377945590684347, 
    0.00067288684906142418, 0.00085441604045068164, 0.0010071904855014618, 
    0.0011312012343268479, 0.0012273857899007981, 0.0012973808030155493, 
    0.0013432569624133677, 0.0013672750854662756, 0.0013716864542988073, 
    0.0013585901321069159, 0.0013298425098974926, 0.0012870268695318599, 
    0.0012314566257694182, 0.001164204715450218, 0.0010861438131907295, 
    0.00099799715662565605, 0.00090039909172123507, 0.00079397960910433608, 
    0.00067945703748324129, 0.00055775868269848693, 0.00043011920114321793, 
    0.0002981680876279403, 0.0001639555091087451, 2.9921740345668912e-05, 
    -0.00010120270946405949, -0.00022654822522708815, 
    -0.00034328933735933652, -0.00044884320217955412, 
    -0.00054103605028997287, -0.00061823119201033071, 
    -0.00067941888283526821, -0.00072424565846945419, 
    -0.00075301559197176815, -0.00076666282104899375, 
    -0.00076670671775771614, -0.00075517930193674419, 
    -0.00073452713771104408, -0.0007074780520855558, -0.0006768851505203823, 
    -0.00064556302184703171, -0.00061611977862619774, 
    -0.00059081011714431073, -0.00057141219622884902, 
    -0.00055912279719969862, -0.00055448880034145718, -0.0005573743808650304, 
    -0.00056695763662063705, -0.00058177473410358409, 
    -0.00059980173236774161, -0.00061858790124407891, 
    -0.00063541759933950889, -0.00064751469104381838, 
    -0.00065226717441020708, -0.00064746543271554705, -0.0006315307896306631, 
    -0.00060370737839844711, -0.00056420040591113711, 
    -0.00051423167833979707, -0.00045599675354834207, -0.00039252622923968, 
    -0.00032745448890952633, -0.0002647350759306784, -0.00020830038186062062, 
    -0.00016171725681892276, -0.00012785382339893577, -0.0001085961183366143, 
    -0.00010465289253256007, -0.00011546723701891509, 
    -0.00013926772686554138, -0.00017325448980477079, 
    -0.00021389347501470291, -0.00025729401871573771, 
    -0.00029962605447444004, -0.00033752707107295661, 
    -0.00036845982071923201, -0.00039097769067120635, 
    -0.00040488324353451046, -0.00041127196958475477, 
    -0.00041246175349746595, -0.000411827348874865, -0.00041356060244116617, 
    -0.0004223757197421609, -0.00044319051156219678, -0.00048079146090891742, 
    -0.00053949780494683315, -0.00062286952332480717, 
    -0.00073344904795153711, -0.00087258220446926802, -0.0010403009945758282, 
    -0.0012352806435268226, -0.0014548469695096194, -0.0016950459346237747, 
    -0.0019507528660097375, -0.002215847722717205, -0.0024834418342422233, 
    -0.002746176444096385, -0.002996566312240241, -0.0032273693509813459, 
    -0.0034319559354046266, -0.0036046256194920182, -0.0037408911632552905, 
    -0.0038376673941566035, -0.0038933960766192686, -0.0039080804721644486, 
    -0.0038832425576576304, -0.0038217911871486539, -0.0037278403538498215, 
    -0.0036064754724284697, -0.0034634914913078321, -0.0033051273991370313, 
    -0.003137808381353053, -0.0029679127056923141, -0.0028015755831259986, 
    -0.0026445295535380618, -0.0025019753258768056, -0.002378472796508616, 
    -0.0022778443687145118, -0.0022030857127475802, -0.0021563099206615534, 
    -0.002138723313523873, -0.0021506407293667646, -0.002191521662053312, 
    -0.0022600201990831559, -0.0023540403951269238, -0.0024707974646836863, 
    -0.0026068881470386212, -0.002758387113111339, -0.0029209569027750623, 
    -0.0030899781927154163, -0.003260699827620164, -0.0034284037796335643, 
    -0.0035885796981617387, -0.0037371119049806611, -0.0038704482040565211, 
    -0.0039857285027872988, -0.0040808580887990789, -0.0041545075198398083, 
    -0.0042060399183784635, -0.0042353787833831627, -0.0042428515120644487, 
    -0.0042290128847936592, -0.0041945050416725615, -0.0041399455295010722, 
    -0.0040658647796216283, -0.0039726913549705334, -0.0038607604469949102, 
    -0.0037303637245277199, -0.0035818162618118025, -0.0034155406710437166, 
    -0.0032321650216081644, -0.0030325894005296897, -0.0028180306763648504, 
    -0.0025900174846551303, -0.0023503656205056539, -0.0021011316871703115, 
    -0.0018445773853705181, -0.0015831583869400459, -0.0013195247789154346, 
    -0.0010565456159902374, -0.00079730651519903666, -0.00054509490901962399, 
    -0.00030334484564657576, -7.553553092505048e-05, 0.00013492598747669941, 
    0.00032483407745950038, 0.00049129660290603782, 0.00063183331396833217, 
    0.0007444401310191664, 0.00082762960653320959, 0.00088044194498433333, 
    0.00090243566943977904, 0.00089367325738876698, 0.00085470317957829663, 
    0.00078656442450505027, 0.00069080769537623737, 0.00056954715037347528, 
    0.00042551083498150222, 0.00026208575895745684, 8.3322880474582877e-05, 
    -0.00010610869427940295, -0.00030103709305805593, 
    -0.00049595375620857909, -0.00068523486709436165, 
    -0.00086338311544156626, -0.0010252733753568753, -0.0011663846953175348, 
    -0.0012830023886285496, -0.0013723661780943388, -0.0014327844399147881, 
    -0.001463688599401816, -0.0014656492787626606, -0.0014403314505990774, 
    -0.001390417653802246, -0.0013194809438223942, -0.001231818605784114, 
    -0.0011322324701698856, -0.0010257668269982967, -0.00091739664471483231, 
    -0.00081168692793532119, -0.00071244496767462252, -0.0006223956359798779, 
    -0.00054290490982687658, -0.00047379769346313639, 
    -0.00041327946146355282, -0.00035798941626843863, 
    -0.00030317842127227767, -0.00024300924058151747, 
    -0.00017095256973835506, -8.0271100345111375e-05, 3.5446272162590383e-05, 
    0.00018173407704742467, 0.00036271469874979965, 0.00058064246566304917, 
    0.0008355484172835291, 0.0011250311694947679, 0.0014441991208017793, 
    0.0017857850147863046, 0.0021404247786977028, 0.0024970850297845151, 
    0.0028436401807695106, 0.0031675311126794403, 0.0034564894349642023, 
    0.0036992566504499601, 0.0038862592534167806, 0.0040101788177758814, 
    0.0040663854551316542, 0.0040531874977541077, 0.00397189998059064, 
    0.0038267127019921787, 0.0036243813319307514, 0.0033737429481718218, 
    0.0030851247349455561, 0.0027696918255702379, 0.002438786956803165, 
    0.0021033344023881025, 0.0017733357099252319, 0.0014575020795184045, 
    0.0011630183623987209, 0.00089544995932762546, 0.0006587602448943151, 
    0.00045544701749982406, 0.00028674062070393151, 0.00015287107354853142, 
    5.334520720243045e-05, -1.2770418867190771e-05, -4.6606998356018252e-05, 
    -4.9318380477272319e-05, -2.1986693610482488e-05, 3.439205102048694e-05, 
    0.00011883345803138655, 0.00023022815233786657, 0.00036716150577227884, 
    0.00052772007434567542, 0.0007093236430477756, 0.0009085864838352469, 
    0.0011212589615284801, 0.0013422493403415382, 0.00156573981368476, 
    0.0017854017468079545, 0.0019946844220221148, 0.0021871694032220283, 
    0.0023569499606929827, 0.002498978282778383, 0.0026093763327421156, 
    0.0026856596714539055, 0.0027268720772239069, 0.0027336130492530792, 
    0.002707972346325067, 0.0026533670452142748, 0.0025743144548008214, 
    0.0024761349872125748, 0.0023646474455850139, 0.0022458300868898992, 
    0.0021255023589884553, 0.0020090265187806479, 0.0019010443943202136, 
    0.0018052705291006727, 0.0017243634364877108, 0.0016598952150270814, 
    0.0016123967733869312, 0.0015814774620909256, 0.0015659732584345756, 
    0.0015641254788684295, 0.0015737520619930354, 0.001592401591334718, 
    0.0016175004694408777, 0.0016464949352531786, 0.0016769779157356887, 
    0.001706799100409532, 0.001734154125903423, 0.0017576175245711885, 
    0.0017761437061727993, 0.0017889995319979772, 0.0017956548754711078, 
    0.0017956592594986478, 0.0017885069540010245, 0.0017735131583868937, 
    0.0017497276723623929, 0.0017158953255997176, 0.0016704859758450684, 
    0.001611771356951325, 0.0015379714972356506, 0.001447447320155177, 
    0.0013389325756726479, 0.0012117835158841641, 0.0010662347674495576, 
    0.00090361391840007859, 0.00072650424375819722, 0.00053880763322531689, 
    0.00034568262951207879, 0.00015334834402227712, -3.126181742229314e-05, 
    -0.00020096579117991975, -0.00034887915577138111, 
    -0.00046897885636836467, -0.00055663943268286029, 
    -0.00060905170520457593, -0.00062547012893687999, 
    -0.00060728404527901441, -0.00055786987545101161, -0.0004822719770707026, 
    -0.000386743671718119, -0.00027821622552393429, -0.000163761574659818, 
    -5.0104927295559491e-05, 5.6754921038861531e-05, 0.00015181153675737849, 
    0.0002312010420251315, 0.00029223274360751748, 0.00033333225493169071, 
    0.00035390598148981754, 0.00035416316811121701, 0.00033490249500784931, 
    0.0002973078071658846, 0.0002427480963272431, 0.00017264934129883314, 
    8.8426216124009595e-05, -8.490627021355134e-06, -0.00011656489969140351, 
    -0.00023402202515230625, -0.00035871168187998911, 
    -0.00048801084853052019, -0.00061877996789250613, 
    -0.00074738522530373871, -0.00086978082291549888, 
    -0.00098160447197267434, -0.001078288864802145, -0.0011552026381954205, 
    -0.0012078134256938583, -0.0012318896322148375, -0.0012237205793100372, 
    -0.0011803431943454876, -0.0010997553410704425, -0.00098108577303182391, 
    -0.00082471248726422486, -0.00063232510429317272, 
    -0.00040691377279261697, -0.000152701836428859, 0.00012498251649184754, 
    0.00041988722974217567, 0.00072506428960515245, 0.0010331404985580936, 
    0.0013366131323766239, 0.0016281458023080834, 0.0019008659803562919, 
    0.0021486292046543945, 0.0023662484757568636, 0.0025496683120738487, 
    0.0026960760585183772, 0.002803950838168548, 0.0028730635128415569, 
    0.0029044204261522133, 0.002900167890801528, 0.0028634420172443664, 
    0.0027981689717718593, 0.0027088215535339332, 0.0026001267272279622, 
    0.0024767600543031624, 0.0023430141980727574, 0.0022025149587190681, 
    0.0020579831518113306, 0.0019110798990607234, 0.0017623603929846059, 
    0.0016113347889829147, 0.0014566220196050692, 0.0012961916152587532, 
    0.0011276593719929632, 0.00094861404120600104, 0.00075694269788004578, 
    0.00055114128652164257, 0.00033055751758637847, 9.5562808801255453e-05, 
    -0.00015237018127211329, -0.00041068375107482756, 
    -0.00067583135626307666, -0.0009434519433296467, -0.0012085851574479762, 
    -0.0014659065572088768, -0.0017099769479823499, -0.001935455353192106, 
    -0.0021372716155977321, -0.0023107800297534837, -0.0024518891237869656, 
    -0.0025571906538432473, -0.0026241038440540823, -0.0026510285767174465, 
    -0.0026375056360134473, -0.0025843649538476788, -0.0024938441884110474, 
    -0.0023696354961155693, -0.0022168417033742267, -0.0020418388397542985, 
    -0.0018520345054265645, -0.001655522388494536, -0.0014606585667720803, 
    -0.0012755941563650627, -0.0011077779281246623, -0.00096349886273051173, 
    -0.00084748498859188697, -0.00076261760146420108, 
    -0.00070976894722257202, -0.00068780335487220092, 
    -0.00069372340632036671, -0.0007229624802552189, -0.00076977334653236017, 
    -0.00082769688053880089, -0.00089004399269084389, 
    -0.00095035578542956704, -0.0010028235165729217, -0.0010426140897867816, 
    -0.0010660847572768694, -0.0010709031251371398, -0.0010560534346205853, 
    -0.00102176337031867, -0.00096938271261426303, -0.00090121511608254096, 
    -0.000820340131131146, -0.00073042953252846121, -0.00063553883990570353, 
    -0.00053989765462718331, -0.00044768080821902463, 
    -0.00036278150187787916, -0.00028858188821517258, 
    -0.00022776657824599448, -0.00018217405882230649, 
    -0.00015271504260665539, -0.00013935378078786773, 
    -0.00014115521987344683, -0.00015639087691512104, 
    -0.00018268048173729736, -0.00021717834517711741, 
    -0.00025676597426937633, -0.00029826531405033785, 
    -0.00033862127526142308, -0.00037508253570554524, 
    -0.00040531619945029511, -0.00042751168014381371, 
    -0.00044042177197691575, -0.00044337425615023282, 
    -0.00043624483050562463, -0.00041939998449793726, 
    -0.00039362550096866492, -0.00036004208483700323, 
    -0.00032000815875043022, -0.00027503377418999254, -0.0002266845844334627, 
    -0.00017648337462831793, -0.00012581706089838127, 
    -7.5843738214291629e-05, -2.7421073233389554e-05, 1.8937306653917996e-05, 
    6.307943090786558e-05, 0.00010519253907107198, 0.00014574273314824367, 
    0.0001853951967821858, 0.00022493270194063253, 0.00026517515292922086, 
    0.00030692357716796117, 0.00035094139467942544, 0.00039796280227677851, 
    0.0004487349605816638, 0.00050405806444822816, 0.00056482236477694366, 
    0.00063200534542636898, 0.00070663239813346566, 0.00078969024731262623, 
    0.00088200985656059958, 0.00098413249770732975, 0.0010961989323377513, 
    0.0012178795317011883, 0.0013483719563552156, 0.0014864599591322147, 
    0.0016306262248057955, 0.0017791673130077761, 0.0019302873062999831, 
    0.0020821189857643304, 0.0022326933267385581, 0.002379860548453446, 
    0.0025212131017952029, 0.0026540256488473738, 0.0027752699973380901, 
    0.0028816962495599461, 0.0029700051071092992, 0.0030370685505057668, 
    0.0030801792154668559, 0.0030972891460619668, 0.0030872201641421442, 
    0.0030498112999381953, 0.0029860133746802951, 0.002897899975828211, 
    0.0027886330171818297, 0.0026623281280543196, 0.0025238579647452442, 
    0.0023785841924858354, 0.0022320104804722791, 0.002089398170873526, 
    0.0019553582961223657, 0.0018334682347595666, 0.0017259638371974093, 
    0.0016335321422900708, 0.0015552603495994411, 0.0014887216116673146, 
    0.0014301943254651204, 0.001374985318877475, 0.0013178164729335407, 
    0.0012532468822384622, 0.0011760934548830414, 0.0010818507458645607, 
    0.00096707035016685449, 0.00082969603788740631, 0.00066931227115771133, 
    0.0004872859998527626, 0.00028678277035632763, 7.2633595085689934e-05, 
    -0.00014892717342404388, -0.00037062724476145947, 
    -0.00058459453836047189, -0.00078279445454399821, 
    -0.00095745834005246254, -0.0011014435287710783, -0.0012085360966458368, 
    -0.0012736707202165673, -0.0012930951315777294, -0.0012644990479678446, 
    -0.0011870932126584028, -0.0010616685272009478, -0.00089059885926802277, 
    -0.00067778577970147654, -0.00042850986374096036, 
    -0.00014919980890918766, 0.0001528774228511857, 0.00046997960483958286, 
    0.00079425127576758601, 0.001118067122831749, 0.0014343190306892351, 
    0.0017366070056012584, 0.0020193627583536262, 0.0022778703243969685, 
    0.0025082409861558203, 0.00270734956628047, 0.0028727447355288327, 
    0.0030025926482772944, 0.0030956391399439057, 0.0031512061705532687, 
    0.00316922966562497, 0.003150296242781504, 0.0030956895866527984, 
    0.0030074007410770078, 0.0028880844178330429, 0.0027409439546681727, 
    0.0025695336603194759, 0.0023774937625854874, 0.0021682693594485113, 
    0.0019448458972121084, 0.001709609976625245, 0.0014643487181279667, 
    0.0012104097740868612, 0.00094898207365934394, 0.00068139909748767338, 
    0.00040937177071856564, 0.0001350739525148556, -0.00013894242962910299, 
    -0.00040998726666208489, -0.00067554772332520331, -0.00093361133602441358, 
    -0.001182921250682097, -0.0014230992536001194, -0.0016546758710128677, 
    -0.0018789841883410526, -0.0020979856729973273, -0.0023140431921505676, 
    -0.0025296473716478192, -0.0027471577244292575, -0.0029685372073827519, 
    -0.0031951205292575996, -0.0034274338055227112, -0.0036650654749197892, 
    -0.0039066161784413076, -0.0041497105225008586, -0.0043910675745347438, 
    -0.0046266452588377268, -0.0048518323698678537, -0.0050617057291477774, 
    -0.0052512966524428774, -0.00541585810430427, -0.0055510899785555581, 
    -0.005653285431201689, -0.0057194380412272927, -0.0057473098486575218, 
    -0.0057354835628277874, -0.0056834187468399666, -0.0055915027188560467, 
    -0.0054610617344033729, -0.0052943312536287077, -0.0050943454082186179, 
    -0.0048647804668645401, -0.0046097340240723586, -0.0043334892941509339, 
    -0.0040402912361275026, -0.00373415291998082, -0.0034187223325397899, 
    -0.0030972256361776964, -0.0027724712619383949, -0.0024469030110162784, 
    -0.0021226631072010036, -0.0018016413250600035, -0.0014855031254928082, 
    -0.0011756869586907034, -0.00087341473455257554, -0.00057972745154120735, 
    -0.00029558344458732803, -2.1992852322199359e-05, 0.00023981524702692392, 
    0.0004882368294443439, 0.00072119262907571096, 0.00093609013782822853, 
    0.0011298786597023912, 0.0012991682626197348, 0.0014403755337773359, 
    0.0015499109962022204, 0.0016243589718662934, 0.0016606669577949914, 
    0.0016563648021782646, 0.0016098212321471895, 0.001520518209956607, 
    0.0013893189460172147, 0.0012186691648672376, 0.0010127106723326256, 
    0.00077727462104516787, 0.00051975858504726394, 0.00024891054541674494, 
    -2.5497491809408387e-05, -0.00029308924582402039, 
    -0.00054338306596329519, -0.00076636861503026729, -0.0009531193230217646, 
    -0.00109637196515031, -0.0011910281374028372, -0.0012345081815998422, 
    -0.0012269152531382604, -0.001170957287739556, -0.0010716636405693196, 
    -0.00093588800218449624, -0.00077167510114239967, 
    -0.00058757430428327522, -0.00039196724471198186, 
    -0.00019250109241179984, 4.3329693927326562e-06, 0.00019343843877862762, 
    0.00037118424269452348, 0.00053530170322370124, 0.00068467278397874693, 
    0.00081903191013905853, 0.00093863352195990815, 0.0010438916607428341, 
    0.001135036550617853, 0.0012118318047546692, 0.0012733564632511881, 
    0.0013179259067652978, 0.0013431614301130735, 0.0013462047211060153, 
    0.0013240689764089833, 0.0012740448885518389, 0.0011941195212720795, 
    0.0010833468918191279, 0.00094214671435754755, 0.00077248316327491, 
    0.00057790681456218072, 0.00036346998318780759, 0.00013550934558284383, 
    -9.8692685949269563e-05, -0.00033131339872221661, 
    -0.00055444117819944318, -0.00076054010031717252, 
    -0.00094287931593882196, -0.0010958908106352085, -0.0012154439635968966, 
    -0.0012990135466127218, -0.0013457521608174765, -0.0013564454695106105, 
    -0.0013333654179378883, -0.001280070204095908, -0.0012011217341449255, 
    -0.0011017700422799254, -0.00098762891102720891, -0.00086437515088485183, 
    -0.00073745199220028035, -0.0006117853089663461, -0.00049153542051686447, 
    -0.00037988374763675461, -0.00027888498775002004, 
    -0.00018940898646622973, -0.00011119651364840358, -4.30141525749953e-05, 
    1.7119167958659198e-05, 7.1690809999412229e-05, 0.00012347051833674238, 
    0.00017532318007901514, 0.00023007197160653946, 0.00029040044822190394, 
    0.00035878708734157696, 0.0004374620536132806, 0.00052836056298902938, 
    0.00063308467175859017, 0.00075285124026752605, 0.00088843193979408226, 
    0.0010400979855587911, 0.0012075558995822354, 0.0013899006824691675, 
    0.0015855591079801999, 0.0017922470904700857, 0.0020069487872484311, 
    0.002225937552605339, 0.0024448630176516564, 0.0026589146510586073, 
    0.0028630503963120043, 0.0030522853376635482, 0.0032219896517389538, 
    0.0033681768104744875, 0.0034877400911657464, 0.0035786216497374519, 
    0.0036399137576767385, 0.0036718898256914204, 0.0036759866461624525, 
    0.0036547223318108045, 0.0036115652106733492, 0.0035507458017820992, 
    0.0034770297176780185, 0.0033954481207577008, 0.0033109839869549947, 
    0.0032282822710220172, 0.003151356746831585, 0.0030833489295693651, 
    0.0030263361920868379, 0.0029812000906832719, 0.0029475822862704672, 
    0.0029239415809020316, 0.0029077201709712388, 0.0028955987260239854, 
    0.0028838074760951867, 0.0028684583770042923, 0.0028458692283764497, 
    0.0028128118004149359, 0.0027666992941348841, 0.0027056658159178965, 
    0.0026285657416244301, 0.0025349174951732286, 0.0024247971171339699, 
    0.0022987470304286842, 0.0021576891950842725, 0.002002874617676194, 
    0.0018358609272790738, 0.0016585099268397086, 0.0014729832814328835, 
    0.0012817191029446187, 0.0010873858488369662, 0.00089281255371394383, 
    0.000700872935030304, 0.00051435597851755732, 0.00033582769296256246, 
    0.00016751262326443353, 1.12075880195282e-05, -0.00013176514944030881, 
    -0.00026058177971363498, -0.00037489626377318656, 
    -0.00047482545559509855, -0.00056092914378529524, -0.0006341798913458216, 
    -0.00069590282548497517, -0.00074769124295298117, 
    -0.00079127769495568865, -0.00082835416916306507, 
    -0.00086036512971299694, -0.00088829824972761449, 
    -0.00091250809048921131, -0.00093260412442340416, 
    -0.00094745325734673237, -0.0009552794897171212, -0.00095387842651740323, 
    -0.00094088348884526168, -0.00091406792630812056, 
    -0.00087159318349944138, -0.00081225337326567453, 
    -0.00073561507822348824, -0.00064210567312194926, 
    -0.00053305166681192858, -0.00041065093101016689, 
    -0.00027789249807987429, -0.00013844032916838069, 3.5274624727709846e-06, 
    0.00014351019274541253, 0.0002768973934168094, 0.00039918165604253141, 
    0.00050614906970402804, 0.00059403713659063524, 0.0006596502553765539, 
    0.00070042353697504032, 0.00071444196521971385, 0.00070043880246930027, 
    0.00065776826941462492, 0.00058638680790496379, 0.00048682698545904834, 
    0.00036020083712251657, 0.00020820109322486097, 3.3126987833895271e-05, 
    -0.00016210347720857163, -0.00037397996602291512, 
    -0.00059848012544297131, -0.00083120936634869776, -0.0010676120294308014, 
    -0.00130321513167724, -0.0015338881278525579, -0.0017560599978849898, 
    -0.0019668858619987517, -0.0021643368237530955, -0.002347233557918852, 
    -0.0025151969399111471, -0.0026685750700093541, -0.002808329271982568, 
    -0.0029358978984669738, -0.0030530215244019623, -0.0031615459371169418, 
    -0.0032632196999035747, -0.0033594905771164489, -0.0034513408850172641, 
    -0.0035391736149635103, -0.0036227159113113054, -0.0037009643409758753, 
    -0.0037721674949385722, -0.0038338511624181962, -0.0038829176207983147, 
    -0.0039158170451991936, -0.0039287849977565582, -0.003918158417583131, 
    -0.003880709819603268, -0.0038139644505092245, -0.0037164712822348712, 
    -0.0035879770824186852, -0.0034295056967192689, -0.0032433177471759039, 
    -0.00303277538416137, -0.002802137520371941, -0.0025563265774458492, 
    -0.0023006847050253813, -0.0020407536618209845, -0.0017820889790891861, 
    -0.0015301045176376404, -0.0012899337910749215, -0.0010662975113223802, 
    -0.00086337180375929288, -0.00068466965755571859, 
    -0.00053292904050210733, -0.00041004512750354076, 
    -0.00031702872148568122, -0.00025402500924400211, 
    -0.00022035812667799072, -0.00021462211819772258, 
    -0.00023477897785180587, -0.0002782559648505697, -0.00034204280664167162, 
    -0.00042276283704790509, -0.00051670381948554754, 
    -0.00061982741740167181, -0.00072776160262382871, 
    -0.00083583873065182657, -0.0009391749970812911, -0.0010328225170310973, 
    -0.0011119701998863018, -0.001172205161290698, -0.0012097912376264727, 
    -0.0012219367052121997, -0.0012070587876526031, -0.0011650038937924523, 
    -0.0010971775459144722, -0.0010065381860016344, -0.00089740381384807862, 
    -0.00077507618917323326, -0.00064533055095015958, 
    -0.00051385050621651569, -0.00038573706590055263, 
    -0.00026518246812080621, -0.00015529510439995603, 
    -5.8112119637316223e-05, 2.5290040598278384e-05, 9.4611378260298334e-05, 
    0.00015013315905699969, 0.00019251148278333726, 0.00022260163510115117, 
    0.00024128925747050444, 0.00024937212354264181, 0.00024746241203683482, 
    0.00023595344177698816, 0.00021504333271953345, 0.0001848279174280533, 
    0.00014546047271616583, 9.736496796419923e-05, 4.1469758487452973e-05, 
    -2.0566845320237195e-05, -8.6225076090865266e-05, 
    -0.00015207691927919214, -0.00021387765372680501, -0.0002667435716241419, 
    -0.0003054057081898733, -0.00032448503013588289, -0.00031876916089279041, 
    -0.00028347082577654916, -0.00021446981111169507, 
    -0.00010853885300491446, 3.6419545283114985e-05, 0.00022114992144334455, 
    0.00044483130867041938, 0.00070490948216029225, 0.000997007521410926, 
    0.0013149894947282852, 0.0016511504982587863, 0.0019965860722126567, 
    0.0023416872446196391, 0.0026767332319964808, 0.0029925046719560221, 
    0.0032808893472856342, 0.0035354017822000678, 0.0037515684060001331, 
    0.0039271535110490322, 0.0040621784897211669, 0.0041587590716664329, 
    0.0042207637494004416, 0.0042533176065266964, 0.0042622508498075303, 
    0.0042535019444255827, 0.0042325686662554162, 0.0042039954896496024, 
    0.0041709787897570754, 0.0041350870503401331, 0.0040960999280724216, 
    0.0040520302119009931, 0.0039993202412934512, 0.0039332231751079832, 
    0.0038483385687572281, 0.0037392568574948484, 0.0036011767870451311, 
    0.0034304709549775581, 0.0032250525243316145, 0.0029845726064111526, 
    0.0027104442401929291, 0.0024057139769836098, 0.0020747830323460436, 
    0.0017230230799855873, 0.001356362625963, 0.00098079596173464073, 
    0.00060195331869410107, 0.00022471677286098172, -0.00014704562341763566, 
    -0.0005106202249598365, -0.00086442843367002414, -0.0012078888548728295, 
    -0.0015411695698687544, -0.0018648977114648509, -0.0021798560717155766, 
    -0.002486730560258795, -0.0027859232610598509, -0.0030774663820831672, 
    -0.0033609915632692635, -0.0036357719032067961, -0.0039007732237473329, 
    -0.0041547022876622626, -0.0043960581199483702, -0.0046231843545598665, 
    -0.004834331736752134, -0.0050277704001403835, -0.0052019286222423433, 
    -0.0053555637629628377, -0.0054879463493640486, -0.0055990513415638214, 
    -0.0056896972846557014, -0.0057616666597866085, -0.0058177646677111099, 
    -0.0058617381407476974, -0.0058981029644115989, -0.005931828355205864, 
    -0.0059679558842339548, -0.0060111853935761574, -0.0060655377201240153, 
    -0.0061341102036257464, -0.0062189250194959397, -0.0063208969722378027, 
    -0.0064398610022114479, -0.0065746239038531979, -0.0067230459015986486, 
    -0.0068821685783477552, -0.0070483698386694486, -0.0072175835341978176, 
    -0.0073855251312037228, -0.0075479416132474553, -0.0077008477770028286, 
    -0.0078406957105591844, -0.0079644722071599526, -0.0080697361331155577, 
    -0.0081545650769016473, -0.0082174703351050021, -0.0082572757638110592, 
    -0.0082729795442577306, -0.0082636325398250023, -0.0082282574462195623, 
    -0.0081658305771509752, -0.0080753363294456051, -0.0079559104690658383, 
    -0.0078070336810676195, -0.0076287506237041267, -0.0074218714479740051, 
    -0.0071881241995869639, -0.0069302451900309725, -0.0066519830721060488, 
    -0.0063580407908750249, -0.0060539439041503553, -0.0057458550548817001, 
    -0.0054403780584930811, -0.005144326134745832, -0.004864473075531851, 
    -0.0046072866975336788, -0.0043786820591923143, -0.0041837524003141167, 
    -0.0040265669629170071, -0.0039099781835053443, -0.0038354769935832148, 
    -0.0038030782159728512, -0.0038113029201324363, -0.003857244119532928, 
    -0.0039367321072620552, -0.0040445967416933779, -0.0041749918007310495, 
    -0.0043217240616588203, -0.0044785413901283211, -0.0046393574674403444, 
    -0.0047983906475720156, -0.0049502535739642268, -0.0050900384044069488, 
    -0.0052133936688654649, -0.0053166554144942774, -0.0053969602603424335, 
    -0.0054523522139723665, -0.005481837421448971, -0.0054854062988120142, 
    -0.0054639963337447537, -0.0054194088580997099, -0.0053541447262419059, 
    -0.0052712159318887789, -0.0051739391089331357, -0.0050657547972270418, 
    -0.0049501035347559808, -0.0048303882872717772, -0.0047100119262530197, 
    -0.0045924456960287187, -0.0044812991965074321, -0.0043803181647343254, 
    -0.0042932946176820544, -0.0042238792661413076, -0.004175356279565166, 
    -0.0041503311018239548, -0.0041504601078244299, -0.0041761789128659417, 
    -0.0042264760941196867, -0.0042987221636855569, -0.0043885911287867892, 
    -0.0044900738873856916, -0.0045955955721530941, -0.0046962669440066968, 
    -0.004782232124901406, -0.0048431034523891249, -0.0048684898459863159, 
    -0.004848546981569825, -0.0047745559468783472, -0.0046394679862044579, 
    -0.0044383666654667364, -0.0041688420357155961, -0.0038312293430633202, 
    -0.0034287085393703764, -0.0029672417893933088, -0.0024553459585717028, 
    -0.0019037177428633345, -0.0013247382076796317, -0.00073191690037882748, 
    -0.00013926407001087419, 0.0004393580712376321, 0.00099089027044553914, 
    0.0015037107407974341, 0.0019682047881885083, 0.0023772289117404938, 
    0.0027264202666118739, 0.0030143253525724807, 0.0032423111913514953, 
    0.0034142907935403384, 0.003536294420709993, 0.00361593276702414, 
    0.0036618133738285149, 0.0036829742696845272, 0.0036883953535990156, 
    0.0036865647212399491, 0.0036851467738569814, 0.0036907175200082206, 
    0.0037085755600794416, 0.0037425907366443628, 0.0037951080620822475, 
    0.0038669021344351451, 0.0039571777621126092, 0.0040635849331881165, 
    0.0041823281771294655, 0.0043083517863830448, 0.0044356515473958358, 
    0.0045576840418429711, 0.0046678908533143125, 0.0047602052336747306, 
    0.0048295513761435665, 0.004872214652267246, 0.0048860118176200524, 
    0.0048702739974952058, 0.004825651789561426, 0.0047537656045578882, 
    0.0046568090094184127, 0.0045371414489830814, 0.004396933807082829, 
    0.0042378933619079146, 0.0040611287984012832, 0.003867120660264014, 
    0.0036559436208681208, 0.0034276073620736259, 0.0031824726073340051, 
    0.0029216526561844664, 0.0026472776679652968, 0.0023625679633809912, 
    0.0020717541235515348, 0.0017797918983066096, 0.0014920347358677801, 
    0.0012138659384655047, 0.00095031490655578515, 0.00070578463450070793, 
    0.0004838150489942697, 0.00028690005596171392, 0.00011638789427845117, 
    -2.7573783856599178e-05, -0.00014600279045725776, 
    -0.00024095841895576488, -0.00031530117274843191, 
    -0.00037240805180305676, -0.00041580693831417816, 
    -0.00044883229829661953, -0.00047432750695262878, 
    -0.00049444267035637056, -0.00051048198555295914, -0.000522875493295095, 
    -0.00053119075425479855, -0.00053423827930378445, 
    -0.00053019381467479939, -0.00051673832400153717, 
    -0.00049121943425986915, -0.0004508269998246245, -0.00039279856737562356, 
    -0.0003146571353729626, -0.00021446444941612442, -9.1035920555720463e-05, 
    5.5867166333496156e-05, 0.00022541613468940783, 0.00041567829152748255, 
    0.00062369994011321722, 0.00084565054272868869, 0.0010770628929232663, 
    0.0013130917314685098, 0.0015487836548547158, 0.0017793258169019146, 
    0.0020002653219302396, 0.002207670875360457, 0.0023982614399223673, 
    0.0025695409755614618, 0.0027198526277125018, 0.0028484269125442514, 
    0.0029554109061578565, 0.0030418352210437255, 0.0031095497084287363, 
    0.0031611021653996678, 0.0031995305921410995, 0.0032280946216236379, 
    0.0032500324188853898, 0.0032683906267835486, 0.0032859164267962232, 
    0.0033050204415954847, 0.0033277623220914262, 0.0033558324949963993, 
    0.0033905026504501795, 0.0034325284866166721, 0.0034820163717498389, 
    0.0035383187066043214, 0.0036000069651042862, 0.0036648960982567538, 
    0.0037301416621866395, 0.0037923919152134645, 0.0038479757034159913, 
    0.0038931138236857473, 0.0039241499302472135, 0.0039377574228063135, 
    0.003931141146280139, 0.0039021783285577752, 0.0038494926584494282, 
    0.0037724316888289515, 0.0036709710554312515, 0.0035455885780388808, 
    0.0033971255592676166, 0.0032267099523734209, 0.0030357483775157296, 
    0.0028259793168083909, 0.0025995861825938186, 0.002359279083599061, 
    0.002108308457614852, 0.0018503354281111173, 0.0015892234101973479, 
    0.0013287743222629858, 0.0010724810209024717, 0.00082331233805143307, 
    0.00058356059652213356, 0.00035472743919914417, 0.00013749500433721338, 
    -6.82202269247248e-05, -0.00026314721251046792, -0.00044854158399337091, 
    -0.0006260485045130928, -0.00079756878702029986, -0.00096512928391005205, 
    -0.0011307075566875477, -0.0012960705391729076, -0.0014625702433005306, 
    -0.0016309688197456052, -0.0018013029573371205, -0.0019727935685775353, 
    -0.0021438400711827096, -0.0023120782857409625, -0.0024745073739787259, 
    -0.0026276417606514056, -0.0027676894551131224, -0.0028906910165807584, 
    -0.0029926710620571512, -0.0030697176813210521, -0.0031180158986910443, 
    -0.0031338700133403358, -0.0031137042790429794, -0.0030540459808462077, 
    -0.0029515791002528804, -0.0028032591318048745, -0.0026065055549632809, 
    -0.0023594689841285677, -0.0020613365877771819, -0.0017126246075456473, 
    -0.001315503054072441, -0.00087402686563460617, -0.0003943276353728678, 
    0.00011533994018277636, 0.00064467111861692757, 0.0011815752210949972, 
    0.0017126635452773863, 0.0022239503589008914, 0.0027017614370644805, 
    0.0031335632442392042, 0.0035086555288067617, 0.003818565120079932, 
    0.0040572314322059651, 0.0042210558349169893, 0.0043090339820760215, 
    0.0043229052752877285, 0.0042672923878780645, 0.0041496309562585251, 
    0.0039798876761709115, 0.0037700238838322456, 0.0035333309738170273, 
    0.0032836680523958702, 0.0030347198985170355, 0.0027993223878872786, 
    0.0025889084557893247, 0.0024130380658945105, 0.0022791053622516653, 
    0.0021921747090959346, 0.002155020077289219, 0.0021682981865393702, 
    0.0022308633090537253, 0.0023402478747716138, 0.0024931152986479286, 
    0.0026856717631493017, 0.0029139353482814968, 0.0031738433203346269, 
    0.0034611380834049616, 0.0037711337010377776, 0.0040984029375009667, 
    0.0044364643064526647, 0.0047775772893095727, 0.0051126646377716032, 
    0.0054313821975988013, 0.0057224109215864736, 0.005973892395621164, 
    0.0061740131118413928, 0.0063116986107617581, 0.0063773860090129654, 
    0.0063637876423116293, 0.0062665189168267538, 0.0060845647624937771, 
    0.0058205041735442846, 0.0054804071871850952, 0.0050735526572844945, 
    0.0046118603392315029, 0.0041093024898820277, 0.0035811465251934932, 
    0.0030432497938157228, 0.0025113778964648047, 0.00200065212707436, 
    0.0015249981382847123, 0.0010967486934045714, 0.00072628272431853633, 
    0.00042175689673859952, 0.00018891705532421746, 3.1002203845701196e-05, 
    -5.1289521825069635e-05, -5.9746060719496766e-05, 1.4358264471430772e-06, 
    0.00012573301581486032, 0.00030442704983310218, 0.00052674718134470546, 
    0.00078012985837500721, 0.0010506718669627663, 0.0013237727291672678, 
    0.001584943889740957, 0.0018207434798310836, 0.0020196760230657708, 
    0.0021729152624955271, 0.0022747950466699392, 0.0023229953596923553, 
    0.0023185169033316535, 0.0022654445819749592, 0.0021705839526287908, 
    0.0020430547275885145, 0.0018937810002560861, 0.0017350055089030902, 
    0.0015796531465265234, 0.0014406966611836053, 0.0013304414743230126, 
    0.0012597938053970545, 0.0012376059286352465, 0.0012701092225587047, 
    0.0013605416496699067, 0.0015090479895901697, 0.0017129056428121289, 
    0.0019671016957093085, 0.0022651450712704658, 0.0026000082327327549, 
    0.0029650907200843555, 0.0033550098327266532, 0.0037661275886132339, 
    0.004196772106744886, 0.004647146305788049, 0.0051189320036516793, 
    0.0056146510548785583, 0.0061368497433252466, 0.0066872100829265153, 
    0.0072656900023595943, 0.0078697595447038901, 0.00849392337102336, 
    0.0091295633661702853, 0.0097651589030928933, 0.010386929880907701, 
    0.010979791510275814, 0.011528511385439814, 0.012018927571747984, 
    0.012439042612535093, 0.012779804529860505, 0.013035649339995386, 
    0.013204645409364536, 0.013288397488664106, 0.013291711958654567, 
    0.013222059395760811, 0.013088870716959454, 0.012902638691408636, 
    0.012673990322926348, 0.012412771480475492, 0.012127256724524088, 
    0.011823626182610947, 0.011505774478977887, 0.011175381948308232, 
    0.010832376891936566, 0.010475404111873338, 0.010102469562233977, 
    0.0097114304780255133, 0.0093003567733152357, 0.0088678160610129973, 
    0.0084130253984625366, 0.0079360675722039888, 0.0074380945868958229, 
    0.0069213583019185794, 0.0063891002645613208, 0.0058451950332860858, 
    0.0052935780073394573, 0.0047377514458539181, 0.0041802299639558871, 
    0.0036223715422926211, 0.0030642630272723461, 0.0025047629108565428, 
    0.0019416013155129971, 0.001371554859452037, 0.00079073013483239472, 
    0.00019488396498884867, -0.00042026071721419818, -0.0010587357879892263, 
    -0.0017240697372081226, -0.0024189646199956455, -0.0031447866129093922, 
    -0.003900832348583105, -0.0046834965867360301, -0.0054854846141298135, 
    -0.0062953716642015246, -0.0070977356793376425, -0.0078738892840555536, 
    -0.0086031095207950645, -0.0092642201779852551, -0.0098372445791098176, 
    -0.010304935279430116, -0.010654008978755391, -0.010876002882426164, 
    -0.010967747166229017, -0.010931351891350425, -0.010773849812889303, 
    -0.010506500214457587, -0.010143916956424217, -0.0097030638669826693, 
    -0.0092023256425507217, -0.0086606635516770329, -0.0080970376380044892, 
    -0.007529847687400633, -0.0069765420049331681, -0.0064531355096828251, 
    -0.0059738553735878865, -0.0055507750425720145, -0.0051934358000840126, 
    -0.0049086410350004262, -0.0047004304382896687, -0.0045701359446498595, 
    -0.0045166482372945944, -0.004536753299082907, -0.0046255095121556155, 
    -0.0047765535964945441, -0.0049824419613099793, -0.0052348861522239411, 
    -0.005524801127285932, -0.0058422151354888185, -0.0061760385635050092, 
    -0.0065138059234122522, -0.0068415019201828308, -0.0071437039433699442, 
    -0.0074042957539030086, -0.007607577377712435, -0.0077395612873732032, 
    -0.007789287019249698, -0.0077497217252764858, -0.0076182730144671029, 
    -0.0073968180119960035, -0.007091371515016702, -0.0067115019440934674, 
    -0.0062694794408246655, -0.0057793108273978128, -0.0052558217341723947, 
    -0.0047138230492393624, -0.0041674918397343677, -0.0036299964409114813, 
    -0.0031132966211654721, -0.00262801485035981, -0.002183375084545869, 
    -0.0017868374300897057, -0.001443678068497882, -0.0011562439740905725, 
    -0.00092325756854491018, -0.00073947750250970246, 
    -0.00059568928032369909, -0.00047949029277782261, 
    -0.00037667242586724651, -0.00027307018589303999, 
    -0.00015636599624273547, -1.7714564874244548e-05, 0.00014749257297048496, 
    0.00033950824751429463, 0.00055490040542025573, 0.00078774639954411999, 
    0.0010310860655060559, 0.0012782093155996367, 0.0015236402989087221, 
    0.0017633312763510245, 0.0019944550706584244, 0.0022143667085421474, 
    0.002419594749240154, 0.0026047040616467847, 0.0027616195662729637, 
    0.0028796800882109554, 0.0029464313276311568, 0.0029490883820923724, 
    0.0028762918047605134, 0.0027196815473860408, 0.002474870944404817, 
    0.002141653032297092, 0.0017234033865945408, 0.0012262744093143214, 
    0.00065806847262147358, 2.7418332306027151e-05, -0.00065671152432305072, 
    -0.0013852886315718696, -0.0021490659479118423, -0.0029383026266095675, 
    -0.0037424890863445195, -0.0045504561374621385, -0.0053508528987073123, 
    -0.0061331350410004605, -0.0068887372679729535, -0.0076123267120562022, 
    -0.0083027059894288172, -0.0089632525276187591, -0.0096016722447461941, 
    -0.010229369403380564, -0.010860213258638908, -0.011509243711324446, 
    -0.012191167114187672, -0.012919051575468158, -0.013703071656669622, 
    -0.014549754196711848, -0.015461235213174015, -0.016434708724574969, 
    -0.017462085931310378, -0.018529973055600328, -0.019620133575763157, 
    -0.020710190957691388, -0.021774777290205882, -0.022786633157269982, 
    -0.023717800922581227, -0.024540558894075616, -0.025227994401153427, 
    -0.025754200791176549, -0.026094487431220472, -0.026225768563274108, 
    -0.026127791832603667, -0.025784771273327789, -0.02518783242610451, 
    -0.02433745060186316, -0.023245572886004342, -0.021936451273802716, 
    -0.020446951666322689, -0.018825297634565672, -0.017129302560849647, 
    -0.015423542384670655, -0.01377549283908458, -0.012250380203544834, 
    -0.010906286231526551, -0.0097895503595090434, -0.008931457718110658, 
    -0.0083462282716855081, -0.008030858862588237, -0.0079665234819898591, 
    -0.0081202369625449581, -0.0084479680906448355, -0.0088985411459949707, 
    -0.0094178611924283766, -0.0099525384010576024, -0.010453640208455201, 
    -0.010877504999019653, -0.011187208444000053, -0.011351552154457909, 
    -0.011344410932258023,
  // Fqt-F(7, 0-1999)
    1, 0.99295674792830069, 0.97217746049057585, 0.93868230264000085, 
    0.89406592021873577, 0.84035329391669511, 0.77982782837543096, 
    0.71485407234363518, 0.64771547992622369, 0.58048257680575099, 
    0.51492028332680273, 0.45243644705376118, 0.39406816046054677, 
    0.34049864522638523, 0.29209582753350427, 0.24896360726407388, 
    0.21099795972539792, 0.17794190936649945, 0.1494352594497817, 
    0.12505683171713475, 0.10435844562471509, 0.086890795899675327, 
    0.072222066706850954, 0.059950402310401843, 0.049711392985467749, 
    0.041181713862058579, 0.034079787735644365, 0.028164329572388683, 
    0.023231407467657325, 0.019110594789040335, 0.015660717588594275, 
    0.012765541819952467, 0.010329702404210307, 0.0082750464637639902, 
    0.0065375033778991339, 0.005064492885972955, 0.0038128486631979095, 
    0.0027472002261154506, 0.0018387252266561102, 0.0010642047247407486, 
    0.0004052904408019242, -0.00015209951226282298, -0.00061835183579257171, 
    -0.0010007417351794625, -0.0013041280589709977, -0.0015317355141106876, 
    -0.0016860044573508105, -0.0017694068601447472, -0.0017851428649538277, 
    -0.0017376158670968759, -0.0016326864954584715, -0.0014776580250184849, 
    -0.0012810811401934733, -0.0010523952081055363, -0.00080152798526057301, 
    -0.00053847456306942241, -0.0002729464806133688, -1.4097196097009857e-05, 
    0.00022969992840041995, 0.00045100072238708723, 0.00064341552927617588, 
    0.00080173167184642265, 0.00092201949528327787, 0.0010017367723739229, 
    0.0010398139617106936, 0.0010367028978315062, 0.00099437898659371425, 
    0.00091626956252835597, 0.00080709758495222457, 0.00067262314509222623, 
    0.00051929187392768853, 0.0003538030185741667, 0.00018264276497419657, 
    1.1617553310852547e-05, -0.0001545592889799537, -0.00031255250504805688, 
    -0.00046052001872860337, -0.00059805362444581708, 
    -0.00072594875035301043, -0.00084586721058678449, 
    -0.00095995382987617921, -0.0010704608066152586, -0.0011794048696972996, 
    -0.0012882973204471474, -0.0013979248693852082, -0.0015082203302000136, 
    -0.0016182021238670635, -0.0017260172475774226, -0.0018290626489077121, 
    -0.0019242054162886032, -0.002008056382626858, -0.0020773033049035165, 
    -0.002129042090857524, -0.0021610823104398062, -0.0021721838506760004, 
    -0.0021622167069432984, -0.0021322158735286281, -0.0020843435594048183, 
    -0.0020217596042755941, -0.001948425903792067, -0.0018688579663480344, 
    -0.0017878161885986213, -0.0017099810643168337, -0.0016396221768471848, 
    -0.0015802884466703214, -0.0015345515297411189, -0.0015038332675579571, 
    -0.0014883289128948133, -0.0014870429787023297, -0.0014979337475299228, 
    -0.0015181382252325419, -0.0015442725471947654, -0.0015727527018003975, 
    -0.0016001192112297135, -0.0016233137901578609, -0.0016398726314142036, 
    -0.001648029988906184, -0.0016467253929673149, -0.0016355218012061401, 
    -0.0016144633135459893, -0.001583902246562615, -0.0015443205281298932, 
    -0.0014962079922968582, -0.0014399945449212618, -0.0013760562511958665, 
    -0.0013047823629376675, -0.0012266562135488984, -0.0011423297440245387, 
    -0.001052650176504775, -0.00095863036145612493, -0.00086135630718147738, 
    -0.00076186166397573677, -0.00066098574802366319, 
    -0.00055925612261672336, -0.00045681560105772297, 
    -0.00035341506209109707, -0.00024847392954504009, 
    -0.00014120306739355152, -3.0768735453089651e-05, 8.352725831018413e-05, 
    0.00020206971515431346, 0.00032480306488915527, 0.0004511516981481349, 
    0.00058002805538231192, 0.0007099129104223478, 0.00083901309094168213, 
    0.00096544046724872097, 0.0010874052657292839, 0.0012033527889310145, 
    0.0013120291106415115, 0.0014124612401125696, 0.0015038614687723972, 
    0.0015855029396525627, 0.0016566175715936188, 0.001716387682813467, 
    0.0017640589080757741, 0.0017991790771030823, 0.0018219143064177698, 
    0.0018333537322960786, 0.0018357187871697993, 0.0018323950953366801, 
    0.0018277631052844626, 0.0018268433292962666, 0.0018348050624099491, 
    0.0018564126907870272, 0.0018954991557120719, 0.0019545163829762214, 
    0.0020342463998699119, 0.002133651247897367, 0.00224988696919099, 
    0.002378423081903047, 0.0025132556485577048, 0.0026471840496597983, 
    0.0027721664310514571, 0.0028797693187751546, 0.0029616653731809263, 
    0.0030101446428659347, 0.0030185644944478456, 0.0029817216437241422, 
    0.0028961268262029179, 0.0027602172220624792, 0.0025745183301524436, 
    0.0023417682612306254, 0.0020669756629202959, 0.0017573562101939281, 
    0.0014220985323057423, 0.0010719224661377359, 0.0007184669512912674, 
    0.00037353258989360785, 4.8296886373533734e-05, -0.00024743115348378086, 
    -0.00050580738364480304, -0.00072135528885693243, 
    -0.00089111412257405489, -0.0010145445152384414, -0.0010932079268782206, 
    -0.0011302833268873025, -0.0011299983295804052, -0.0010970468620638721, 
    -0.0010360835284562164, -0.0009513599718807518, -0.00084653850890514348, 
    -0.00072469035147761421, -0.00058845813684811046, 
    -0.00044031531319553509, -0.00028285901112251914, 
    -0.00011906090754475369, 4.7584480635131775e-05, 0.00021304270184979127, 
    0.00037285198854015197, 0.00052235208085561779, 0.00065698371536211696, 
    0.0007726195317407724, 0.00086586885738627222, 0.00093429969767765955, 
    0.00097657409173032106, 0.0009924678782085878, 0.00098279401588405486, 
    0.00094925827509300688, 0.00089427786553812844, 0.00082080954726148703, 
    0.000732218953261186, 0.00063220463340995137, 0.00052476490787766274, 
    0.00041420359660657624, 0.00030512612290251365, 0.00020241265777389228, 
    0.00011111839799312343, 3.6311359402084833e-05, -1.7171492160847411e-05, 
    -4.5020377120293922e-05, -4.3785309856539368e-05, 
    -1.1197023247750413e-05, 5.3556574517838211e-05, 0.00014965492041552856, 
    0.00027459294552704603, 0.0004242767686567484, 0.00059326527124639844, 
    0.00077513523801023862, 0.00096294604279795507, 0.0011497493679594676, 
    0.0013290942300526402, 0.0014954778504191939, 0.0016446913170724592, 
    0.0017740218954002268, 0.0018823062550993542, 0.0019698317905267305, 
    0.002038105995325082, 0.0020895366877978988, 0.0021270540060210324, 
    0.0021537384842693626, 0.0021724816757187505, 0.0021857029135535794, 
    0.002195158363764103, 0.0022018408483224336, 0.00220596812986836, 
    0.002207076114889437, 0.0022041866616711232, 0.0021960381345580973, 
    0.0021813546466677987, 0.0021591197077779701, 0.0021288097815924645, 
    0.0020905662188367242, 0.0020452642382612759, 0.0019944688829912757, 
    0.0019402864338146702, 0.0018851322434174944, 0.0018314369025010896, 
    0.0017813664249595508, 0.0017365743584081175, 0.0016980465134171282, 
    0.0016660772098525194, 0.001640348247635216, 0.0016201189530537857, 
    0.001604461739399934, 0.0015925129396613404, 0.0015836634214310545, 
    0.0015776679554827015, 0.0015746527395548787, 0.001575006014492243, 
    0.0015791795510027517, 0.0015874469094576619, 0.0015996560199167292, 
    0.0016150419713779379, 0.0016321212002675632, 0.0016487030239496683, 
    0.001662010478324386, 0.0016688670642722361, 0.0016659369859195357, 
    0.0016499402170705958, 0.0016178186792177582, 0.0015668252487539532, 
    0.0014945466637542918, 0.0013988848519897012, 0.001278047538394755, 
    0.0011305775182427369, 0.00095545753576889631, 0.00075228819413710748, 
    0.00052150466394513813, 0.00026458771681505202, -1.5787063622992735e-05, 
    -0.00031574258425119239, -0.0006303432288002691, -0.00095392165522984037, 
    -0.0012805610339970688, -0.0016046425845634735, -0.0019213733399300597, 
    -0.0022271732762693328, -0.0025198136066514223, -0.002798278077561233, 
    -0.0030623954322226044, -0.0033123413388024894, -0.0035481512400183301, 
    -0.0037693503098342536, -0.0039747635298757814, -0.0041625142219505898, 
    -0.0043302007027143435, -0.0044751980304788049, -0.0045950296290371302, 
    -0.0046877504237849681, -0.0047522773464631751, -0.0047886167570895116, 
    -0.0047979566766860448, -0.004782629129442174, -0.0047459269365714993, 
    -0.004691834931193517, -0.0046246719642854747, -0.0045487040585912471, 
    -0.0044677790287682585, -0.0043850094718449438, -0.004302553857222273, 
    -0.0042215380987788509, -0.0041421022131713225, -0.0040635860455290112, 
    -0.0039848038529193925, -0.0039043581238420717, -0.0038209559723733086, 
    -0.0037336625461663452, -0.00364206782587912, -0.0035463621092568336, 
    -0.0034473104526377722, -0.0033461575762840094, -0.0032444801419231387, 
    -0.0031440036514721152, -0.0030464238030019869, -0.0029532310465821901, 
    -0.0028655573104254396, -0.0027840624861425979, -0.0027088673448442476, 
    -0.0026395524227657398, -0.0025752163859053077, -0.0025145958324690192, 
    -0.0024562428232999573, -0.0023987109707952299, -0.0023407169797538931, 
    -0.0022812526951808583, -0.002219623843925309, -0.0021553994255105896, 
    -0.0020882742224101257, -0.0020178785212898488, -0.0019435451632280748, 
    -0.0018641289578050649, -0.0017778973121089494, -0.0016825575169423892, 
    -0.0015754116979798494, -0.001453648022799209, -0.0013146820032296398, 
    -0.0011565370345182576, -0.00097817304339339189, -0.00077974237927625769, 
    -0.00056272175363334374, -0.00032994574873564689, 
    -8.5523524249647519e-05, 0.0001653312838550804, 0.00041652191549652033, 
    0.00066134379631198207, 0.00089277073514815522, 0.001103753089727525, 
    0.0012874963245314282, 0.001437711426538263, 0.0015488225304361406, 
    0.0016161441937793701, 0.0016360353680886816, 0.0016060402572737836, 
    0.0015250230690262135, 0.0013932691996788107, 0.001212528260394471, 
    0.00098598134765161142, 0.00071812501442878609, 0.00041457059288587251, 
    8.1801301071615499e-05, -0.0002731455633758228, -0.00064302565609847641, 
    -0.0010207780434606504, -0.0013998890574325371, -0.0017746764825087116, 
    -0.0021404559968157917, -0.0024935899211935382, -0.002831443747324486, 
    -0.0031522637850537666, -0.0034550036049154765, -0.0037391237216820913, 
    -0.0040043767370282314, -0.0042506013643162036, -0.0044775438603286734, 
    -0.0046847230415189688, -0.0048713569244003795, -0.0050363453501584832, 
    -0.0051783003608485631, -0.0052956216638942889, -0.005386588087923477, 
    -0.0054494805559252056, -0.0054827238203855834, -0.0054850646724767674, 
    -0.0054557678970133094, -0.0053948297607687139, -0.0053031480389324516, 
    -0.0051826264032092811, -0.0050361660269010603, -0.0048675549975313714, 
    -0.004681221602440477, -0.0044819120446024938, -0.0042742960482835234, 
    -0.0040625649027464829, -0.0038500726880275437, -0.0036390765222158289, 
    -0.00343061841881324, -0.003224571922247078, -0.0030198409013145432, 
    -0.0028146977602181, -0.0026072019778641282, -0.0023956368932164722, 
    -0.00217889473307785, -0.0019567407851192576, -0.0017299061084183969, 
    -0.001500028556804664, -0.0012694383204289131, -0.0010409076033233745, 
    -0.00081739403061983885, -0.0006018712079550292, -0.00039724400300991333, 
    -0.0002063341765707756, -3.1873533773838983e-05, 0.00012353816803006967, 
    0.00025756725862930861, 0.00036834965694880337, 0.00045471310439381156, 
    0.00051632758752619438, 0.00055372539704723464, 0.00056817932967471551, 
    0.00056148253634163774, 0.00053571819451373164, 0.00049307170614716189, 
    0.00043570453356761986, 0.00036570209105704529, 0.00028508565578250499, 
    0.00019586276382140612, 0.00010010335367162778, 1.6075625608946102e-08, 
    -0.00010200139775101317, -0.00020337721185482034, 
    -0.00030142079673102723, -0.00039344066880558519, 
    -0.00047690708335921807, -0.00054963736111998424, 
    -0.00060996705770949701, -0.00065690160952794124, 
    -0.00069020556553913196, -0.00071043690062304429, -0.000718912170582849, 
    -0.00071761343319410122, -0.00070905733205728805, -0.0006961280457246817, 
    -0.00068189271214929171, -0.00066939401637354263, 
    -0.00066143829228294663, -0.00066039205358625836, 
    -0.00066800036773496756, -0.00068526630478389779, 
    -0.00071239267367800916, -0.0007488074261631989, -0.00079326894077396261, 
    -0.00084402642468637992, -0.00089902010802423164, 
    -0.00095607545853919492, -0.0010130530296332835, -0.0010679388376678219, 
    -0.0011188585149760513, -0.00116403063421179, -0.0012016910601508582, 
    -0.0012300266934836797, -0.0012471402884788158, -0.0012510914648559282, 
    -0.0012400043102184627, -0.0012122316732471746, -0.0011665266370611653, 
    -0.0011021837880570116, -0.0010190922148743521, -0.00091768876558471308, 
    -0.00079879628004900206, -0.00066341669816883352, 
    -0.00051251559168774194, -0.00034688457247382517, 
    -0.00016709461244851823, 2.6418439053743289e-05, 0.00023319538230117624, 
    0.00045254282597114511, 0.00068334265212848942, 0.00092389724001650875, 
    0.0011718353399242749, 0.0014241036148369163, 0.0016770400281258609, 
    0.0019265461588027137, 0.0021683288013262464, 0.0023981779463972588, 
    0.0026122138292817097, 0.0028070798221786052, 0.0029800270394558098, 
    0.0031289129349786199, 0.0032521163288903266, 0.0033484359659367016, 
    0.0034169933403621166, 0.0034571937468007136, 0.0034687493543994596, 
    0.0034517559411721124, 0.0034068131656675004, 0.0033351612870810301, 
    0.0032388214100764704, 0.0031207193321238979, 0.0029847650161438526, 
    0.0028358699423357103, 0.0026798634813188144, 0.0025233076997055004, 
    0.0023732134846245552, 0.0022367140685567535, 0.0021207315380098271, 
    0.002031685701134205, 0.001975271358604739, 0.001956295154447482, 
    0.0019785543679346628, 0.0020447476911246024, 0.0021563885071869187, 
    0.0023137210185347826, 0.0025156042504575183, 0.0027593747592034429, 
    0.003040698121752223, 0.0033534411175086425, 0.0036896122112630601, 
    0.0040394313265949564, 0.0043915536673772848, 0.0047334739035166627, 
    0.0050520737659614625, 0.005334277062354436, 0.005567758100670896, 
    0.0057416165718717693, 0.005846998529336042, 0.0058775740484816328, 
    0.0058298669252033145, 0.0057034269148017883, 0.0055008431798462395, 
    0.0052276274696362382, 0.0048919602023854937, 0.004504307177612423, 
    0.0040769231886997751, 0.0036232534360948242, 0.0031572817830759626, 
    0.0026928529486918156, 0.002243012168931489, 0.0018193876288500814, 
    0.0014316473108312081, 0.0010870349772970701, 0.00079004085945075394, 
    0.00054222588146711492, 0.00034222839566263002, 0.00018597274306534283, 
    6.7061551490082592e-05, -2.2675930981777722e-05, -9.2553498806077761e-05, 
    -0.00015235127381103012, -0.00021167180161794263, 
    -0.00027937069918474187, -0.0003630841356437952, -0.00046885610846873478, 
    -0.00060087278480159048, -0.00076128606754197637, 
    -0.00095014058969739316, -0.0011653844294236982, -0.0014029751555846102, 
    -0.0016570766540855977, -0.0019203292724022864, -0.0021842214548807946, 
    -0.0024395116795374898, -0.0026766931805427964, -0.0028864821890347788, 
    -0.0030602803144625388, -0.0031905888388400272, -0.0032713240767522013, 
    -0.0032980407522703969, -0.0032680216614374212, -0.003180275114482713, 
    -0.0030354372478884261, -0.002835628329657479, -0.0025842754182717215, 
    -0.0022859362427695004, -0.0019461053054673314, -0.0015710362740026195, 
    -0.0011675586540646069, -0.00074290915849628753, -0.00030456640996465644, 
    0.00013989472093040085, 0.00058294497849741575, 0.0010172178007067331, 
    0.0014356033890683829, 0.0018313275816723284, 0.0021979931148957349, 
    0.0025296181420568827, 0.0028206944728868927, 0.0030662842968731093, 
    0.0032621826475105415, 0.0034051547102482214, 0.0034932036738703392, 
    0.0035258478388036263, 0.0035043278027032682, 0.0034317152528166822, 
    0.0033128677993569731, 0.0031542256483643354, 0.0029634567553678769, 
    0.0027489915579169272, 0.002519494413042769, 0.0022833265022639093, 
    0.0020480667666881408, 0.0018201322443764996, 0.0016045387014659857, 
    0.0014047910397568951, 0.0012228968088364379, 0.001059468418456423, 
    0.00091387784007490938, 0.00078442978875638313, 0.00066855759301221037, 
    0.00056303771442813564, 0.00046424748589544561, 0.00036849931125390855, 
    0.00027242198976986553, 0.00017339951789221238, 6.9975830732072169e-05, 
    -3.779733168192752e-05, -0.00014816181085254031, -0.0002576328376987882, 
    -0.00036118960921611694, -0.0004526820807132418, -0.00052539387281041235, 
    -0.00057272688203095865, -0.0005888908817701015, -0.00056952952323659602, 
    -0.00051218948915935703, -0.00041659164857544699, 
    -0.00028466637357242412, -0.00012038193817163979, 7.06129537926518e-05, 
    0.00028147037009377846, 0.00050469288183187841, 0.00073266415803926793, 
    0.00095812020550806848, 0.0011745086721576437, 0.0013762108142174781, 
    0.0015586494390029571, 0.0017182815785550946, 0.0018525355234162643, 
    0.0019597181407767007, 0.0020389394549149165, 0.002090081151500603, 
    0.002113805809656537, 0.0021115985398231741, 0.0020858179435986513, 
    0.0020396787691354459, 0.0019771619119193324, 0.0019028293197439869, 
    0.0018215490703396252, 0.0017381647250508294, 0.0016571510502064533, 
    0.001582317647657097, 0.0015165651329377122, 0.0014617269988166622, 
    0.0014185056212335048, 0.0013864983503482527, 0.0013643161684704784, 
    0.0013498038284380891, 0.0013403276523641862, 0.0013330894558266355, 
    0.0013254578936344253, 0.0013152528155506683, 0.0013010107293311922, 
    0.0012822041659051272, 0.0012593851690156684, 0.0012342219812576829, 
    0.0012093919259562132, 0.0011883412440510353, 0.0011749534623999643, 
    0.0011731750409019973, 0.0011866393168700326, 0.0012183092498392861, 
    0.0012701490798962905, 0.0013428547589027153, 0.0014356848796927913, 
    0.0015464407823279117, 0.0016716262433037134, 0.0018068037884703561, 
    0.0019470995102339637, 0.0020877673009059377, 0.0022247294969773563, 
    0.0023549929298125496, 0.0024768601755377245, 0.0025899243790172793, 
    0.0026948480495898011, 0.0027929823365655092, 0.0028858656790644774, 
    0.0029747072432193722, 0.0030599012127932022, 0.0031406374004282422, 
    0.0032146629025225117, 0.0032782110055995703, 0.0033261144057201166, 
    0.0033521048589769328, 0.0033492572870040932, 0.003310567363212506, 
    0.0032296065317146184, 0.0031011778582335299, 0.0029219162052821412, 
    0.002690769371013777, 0.0024092682741224192, 0.0020815748955098504, 
    0.0017142813915971024, 0.0013159941408956255, 0.00089674425965858076, 
    0.0004672860197575203, 3.8374892773227181e-05, -0.00037991504263425646, 
    -0.00077877238898925623, -0.0011510764402425007, -0.0014916578285829474, 
    -0.0017973879047393964, -0.0020671068151813217, -0.0023014192802538248, 
    -0.0025023889493040272, -0.0026731785904112113, -0.0028176829491018832, 
    -0.0029401938021234625, -0.0030451060768018436, -0.0031366793985349523, 
    -0.0032188375138467256, -0.0032949997169504238, -0.0033679126078169212, 
    -0.0034394869435223864, -0.0035106527229028846, -0.0035812233731506802, 
    -0.0036498192193143903, -0.0037138437142004033, -0.0037695630026232368, 
    -0.0038122864216166971, -0.0038366724671245254, -0.0038371291113221766, 
    -0.0038082844597813869, -0.0037454904947995847, -0.0036452865819477133, 
    -0.0035057996366674835, -0.0033270085628462876, -0.0031108524491803295, 
    -0.0028611897557287774, -0.0025835918832970554, -0.0022850027585438115, 
    -0.0019732840966859761, -0.001656672367581468, -0.0013431889434398819, 
    -0.0010400310299544995, -0.00075303991388577776, -0.00048627800445314909, 
    -0.0002418014247246292, -1.965090231193531e-05, 0.00018195357597082496, 
    0.00036623017160029793, 0.00053734517206769034, 0.00069989353639809276, 
    0.00085839231593212988, 0.0010168564181417578, 0.0011784537878306413, 
    0.0013452445034839583, 0.0015179851591971716, 0.0016959981695327051, 
    0.0018771073314865225, 0.0020576679200307955, 0.0022327053744987837, 
    0.0023962121512130061, 0.0025415946176636189, 0.0026622701039781828, 
    0.0027523511347775304, 0.0028073483095220082, 0.0028247905299058516, 
    0.0028046723683341863, 0.0027496172448800765, 0.002664740150600317, 
    0.0025572274232454097, 0.0024356811113459085, 0.002309351079755407, 
    0.0021873550709294244, 0.0020779916090999705, 0.0019882087399552043, 
    0.001923258572544894, 0.0018865489520509273, 0.0018796363808098915, 
    0.0019023521852399301, 0.001953000467926969, 0.0020285970354819425, 
    0.0021251390551530248, 0.0022378592558407436, 0.002361457177749758, 
    0.0024903039109271745, 0.0026186059013994802, 0.0027405391210294635, 
    0.0028503754975236083, 0.002942589516828735, 0.00301198376988933, 
    0.0030538184193962354, 0.003063963716218789, 0.0030390644042199355, 
    0.0029767382787877564, 0.0028757708602409728, 0.0027362999663329188, 
    0.0025599653393791654, 0.0023499758239281148, 0.0021110792543177488, 
    0.0018494026384847594, 0.0015721483131070938, 0.00128716307359427, 
    0.0010024364803109455, 0.0007255723800078769, 0.0004633076498977162, 
    0.00022114622569497782, 3.1141375331315553e-06, -0.00018835787983060903, 
    -0.00035242658711069652, -0.00048976290597923838, 
    -0.00060239916645867886, -0.00069352563345166185, 
    -0.00076722170305227461, -0.0008281216858190215, -0.0008810172485327753, 
    -0.00093042626854198513, -0.00098016806003345999, -0.0010329645838629111, 
    -0.0010901349571589549, -0.0011514164260394966, -0.0012149265726675426, 
    -0.0012772759194145933, -0.0013338090949666364, -0.0013789619060035182, 
    -0.0014066977916318629, -0.0014109865433084273, -0.0013862895882395781, 
    -0.0013280245137137566, -0.0012329631995849689, -0.0010995528065329771, 
    -0.00092815526444041006, -0.00072116285386144663, 
    -0.00048298669243557494, -0.00021992212722983718, 6.0140853326797492e-05, 
    0.00034811396787212624, 0.00063418883910760582, 0.00090834547589939093, 
    0.0011608579554745245, 0.001382722959425046, 0.0015660067979483664, 
    0.0017041142826493157, 0.0017919691645600761, 0.001826131776417429, 
    0.0018048880478288665, 0.0017282963211798202, 0.0015981889786019772, 
    0.0014181389637600243, 0.0011933564811226903, 0.00093051960292308742, 
    0.0006375437252527942, 0.00032327317796110902, -2.8752212871862768e-06, 
    -0.00033132052025412029, -0.00065274180909551105, 
    -0.00095850592472945654, -0.0012410629839891931, -0.0014942935741755418, 
    -0.0017137515848070618, -0.0018968012987482378, -0.0020426231168204027, 
    -0.0021520767015235252, -0.0022274443388226347, -0.0022720722235373618, 
    -0.0022899806393020744, -0.0022854935591833316, -0.0022629368494209443, 
    -0.0022264381190400702, -0.0021798361244970664, -0.0021266872756603552, 
    -0.002070312760773357, -0.0020138586682369834, -0.0019603187507395291, 
    -0.0019124723301657944, -0.0018727459530749142, -0.0018429835675485941, 
    -0.001824199189246195, -0.0018163440911358436, -0.0018181564755301559, 
    -0.001827148128515694, -0.0018397312069631884, -0.0018514893593150666, 
    -0.0018575683092432779, -0.0018531346737899982, -0.0018338651126234725, 
    -0.0017964235848935881, -0.0017388783414576964, -0.0016610249501875531, 
    -0.0015645500656897406, -0.0014530262989341449, -0.0013317045354035231, 
    -0.0012071453060634044, -0.0010867568891664487, -0.00097829548601238042, 
    -0.00088938087668886858, -0.00082708267607676232, 
    -0.00079755771588453856, -0.00080576577473731863, 
    -0.00085522343865655943, -0.00094778927173331791, -0.0010834879323478059, 
    -0.0012603798717623058, -0.0014744864354316412, -0.0017198095981932593, 
    -0.0019884780429089252, -0.0022710396855175055, -0.0025569293069051305, 
    -0.0028350918081254902, -0.0030947352878109191, -0.0033260996122372421, 
    -0.0035211995860922173, -0.0036744106162849822, -0.003782845600982329, 
    -0.0038464584065241768, -0.0038678484790955914, -0.0038517954556199796, 
    -0.0038045611605226981, -0.003733081384468746, -0.0036441470383634625, 
    -0.0035436823648810306, -0.0034362091351167225, -0.003324540828087157, 
    -0.0032097412739536578, -0.0030913426198744334, -0.0029677843974454973, 
    -0.0028369991701724414, -0.0026970482057382048, -0.0025466839737782092, 
    -0.0023857333088984616, -0.0022152603197449485, -0.0020375120315008132, 
    -0.001855679708800336, -0.0016735691373161153, -0.0014952251469980945, 
    -0.0013245920490913396, -0.0011652411505983992, -0.0010201772831813574, 
    -0.00089172574093962064, -0.00078151057117726349, 
    -0.00069049957083468433, -0.00061913448615800342, 
    -0.00056748532687440293, -0.00053542737422032454, 
    -0.00052277188421061228, -0.00052930339082911545, 
    -0.00055474117613942703, -0.00059863066347324526, 
    -0.00066023049416246099, -0.00073845536247486767, 
    -0.00083189544833401437, -0.00093890699122994067, -0.0010577099164491212, 
    -0.0011864466689582188, -0.0013231465421209121, -0.0014655957578965306, 
    -0.0016111612400628386, -0.0017566457185586347, -0.0018982685043111005, 
    -0.0020318379151938932, -0.0021531084580603196, -0.002258265120466479, 
    -0.0023444247673996017, -0.0024100063337749579, -0.0024548864056385521, 
    -0.0024803313916929486, -0.0024887303772115339, -0.0024832046984093938, 
    -0.0024671851908969812, -0.0024440362263103027, -0.0024167999743577423, 
    -0.0023880467616644477, -0.002359804606726335, -0.002333540479030042, 
    -0.0023101472121141897, -0.002289961171981885, -0.002272814883846013, 
    -0.0022581282207173843, -0.0022449939389418299, -0.0022322520257794546, 
    -0.0022185246275920199, -0.0022021974542426109, -0.002181377389582653, 
    -0.0021538234950566515, -0.0021168661960701595, -0.0020673261581125452, 
    -0.0020014911313527891, -0.0019152124746910824, -0.0018041773466498916, 
    -0.0016643648233177644, -0.0014926277465120085, -0.0012872540877749818, 
    -0.001048401013292261, -0.00077828717282053795, -0.00048112947702145967, 
    -0.00016283909720099006, 0.00016943490537016902, 0.00050784219550289978, 
    0.00084438538357424053, 0.0011714288838809601, 0.0014821393962645879, 
    0.0017708264183126433, 0.0020331723763490832, 0.0022663479636965333, 
    0.0024689982493673402, 0.0026411202054912445, 0.0027838562892404718, 
    0.0028991952719726547, 0.0029896555372356812, 0.0030579345237332499, 
    0.0031066084696732468, 0.0031378792634638307, 0.0031534098469836107, 
    0.003154244315878236, 0.0031408227308077682, 0.00311304982062481, 
    0.0030704099559934095, 0.0030120949274217634, 0.0029371310213236967, 
    0.0028445095465923602, 0.002733326856765157, 0.0026029253449735236, 
    0.0024530661209476831, 0.0022841261706588326, 0.0020973275042546263, 
    0.0018949593522941768, 0.0016805551876880164, 0.0014589802612595881, 
    0.001236352463709226, 0.001019773398961652, 0.00081689663892490225, 
    0.00063539304278596742, 0.00048238160804766456, 0.00036388661772678656, 
    0.00028437289213183241, 0.00024639705845377218, 0.00025036340221327384, 
    0.00029441830521059802, 0.00037447947148063984, 0.00048439451863223424, 
    0.00061625713891769814, 0.00076090693770103411, 0.00090858759957703297, 
    0.0010497146004407095, 0.0011756763277061264, 0.0012795445734342494, 
    0.0013565938444776214, 0.0014045229281320617, 0.0014233248588152384, 
    0.0014148430780352187, 0.0013820671791425761, 0.0013283202692908861, 
    0.001256498473903858, 0.0011685133840670732, 0.0010650295004620257, 
    0.00094555550893452066, 0.0008088343373822347, 0.00065342961656886288, 
    0.00047834426776773996, 0.00028351802201580874, 7.0080764446640381e-05, 
    -0.00015967158721932957, -0.00040252458007460984, 
    -0.00065471111933294401, -0.00091231201474164961, -0.0011715665806317571, 
    -0.0014290679895753674, -0.0016818086836815544, -0.0019271108520600921, 
    -0.0021624800925521314, -0.0023854326196988142, -0.0025933683764176501, 
    -0.002783498544116652, -0.0029528822749701148, -0.0030985651347080916, 
    -0.0032178060984465687, -0.0033083360596467275, -0.0033686315244358979, 
    -0.0033981087704077883, -0.0033972470233733453, -0.0033675812508664848, 
    -0.0033115654382820745, -0.0032323375820061686, -0.003133422106017773, 
    -0.0030184175933352514, -0.0028907050595613397, -0.0027532305052193357, 
    -0.0026083583832251112, -0.0024578281805512667, -0.0023027550455625317, 
    -0.0021436993468179825, -0.0019807482001660552, -0.0018136185748666017, 
    -0.0016417366642594933, -0.00146430237783093, -0.0012803122778574519, 
    -0.0010886022786269574, -0.00088788005935175167, -0.00067680457824866036, 
    -0.00045411468166365226, -0.00021879824577318964, 2.9737936747276539e-05, 
    0.00029154806611750598, 0.00056609087332663898, 0.00085228277926584998, 
    0.0011486382792926756, 0.0014534486091833309, 0.0017649665352930349, 
    0.0020815540795198133, 0.0024017463699872372, 0.0027242309106325462, 
    0.0030477384299270518, 0.0033708430782525144, 0.0036917205124797421, 
    0.0040078993865542752, 0.0043160509863964152, 0.0046118908411519593, 
    0.004890215396863613, 0.0051450953028365325, 0.0053702161416071727, 
    0.005559326974895481, 0.0057067551109639377, 0.0058079055851913445, 
    0.0058597283884918305, 0.0058610977442461881, 0.0058130711264206191, 
    0.0057189849814935278, 0.0055843696508781106, 0.0054166587793049968, 
    0.0052246953848730697, 0.0050180593722276455, 0.0048062771602008052, 
    0.0045979852437878698, 0.0044001671833595853, 0.0042175258718695763, 
    0.0040520901910408771, 0.00390308011244367, 0.0037670507395625771, 
    0.0036382937780263958, 0.0035094607913409102, 0.0033723353143137965, 
    0.0032186833650608964, 0.0030410547638277208, 0.0028334697204460422, 
    0.0025919221467316238, 0.0023146294750647483, 0.0020020880612163202, 
    0.0016569027429122946, 0.0012834550606495413, 0.00088749699089125434, 
    0.00047569183354981, 5.5171958623239075e-05, -0.00036685419466726056, 
    -0.00078342187598008195, -0.0011880704976579535, -0.0015750452018382446, 
    -0.0019394245608286458, -0.0022772020293594843, -0.0025852987917005668, 
    -0.0028615064693053548, -0.0031043613314862295, -0.0033130048097527037, 
    -0.003487063167828043, -0.0036266128926038597, -0.0037322284250430071, 
    -0.003805136551567034, -0.0038474104531529283, -0.0038621330391280773, 
    -0.003853443190945046, -0.003826419046694052, -0.0037867799336627813, 
    -0.0037404326084724505, -0.0036929114775236978, -0.0036487874303207301, 
    -0.0036111207893435773, -0.0035810668265506161, -0.003557691301133412, 
    -0.003538044415433878, -0.0035174976008563747, -0.0034902635718916078, 
    -0.0034500543634817904, -0.0033907615785432315, -0.0033070530426862169, 
    -0.0031948316162015286, -0.0030515252339567973, -0.0028761736330317231, 
    -0.0026693478234764466, -0.0024329020364882571, -0.0021696463511366548, 
    -0.0018829740209834035, -0.0015765304897817733, -0.0012539810820196918, 
    -0.00091891255390008251, -0.00057487117129523583, 
    -0.00022548600310351528, 0.00012535790106042472, 0.00047339841967366798, 
    0.00081395657933567797, 0.0011420189923552699, 0.0014524197903509743, 
    0.0017400746201194756, 0.0020002332327428872, 0.0022286974663909644, 
    0.0024219803761014163, 0.0025774328298562672, 0.0026932918056062206, 
    0.0027686931351092992, 0.0028036749839817875, 0.002799160630359984, 
    0.0027569339323291774, 0.0026796108078336301, 0.0025706245641736862, 
    0.0024341783793892218, 0.0022751762613454655, 0.002099120512806747, 
    0.0019119853909767971, 0.0017200822162572397, 0.0015299686029965078, 
    0.0013483637689848795, 0.0011820373986793232, 0.0010376552534326158, 
    0.00092155668016044166, 0.00083944509004303799, 0.0007960389195488843, 
    0.00079465798919281885, 0.00083682787328242527, 0.00092192349606527431, 
    0.0010469196150462725, 0.0012063270768930899, 0.0013923521327215145, 
    0.0015952904425758903, 0.001804150606427257, 0.0020074076950144662, 
    0.0021938385298494799, 0.0023533186254288941, 0.0024775184265430376, 
    0.0025604137726256103, 0.0025985958878960657, 0.0025913490765478056, 
    0.0025405362486428181, 0.0024502985921346166, 0.0023266165682957053, 
    0.0021767312491067906, 0.0020084920237367545, 0.001829628309387183, 
    0.0016470279971747739, 0.0014660853506626628, 0.0012901974187810913, 
    0.0011205024342665466, 0.00095588069975871038, 0.00079325598982375701, 
    0.00062813794886105393, 0.00045533436352379858, 0.00026976497193889214, 
    6.7235414785557263e-05, -0.00015487815624745725, -0.00039713120736434532, 
    -0.0006577593716665368, -0.00093268739811290784, -0.0012157894075901948, 
    -0.0014993213398532903, -0.0017745313182481702, -0.0020323054205186875, 
    -0.0022638336028518303, -0.0024612315449258548, -0.0026181275816901644, 
    -0.0027301445126543923, -0.0027952607151198691, -0.0028140073654084122, 
    -0.0027894112708703009, -0.0027267051107260033, -0.002632762330955921, 
    -0.0025153517838922635, -0.0023823113855928986, -0.0022408045066778584, 
    -0.0020967284347179868, -0.0019543388152910629, -0.001816080836562908, 
    -0.0016826110993954473, -0.0015529186878191932, -0.001424571583338989, 
    -0.0012940810669111603, -0.0011574047955634544, -0.0010105926872079091, 
    -0.00085048732757416336, -0.00067535999996772358, 
    -0.00048533347740642614, -0.00028255085697801639, 
    -7.1078173065922459e-05, 0.00014340296125348712, 0.00035406229033898586, 
    0.00055348204956777989, 0.00073423596750067308, 0.00088943083646754234, 
    0.0010131836532633744, 0.0011009599073655242, 0.0011497737194005988, 
    0.0011582508519506363, 0.0011265170359919217, 0.0010559604843225633, 
    0.00094891784398730612, 0.00080828994963252757, 0.00063722701911862007, 
    0.00043887409524763358, 0.0002162915516572032, -2.7487194487846498e-05, 
    -0.00028928374398040516, -0.00056553848321890237, 
    -0.00085208391565062738, -0.0011439807654477707, -0.0014354193278645873, 
    -0.0017197408178309212, -0.0019895393116655465, -0.0022368791315877132, 
    -0.0024536053932719126, -0.0026317003453171367, -0.0027636886763026916, 
    -0.0028430418055205848, -0.0028645569734614459, -0.0028246890395173373, 
    -0.0027218169614752754, -0.0025564227697606997, -0.0023311937742435621, 
    -0.0020509701354258082, -0.0017225991600192687, -0.0013546329731469293, 
    -0.00095692389457266045, -0.00054008478259554515, 
    -0.00011489727809268872, 0.00030829118998405662, 0.00072012802651619549, 
    0.001112734284713107, 0.0014799832770640538, 0.0018176307897249159, 
    0.0021232373536964185, 0.0023959160857875959, 0.0026359408587646499, 
    0.0028442538109538147, 0.0030219045495246746, 0.003169510360657104, 
    0.0032868241120148573, 0.0033725145366446624, 0.0034242864969622937, 
    0.0034392859658957616, 0.0034147693582978764, 0.0033488565317057587, 
    0.0032411760146076152, 0.0030932937218278397, 0.0029088480323665837, 
    0.0026934187151341966, 0.002454171512428592, 0.0021993573040104695, 
    0.0019377527411473456, 0.00167806724704551, 0.0014284100087128134, 
    0.0011958804528247428, 0.00098631242878803615, 0.00080417811397784161, 
    0.0006526531912244924, 0.00053379882209463134, 0.00044876040067801787, 
    0.00039797629433420032, 0.0003812886083506295, 0.00039799679704206892, 
    0.0004468127432134606, 0.00052578156622631368, 0.00063218175875691418, 
    0.000762491943935495, 0.00091242589068370455, 0.001077097930273426, 
    0.0012512957282438775, 0.0014298277733413892, 0.0016078518269006495, 
    0.0017811050823042264, 0.0019460014241080104, 0.0020995758082279731, 
    0.0022393604979703608, 0.0023632699505228946, 0.0024695487467628467, 
    0.0025568176628639884, 0.0026241722651709856, 0.002671295348964211, 
    0.0026984759741364118, 0.0027065147302595335, 0.0026965079635315648, 
    0.002669546830022098, 0.0026264089340446465, 0.0025673117224213234, 
    0.0024917845756610674, 0.0023986861122304156, 0.0022863528274091691, 
    0.002152893132361128, 0.0019966087196171228, 0.0018164811259793383, 
    0.0016126960756702171, 0.0013871136314967489, 0.001143592919444111, 
    0.00088808542905190776, 0.00062845484022937183, 0.00037401927226454203, 
    0.0001348587116190165, -7.8968032626708471e-05, -0.00025819859720287511, 
    -0.00039500340156207211, -0.00048341251062409348, 
    -0.00051952157814828229, -0.00050146306146362277, 
    -0.00042923032359371027, -0.00030439082214530559, -0.0001297216538774452, 
    9.1147595860207611e-05, 0.00035405333037332061, 0.00065456945474539241, 
    0.00098818332791246466, 0.0013503826024469589, 0.0017366157016396285, 
    0.002142192103802966, 0.0025621233668597261, 0.0029910203085417599, 
    0.0034230364121173289, 0.0038518902937595594, 0.0042709706833092397, 
    0.0046734683644437582, 0.0050525423627886005, 0.0054014713907361081, 
    0.0057137986854108374, 0.0059834499886899798, 0.0062048839869432819, 
    0.0063732243089437892, 0.006484487805281762, 0.0065358286897676792, 
    0.0065258294406986004, 0.0064547629398588845, 0.0063248253997478538, 
    0.0061402404320171832, 0.0059071822269209737, 0.0056335499102822938, 
    0.0053285712648807404, 0.0050023200093219375, 0.0046652212072584116, 
    0.0043276190639826339, 0.0039994246346430661, 0.0036897930006778755, 
    0.0034067603580309495, 0.0031568511616738471, 0.0029446872437755419, 
    0.0027727860806785391, 0.0026415946669479723, 0.0025497768183909827, 
    0.0024947373845652463, 0.0024731592451076685, 0.0024815173037161485, 
    0.0025164099008428689, 0.0025747007481702498, 0.0026534420552995377, 
    0.002749755730661304, 0.0028606681062431616, 0.0029830496413559004, 
    0.0031136662262290422, 0.0032493127398042949, 0.0033869470195191163, 
    0.0035237818858633251, 0.0036572993518150213, 0.0037851753064041347, 
    0.0039051520175832442, 0.0040149142232256468, 0.0041119712796983086, 
    0.0041935844149517641, 0.0042567060500693886, 0.0042979683887168739, 
    0.0043137194152565294, 0.0043001186934626782, 0.0042533656353833469, 
    0.0041700092295255285, 0.0040473627196323941, 0.0038839266658912798, 
    0.0036798011106118061, 0.0034369911027482174, 0.0031595682868648988, 
    0.0028536529178087707, 0.0025271663071587576, 0.0021893805866621918, 
    0.0018502183803434523, 0.0015194501922497911, 0.0012058394779392075, 
    0.000916402451717154, 0.00065585581313017029, 0.00042641195410089521, 
    0.00022792184244145954, 5.830568462628625e-05, -8.5771575558121348e-05, 
    -0.00020818061221288616, -0.00031263752580468099, 
    -0.00040217992388866307, -0.00047883655490617945, 
    -0.00054348859843984419, -0.00059592910247362153, 
    -0.00063503770889788242, -0.00065906619139788781, 
    -0.00066598555618570861, -0.00065385460752341552, 
    -0.00062113171594059731, -0.00056692218431567533, 
    -0.00049111235793274826, -0.00039440186517027251, 
    -0.00027827891216211051, -0.00014493827836892177, 2.8372133087443659e-06, 
    0.0001618557052127463, 0.0003286872829678316, 0.00049985156129477633, 
    0.00067198432021026199, 0.00084193170677006714, 0.0010067495707274075, 
    0.0011636312232316149, 0.0013097742295799125, 0.0014422174398731494, 
    0.0015577396203412515, 0.0016527851827272159, 0.0017234708671474402, 
    0.001765722250602334, 0.0017754782860831646, 0.0017490332969173213, 
    0.0016834517710326647, 0.0015770091258934303, 0.0014296964861134902, 
    0.0012436757125633567, 0.0010235403669360038, 0.00077629700838219122, 
    0.00051096383811541509, 0.00023786639391253935, -3.2188150411365597e-05, 
    -0.00028883889263877093, -0.00052291248024257742, 
    -0.00072699441884078574, -0.00089582339245615765, -0.0010264545511681536, 
    -0.0011182561737774724, -0.0011727599973120524, -0.0011932809957087437, 
    -0.0011843423262733552, -0.0011510201581363629, -0.001098211340004229, 
    -0.0010300086610176709, -0.00094922933199326903, -0.00085723110928685644, 
    -0.00075400889022426705, -0.00063853261828397526, 
    -0.00050925850295490413, -0.00036471120059370071, 
    -0.00020407204814883607, -2.762456996763907e-05, 0.00016295332866359306, 
    0.00036449844657482561, 0.00057249004303597619, 0.00078133126863180269, 
    0.00098482033996870897, 0.001176735283221332, 0.0013515472488145473, 
    0.0015051304708634042, 0.0016353598834336208, 0.0017424634243049283, 
    0.0018290957009790196, 0.0018999849080759204, 0.0019612887108294411, 
    0.0020197230173823462, 0.0020815621332912924, 0.0021516728211332966, 
    0.0022327005118715584, 0.0023245017958079062, 0.0024239360818786183, 
    0.0025250064313491697, 0.0026193371804302768, 0.002696868175512119, 
    0.0027467261270227856, 0.0027580950491414287, 0.0027210543162930929, 
    0.0026273816832122999, 0.0024712558422538525, 0.0022499250515846171, 
    0.0019642822244313714, 0.0016192019870152744, 0.0012235978805719156, 
    0.00079015142422602237, 0.00033463398511487469, -0.00012509500785467184, 
    -0.00057036786408829572, -0.00098312769727004843, -0.0013473546549529619, 
    -0.001650327919660467, -0.0018835496542069542, -0.0020432361741756421, 
    -0.0021302411955037744, -0.0021495271534214132, -0.0021092688071301649, 
    -0.0020197564212928024, -0.0018922979430235349, -0.0017382289552556889, 
    -0.0015681463606964235, -0.0013913721596961353, -0.001215658971699863, 
    -0.001047080033157689, -0.00089003752306201838, -0.00074738530845014513, 
    -0.00062057376633681456, -0.00050980539256347663, 
    -0.00041419799312372978, -0.00033192816294641265, 
    -0.00026041442241997827, -0.00019643524532545528, 
    -0.00013631531897132486, -7.6078825282798845e-05, 
    -1.1638034376600646e-05, 6.1053004263093825e-05, 0.0001458491289952628, 
    0.00024635301229561282, 0.00036584601163292126, 0.00050719225407429432, 
    0.00067265457080466478, 0.00086363602169988005, 0.0010804808994266694, 
    0.001322391744515419, 0.001587512643252121, 0.0018730877895287862, 
    0.0021757359303545849, 0.0024916929539779979, 0.002817042671338487, 
    0.0031478518461869956, 0.0034802003622463641, 0.0038101133800221374, 
    0.0041334329597025972, 0.00444572037946809, 0.0047421919398400363, 
    0.0050177397445438044, 0.0052670499540461452, 0.0054847594022657351, 
    0.0056656788123102264, 0.0058050578264432278, 0.0058989156025045873, 
    0.0059443929337603604, 0.0059401490468671608, 0.0058867126574385018, 
    0.0057866829838645788, 0.005644726402437213, 0.0054673422494296254, 
    0.0052623119858000071, 0.0050379590131047992, 0.0048022270505671755, 
    0.0045618471388567047, 0.0043216569408985805, 0.0040842238939396572, 
    0.0038498533945356727, 0.0036169443369990506, 0.0033826157130173017, 
    0.0031435211623464434, 0.0028965712346569346, 0.0026394876866799068, 
    0.0023710174589071588, 0.0020907944889552599, 0.0017989935186959699, 
    0.0014958925970069148, 0.0011816356285638918, 0.0008561871981136429, 
    0.00051947517748944429, 0.00017153015405267365, -0.00018748567704753071, 
    -0.0005573720132512523, -0.00093804225459485587, -0.001329716187635161, 
    -0.0017330535006945377, -0.0021491526284913923, -0.0025792970586902119, 
    -0.0030244292633364832, -0.0034844438757599076, -0.0039573411493676125, 
    -0.0044385103703820511, -0.0049203040079588414, -0.0053920814003379286, 
    -0.0058407776618586218, -0.0062519349787246272, -0.0066110281982433745, 
    -0.0069047928260006141, -0.0071224360985327716, -0.0072565045274424513, 
    -0.0073033156143533428, -0.0072630376497845404, -0.0071394046791869413, 
    -0.0069392130923894568, -0.0066716333194705929, -0.0063474138643694489, 
    -0.005977966712910501, -0.0055744673968242909, -0.0051470382419156642, 
    -0.0047041130441699535, -0.0042521018564883372, -0.0037953712698108118, 
    -0.0033365276640472978, -0.0028768383391124621, -0.0024168396170751202, 
    -0.0019568875059383876, -0.0014976402092780161, -0.00104037327669228, 
    -0.00058713004485231603, -0.00014073557148412859, 0.00029538618825614355, 
    0.00071755312509770835, 0.0011222863197567279, 0.0015068195252697391, 
    0.0018695554206802859, 0.0022103526646268272, 0.00253054194400427, 
    0.0028326360715502444, 0.0031198568216857427, 0.0033954262601085627, 
    0.0036618074166475593, 0.0039198805517276017, 0.0041682753589295405, 
    0.0044028498129037785, 0.0046164554746005561, 0.0047991339342515014, 
    0.0049387307266668011, 0.0050219813065927668, 0.005035807896989551, 
    0.0049686965351805595, 0.0048118904893399619, 0.0045602958937845193, 
    0.0042130142305504392, 0.0037735494146664845, 0.0032497783302133706, 
    0.0026536329249298852, 0.0020005569840333337, 0.0013086712485269468, 
    0.00059776507887149472, -0.00011191032832120719, -0.00080082673416608094, 
    -0.0014512770712824365, -0.002048272210213187, -0.0025801319742950178, 
    -0.0030387775410871962, -0.0034197546170955133, -0.0037221090576264157, 
    -0.0039481276607912768, -0.0041031087878990952, -0.0041950780219270475, 
    -0.004234430344162838, -0.0042334722453599722, -0.004205741477755303, 
    -0.0041651637639931148, -0.0041250725115675752, -0.0040971969957257484, 
    -0.0040907013469895859, -0.0041113742916906683, -0.0041611391716136394, 
    -0.0042378353735993586, -0.0043354249613244099, -0.0044445324907238211, 
    -0.0045532989427595058, -0.0046483885229595323, -0.0047160339362367935, 
    -0.0047429954129459013, -0.0047173180511122324, -0.0046288939384286354, 
    -0.0044698546467140778, -0.0042347656281177025, -0.0039207994101261379, 
    -0.0035279131833148652, -0.003059015126200406, -0.0025201980394876315, 
    -0.0019209238071170919, -0.0012742183695249366, -0.00059675705666549072, 
    9.1288391639085011e-05, 0.00076669441090287276, 0.0014041055365190188, 
    0.001977326934645056, 0.0024610647027233654, 0.0028327993366221932, 
    0.0030745053494247057, 0.0031739883070314653, 0.0031256270952998762, 
    0.0029304398300437416, 0.0025955157783636587, 0.0021330640403890103, 
    0.0015591678491166843, 0.00089264170340513471, 0.00015409378358423396, 
    -0.00063465422055889082, -0.0014508964176728747, -0.0022712160221045122, 
    -0.003071683814531065, -0.0038281327795266153, -0.0045166087877585841, 
    -0.0051140507339895594, -0.0055992532309140901, -0.0059542558116274652, 
    -0.0061660770836651588, -0.0062284046622238277, -0.0061428363225614875, 
    -0.0059192923836242509, -0.0055754927020150776, -0.0051356942516548433, 
    -0.0046291293854028356, -0.0040882575350899304, -0.0035468742520913523, 
    -0.0030378955996419503, -0.0025909278762304882, -0.0022300434112663579, 
    -0.0019719098025358052, -0.0018248254212626612, -0.0017886382814701566, 
    -0.0018554403375937558, -0.0020110006429337754, -0.0022365951906396305, 
    -0.0025110834044858271, -0.0028128492586160523, -0.0031214893610062885, 
    -0.0034190159913937601, -0.003690679352082179, -0.0039251756633105015, 
    -0.0041147512056509423, -0.0042549621513874192, -0.0043442440119725598, 
    -0.0043832488402746781, -0.0043740651300123671, -0.0043194645186625724, 
    -0.0042223954122475775, -0.0040857341730698585, -0.0039123828910926795, 
    -0.0037055545071837744, -0.0034690867898119733, -0.0032075994148042472, 
    -0.0029265561248341698, -0.0026321609340840923, -0.0023312525062849751, 
    -0.0020313311318747376, -0.0017406503876097002, -0.0014683778671470723, 
    -0.0012246889787770503, -0.0010207376871959502, -0.00086836614450193274, 
    -0.00077957816501133983, -0.00076581895218175784, 
    -0.00083725531748788718, -0.0010021907003005517, -0.0012667145429252494, 
    -0.0016345067429311014, -0.0021068563312280808, -0.0026827492235851538, 
    -0.0033587117220607939, -0.0041285525442627596, -0.0049827637857332236, 
    -0.005907691216414471, -0.0068847179509141316, -0.0078896759547167905, 
    -0.0088931857489297876, -0.0098619249041611741, -0.010760983024642234, 
    -0.011556683154606432, -0.012219416529943789, -0.012725782018418313, 
    -0.013059942150280109, -0.013213983244754675, -0.013187589348474161, 
    -0.012987221714159551, -0.012625043069822149, -0.012117801630667523, 
    -0.011485778820855146, -0.010751703400910643, -0.0099399153908166157, 
    -0.0090756063466274958, -0.0081842552095918522, -0.0072913676725483668, 
    -0.0064222399310724385, -0.0056016824313880435, -0.0048536296778588827, 
    -0.0042000701755954819, -0.0036597381911126752, -0.0032462504008693013, 
    -0.0029664797110678853, -0.0028193094155333775, -0.002795228021489217, 
    -0.0028769893333596111, -0.0030407145233864578, -0.0032576207326471341, 
    -0.0034957331667563487, -0.0037215245634988911, -0.0039014822772914215, 
    -0.0040032842350977271, -0.0039969412582813481, -0.0038557105898223269, 
    -0.0035571597617840029, -0.0030841716523682529, -0.0024260933216523946, 
    -0.0015796393168825049, -0.00054945215685112819, 0.00065190799398554065, 
    0.0020047781369878855, 0.0034839608194305654, 0.0050606987982898732, 
    0.006704760839446061, 0.0083864006075572619, 0.010077695504160371, 
    0.011753238614464824, 0.013390193582785242, 0.014967809663941362, 
    0.01646644649509079, 0.017866405214117097, 0.019146324470595777, 
    0.020281772141712836, 0.021244562021503127, 0.022002839401263165, 
    0.022522507190035426, 0.022769573377824363, 0.02271273556714172, 
    0.022325733830307538, 0.021588606116392559, 0.020488428254736957, 
    0.019020141315728423, 0.017187726777079894, 0.01500629276430409, 
    0.012504570516365473, 0.0097272517742835844, 0.0067358292260531263, 
    0.0036073980905398369, 0.00043102291866485305, -0.0026981863267825598, 
    -0.0056859790769471161, -0.0084456279136587258, -0.010903355556141248, 
    -0.013002262774741027, -0.014705135238613784, -0.015995808903269695, 
    -0.016879833072177122, -0.017383825888883573, -0.017553101613341674, 
    -0.017447908586744991, -0.017138259254015003, -0.01669771545801137, 
    -0.016197559021316636, -0.015701017846644738, -0.015258853719230627, 
    -0.014906655504055741, -0.014663849461977701, -0.014535000846173011, 
    -0.01451307809211135, -0.01458420397812844, -0.01473293086990678, 
    -0.014945460020226949, -0.015209649997592311, -0.015511490974066721, 
    -0.015830031368277993, -0.016131282932699702, -0.016365927263963631, 
    -0.016471709154731836, -0.01638004872340167, -0.016024210426298958, 
    -0.015347418779698953, -0.014308392476516654, -0.012884500778506801, 
    -0.011074345842700091, -0.0088987783614594765, -0.006401006875634602, 
    -0.0036461239357004644, -0.00071858107880149596, 0.0022833673313506515, 
    0.0052550711875631552, 0.0080950107778271999, 0.010712091086507163, 
    0.013035549480802483, 0.01501402770296025,
  // Fqt-F(8, 0-1999)
    1, 0.99102138416827901, 0.96463576717844379, 0.92243368367988321, 
    0.86686754409292788, 0.80098732787222182, 0.7281351877208414, 
    0.65164491384048828, 0.57458517422061273, 0.49957212731092204, 
    0.42866144635871262, 0.36331576844431585, 0.30443365185044508, 
    0.25242105078117222, 0.20728590183526188, 0.16873914922362168, 
    0.13628998227822828, 0.10932799948737135, 0.087189030069327933, 
    0.069204438578761296, 0.054735601237664175, 0.043195970220226504, 
    0.034063354368881874, 0.026884777834852745, 0.021275941385286292, 
    0.016916975524842958, 0.013545798229439146, 0.010950262495818852, 
    0.0089600121837636309, 0.0074387619245389301, 0.0062775517340094939, 
    0.0053891985830201482, 0.0047040201145118424, 0.0041666841990865089, 
    0.0037339378988998882, 0.0033729127258162557, 0.0030597568059702852, 
    0.0027783882777858812, 0.002519290814837663, 0.0022783171598860078, 
    0.002055516716754253, 0.0018539940001253829, 0.0016788127577049355, 
    0.0015359208872554951, 0.0014310598013276082, 0.0013687189941926697, 
    0.0013511656285307636, 0.0013776806606985259, 0.0014441125245507006, 
    0.0015428367311818728, 0.0016631659851141132, 0.0017922052292964107, 
    0.0019160482963322789, 0.0020211651401428172, 0.002095776015455208, 
    0.0021309998207740496, 0.0021215972802451884, 0.0020662013247084339, 
    0.0019670616239611271, 0.0018293716114432263, 0.001660381316026526, 
    0.0014684757187982316, 0.001262369459468012, 0.0010504924197126558, 
    0.00084058564660195235, 0.00063944428700646772, 0.00045277588136862624, 
    0.00028514136386086092, 0.00013994491061412591, 1.9485724219022067e-05, 
    -7.4941469578468909e-05, -0.00014286030083158607, 
    -0.00018440147451100899, -0.00020007873146046562, 
    -0.00019061364980727468, -0.00015683046805198947, -9.959165071678829e-05, 
    -1.9797201235120256e-05, 8.157827095311022e-05, 0.00020339323668489722, 
    0.00034417110693446312, 0.00050186608453790436, 0.00067358660900291353, 
    0.00085532591795128387, 0.0010417807020143559, 0.0012263191465389448, 
    0.0014011698826092063, 0.0015578271324141228, 0.001687681808008381, 
    0.0017827845192441164, 0.0018366755482055411, 0.0018451350545778487, 
    0.0018067702068779317, 0.0017233236285053458, 0.0015996657118130583, 
    0.0014434207123875428, 0.001264293851246183, 0.0010731563658617242, 
    0.00088101525603355348, 0.00069802915079988676, 0.00053268734987954158, 
    0.00039130330062068375, 0.00027784495247244701, 0.00019409500200712795, 
    0.00014005750173635544, 0.00011449849414062126, 0.00011548016701901004, 
    0.00014081039623283745, 0.00018832017183258816, 0.00025597411525655372, 
    0.00034183796300983512, 0.0004439579285806782, 0.00056022913353436833, 
    0.00068830604764159463, 0.00082559748466647185, 0.00096934961347919647, 
    0.0011167783878365035, 0.0012651972569025316, 0.0014120860860189679, 
    0.001555084945119912, 0.0016919086594021854, 0.0018202070469247934, 
    0.0019374102745162638, 0.0020405977740652597, 0.002126439362905381, 
    0.0021912262364568503, 0.0022310091427427659, 0.0022418356190966877, 
    0.0022200302264919428, 0.0021624889056717027, 0.0020669380676786096, 
    0.0019321214596473093, 0.0017578851962085668, 0.0015451858245213277, 
    0.0012960210697799172, 0.0010133352260854663, 0.00070091074975474408, 
    0.00036329297891795568, 5.7384084722300374e-06, -0.00036581071262757625, 
    -0.00074476574998699199, -0.0011239516413935227, -0.0014957443477233111, 
    -0.0018522755795432962, -0.0021857155293915284, -0.0024885959395458354, 
    -0.0027541664224081789, -0.0029767250585555054, -0.0031519221922433568, 
    -0.0032769923891787412, -0.0033509088303805864, -0.0033744187185798949, 
    -0.0033499462797446566, -0.0032813447906775866, -0.0031735118350563868, 
    -0.00303189465295116, -0.0028619535737774179, -0.0026686597159577582, 
    -0.0024561043457385959, -0.0022272960727688193, -0.0019841610954759604, 
    -0.0017277317003304934, -0.0014584493604665317, -0.0011764996348832522, 
    -0.00088209595147597803, -0.00057563648844792114, 
    -0.00025776435042812874, 7.0661580386943658e-05, 0.00040858107632998073, 
    0.00075467188819022531, 0.0011071617726992708, 0.0014635115746514786, 
    0.0018200399226072775, 0.0021715857977565112, 0.0025113433165606892, 
    0.0028309271319259246, 0.0031207260417683482, 0.0033705056873711441, 
    0.0035702435735098133, 0.0037110842106663497, 0.0037863215311851189, 
    0.0037922725195199316, 0.0037288982957921339, 0.0036000588478935225, 
    0.003413315720347298, 0.0031793077031643893, 0.0029107568346084965, 
    0.0026212635155313446, 0.0023240590196429347, 0.0020308800901633161, 
    0.00175109559604879, 0.001491178167094069, 0.0012545248594780546, 
    0.0010416104986864306, 0.00085040377833156869, 0.00067695955552153945, 
    0.00051610548748668209, 0.00036213619185549578, 0.00020947052504686394, 
    5.3229685156376528e-05, -0.00011029703876883037, -0.00028331800291520894, 
    -0.00046634739273934662, -0.00065817879168527933, 
    -0.00085601240440143721, -0.0010557066946263909, -0.0012521313059697347, 
    -0.0014395696593189284, -0.0016121322507055456, -0.0017641522795704251, 
    -0.0018905426259284814, -0.0019870803104999005, -0.0020506134035446159, 
    -0.0020791739629785013, -0.0020719863570150534, -0.0020293738092580994, 
    -0.0019525886998390859, -0.0018435830182585468, -0.0017047893599582741, 
    -0.0015389241909332407, -0.0013488506417546171, -0.0011374991312001457, 
    -0.00090784899691094935, -0.00066293946166127581, 
    -0.00040588407832388657, -0.00013989851084945346, 0.0001316788351701406, 
    0.00040533439468629724, 0.00067732310487045777, 0.00094360317836752572, 
    0.0011997909352237206, 0.0014411831221352151, 0.001662863499422013, 
    0.001859910428693246, 0.002027677308772262, 0.0021621092167766745, 
    0.0022600419794503424, 0.00231942045524352, 0.0023394182121194004, 
    0.0023204286496144996, 0.0022639549144563872, 0.0021724152772672786, 
    0.0020489307567942766, 0.0018971169704226393, 0.0017209233155235826, 
    0.0015245248989907811, 0.0013122859947568102, 0.0010887626940228236, 
    0.00085873068153219194, 0.00062719693894285489, 0.00039939872985506568, 
    0.00018077099294065902, -2.3102310529410342e-05, -0.00020656101510106945, 
    -0.00036396790298632637, -0.00048985661626839276, 
    -0.00057913660611633915, -0.00062734223866421429, 
    -0.00063093216270674744, -0.00058758879637562343, 
    -0.00049650988464667038, -0.00035864985181705542, 
    -0.00017687361462524816, 4.3975582764065416e-05, 0.00029712995707008164, 
    0.00057406463307068463, 0.00086481954793512204, 0.0011584482304196515, 
    0.0014435939253244282, 0.0017091659010035213, 0.0019450583563868818, 
    0.0021428484070341227, 0.0022964052017990888, 0.0024023417684767155, 
    0.0024602627808337483, 0.0024727777430611172, 0.0024452878400578948, 
    0.0023855438201692124, 0.0023030242430053869, 0.0022081458379909894, 
    0.0021113681892671516, 0.0020222307273985206, 0.0019484090512934241, 
    0.0018948679927775615, 0.0018632243328518192, 0.0018514244694573341, 
    0.0018538098677529447, 0.0018615995697814438, 0.0018637661785361546, 
    0.0018481820484332657, 0.001802922744473956, 0.0017175165277954145, 
    0.0015840094911413456, 0.0013977033400429785, 0.0011575016462940456, 
    0.00086585652697351856, 0.0005283658423721082, 0.00015313789824270834, 
    -0.00024996029917651372, -0.00067003485062033482, -0.0010957765495858776, 
    -0.0015159302985499671, -0.0019196232729866741, -0.0022966267218676832, 
    -0.0026376431149855639, -0.0029346545948816674, -0.0031813397307863369, 
    -0.0033735291364277867, -0.0035095784907796818, -0.0035905741637735715, 
    -0.0036202756677651857, -0.0036047442823675586, -0.0035517392749899526, 
    -0.003470002093543523, -0.003368565416314711, -0.0032561945353896393, 
    -0.0031409938604154909, -0.0030301777350835611, -0.0029299669952970939, 
    -0.002845571262542276, -0.0027811683254172124, -0.0027398881975083116, 
    -0.002723736867294292, -0.0027335104816628517, -0.0027687320921146179, 
    -0.0028276554607886608, -0.002907365098561294, -0.0030039704330186395, 
    -0.0031128941090535632, -0.0032291914114676509, -0.0033478499903774077, 
    -0.0034640348535765566, -0.0035732260590840993, -0.0036712698507365251, 
    -0.0037543540049455645, -0.0038189462846526232, -0.0038617523870155715, 
    -0.0038797047039606323, -0.003870009381298686, -0.0038302497968350935, 
    -0.0037585068572330645, -0.0036534803964553509, -0.0035145663018264889, 
    -0.0033418820941980799, -0.0031362584980488416, -0.0028992014603061922, 
    -0.0026328895136331931, -0.0023402229133662974, -0.0020249404938467268, 
    -0.0016917418138920933, -0.0013463646528446822, -0.00099552702073187559, 
    -0.0006466990017315288, -0.00030770218129549395, 1.3815358193235166e-05, 
    0.00031094989485828576, 0.00057808433101993041, 0.00081128540186412577, 
    0.001008497731002266, 0.0011695056834496711, 0.0012956779588001947, 
    0.0013895205416297762, 0.0014541538245750928, 0.0014927703990030474, 
    0.0015081720701327172, 0.0015024271806037862, 0.0014767254320995271, 
    0.0014314281201552798, 0.0013662989323613463, 0.0012808734975459893, 
    0.0011749118816590039, 0.0010488370731752436, 0.00090413733831597729, 
    0.00074365498036124016, 0.00057174398789667299, 0.0003942694299860093, 
    0.00021844415946982123, 5.2486367420950732e-05, -9.4886314205547972e-05, 
    -0.00021509088353949333, -0.00030040126909029649, -0.0003446412153258159, 
    -0.00034379022939446421, -0.0002964096181813649, -0.00020383589011088314, 
    -7.0155438086532432e-05, 9.8054989528630822e-05, 0.00029217092004412597, 
    0.00050213083426430363, 0.00071715942842164471, 0.00092655951790325585, 
    0.0011204809210490828, 0.0012906057680351036, 0.0014306586746473762, 
    0.0015367230152771758, 0.0016073394466353413, 0.0016434115062493419, 
    0.0016479413407759235, 0.0016256424543774016, 0.0015824681983386377, 
    0.0015251082696581444, 0.0014604849434912226, 0.0013952927867913513, 
    0.0013355905784790221, 0.0012864568184167509, 0.0012517086828582799, 
    0.0012336694889671909, 0.0012329810630386745, 0.0012484704375393197, 
    0.0012770830154189641, 0.0013139281856680443, 0.0013524780101741619, 
    0.0013849390405011822, 0.0014028124775977381, 0.0013976004157583845, 
    0.0013615873695953995, 0.0012885990922957156, 0.0011746506715607141, 
    0.0010184099585468897, 0.00082143614653653252, 0.00058820426922844948, 
    0.00032588724049155101, 4.393488844803479e-05, -0.00024653585948757609, 
    -0.00053349683809256144, -0.00080481072260456363, -0.0010489947212576616, 
    -0.0012558600981284415, -0.0014169544263997187, -0.0015257960769784081, 
    -0.0015779204928874962, -0.0015708157639042384, -0.001503813192839619, 
    -0.0013780271993811685, -0.0011963776831445342, -0.00096369766681004491, 
    -0.00068687693375120516, -0.00037498635961346428, 
    -3.9282236037470027e-05, 0.00030695544409232328, 0.00064881374706789066, 
    0.00097037000386812221, 0.0012555566694098302, 0.0014892336845146409, 
    0.0016583771837264875, 0.0017532397211443625, 0.0017682825157404949, 
    0.0017026901412020511, 0.0015603820288514108, 0.0013495737916966919, 
    0.0010819816640061626, 0.00077183073469075023, 0.00043475953526001237, 
    8.6738565954887171e-05, -0.00025695673674111725, -0.00058261557708059347, 
    -0.00087878585502770801, -0.0011367164730615399, -0.0013505767845434363, 
    -0.0015174202083423874, -0.0016369468877398729, -0.0017111300174988396, 
    -0.0017437326180422771, -0.001739778148186055, -0.0017049983743252541, 
    -0.0016452994473586521, -0.0015662581762542721, -0.0014726911602320958, 
    -0.001368334984724616, -0.0012556621652297835, -0.0011358706982894883, 
    -0.0010090478825123391, -0.00087447768767486684, -0.00073104820201726575, 
    -0.00057770780195734971, -0.00041387755414372174, 
    -0.00023978297810927935, -5.6640556963788159e-05, 0.0001333251878349939, 
    0.00032703547394578446, 0.00052084795484432607, 0.00071092247704064766, 
    0.00089360762933691563, 0.0010657656112927649, 0.0012249783424631015, 
    0.001369600398539086, 0.0014986622361245173, 0.0016116490969779282, 
    0.0017082173541833169, 0.0017879266394154316, 0.0018500813504888746, 
    0.0018937187785908851, 0.0019177712075271053, 0.0019213773485888606, 
    0.0019042799534179234, 0.0018671851992677231, 0.0018120229689115267, 
    0.0017419895888616966, 0.0016613625997473438, 0.0015751451650488895, 
    0.0014885873752643216, 0.0014066856783227961, 0.0013337324267348133, 
    0.0012729706233794542, 0.0012263849991768587, 0.0011946906960251665, 
    0.0011775006639065811, 0.0011736434698745751, 0.0011815610208685901, 
    0.0011996684295978886, 0.0012266006759478764, 0.0012612647097854299, 
    0.0013026900959807047, 0.0013497363724397186, 0.0014007403355216885, 
    0.0014532171787389986, 0.0015037242837263392, 0.001547976699726943, 
    0.0015812234481159869, 0.001598837972380268, 0.0015970126137325846, 
    0.001573409998596835, 0.0015276268644159189, 0.0014613724291454952, 
    0.0013783485605205652, 0.001283848990486118, 0.0011841455558832651, 
    0.0010857421187108075, 0.00099458546890376248, 0.0009153188307507858, 
    0.0008507114924059644, 0.00080135860633344749, 0.00076574631534681538, 
    0.00074066225685236729, 0.00072186953102461283, 0.00070487359417576107, 
    0.00068564628845010499, 0.00066117859787891121, 0.00062981283411039056, 
    0.00059130621175929564, 0.00054667311273479341, 0.0004978158181747302, 
    0.00044704181937354174, 0.00039654450020717974, 0.00034794863924990219, 
    0.000301997522190185, 0.00025843017478594877, 0.00021605169368313029, 
    0.00017295639038686578, 0.00012681086227036908, 7.5130231016319864e-05, 
    1.5450841602969358e-05, -5.4573395420360959e-05, -0.00013714452240314831, 
    -0.00023429779125770948, -0.00034780131536279318, -0.0004789482752053297, 
    -0.00062823161936786259, -0.00079494202657027742, 
    -0.00097680426754991252, -0.0011697295024699402, -0.0013678102595408412, 
    -0.0015635687745859041, -0.0017484366952703956, -0.0019134057032559554, 
    -0.0020497565934432358, -0.0021497683023880554, -0.0022073273407836446, 
    -0.0022183858426132867, -0.0021812107077784975, -0.002096385694399309, 
    -0.0019665878999134984, -0.0017961795486665978, -0.0015906809339946647, 
    -0.0013562352444174922, -0.0010991612142096428, -0.0008256648093302977, 
    -0.00054170601379426638, -0.00025303723883425875, 3.4689419270462932e-05, 
    0.0003157671099384056, 0.00058434282607696102, 0.00083441810385905728, 
    0.0010599672863854091, 0.0012551701751829592, 0.0014147327752874357, 
    0.001534251083525654, 0.0016105773703323021, 0.0016421492414719159, 
    0.0016292500664638206, 0.0015741830532566693, 0.001481319809849938, 
    0.0013570194379246114, 0.0012093893891170135, 0.0010478897681540926, 
    0.00088280912305854818, 0.00072464269815618451, 0.00058343205434886649, 
    0.00046814694828944199, 0.0003861554765601917, 0.00034283809957176385, 
    0.0003413843312337541, 0.00038276678528777311, 0.00046586235471177947, 
    0.00058767111651594783, 0.00074357087273183844, 0.00092756218020035534, 
    0.0011324953936004858, 0.0013503032473175956, 0.001572244927728022, 
    0.0017891964264773641, 0.0019920126400368825, 0.0021719460393854724, 
    0.0023211170179662038, 0.002432988705754906, 0.0025027968037043442, 
    0.0025278564932455592, 0.0025077320634615289, 0.0024442275138556635, 
    0.0023412065100866463, 0.0022043002962040818, 0.0020405283695780836, 
    0.0018578768126179895, 0.0016648619479930301, 0.0014700881058005123, 
    0.0012818222640309609, 0.0011075878409390763, 0.00095379304264852597, 
    0.00082543039302728426, 0.0007258679264883737, 0.00065675132729148657, 
    0.00061798529972978866, 0.00060779925719410912, 0.00062285448006580845, 
    0.00065840779763092167, 0.00070853207411375051, 0.00076639104998231511, 
    0.00082458786010226534, 0.00087556529178920372, 0.00091207443889507048, 
    0.00092766902567440856, 0.00091721943468067962, 0.00087738201309290839, 
    0.00080696947513691033, 0.00070713978176839207, 0.00058136165780829597, 
    0.00043512824700666578, 0.00027542063420379827, 0.00010999119982795008, 
    -5.3450934862759767e-05, -0.00020803049082133635, 
    -0.00034836547218064322, -0.00047100352848244618, 
    -0.00057456898225984661, -0.00065963723812602186, 
    -0.00072833847380585168, -0.00078376992861230611, 
    -0.00082931680972719293, -0.00086794667856883098, 
    -0.00090159820114085526, -0.000930716426231344, -0.00095399601838590047, 
    -0.00096836898269068278, -0.00096923069471599498, 
    -0.00095090655263284384, -0.00090728477030246489, 
    -0.00083257086138469906, -0.00072204266717251536, -0.0005726844895350972, 
    -0.00038360444129889484, -0.00015618539586354164, 0.00010603736784407011, 
    0.00039764648575662116, 0.00071171923820578017, 0.0010402035645683059, 
    0.0013742589070920533, 0.0017046159207824763, 0.0020219678395464813, 
    0.0023174176473766878, 0.0025829837756282158, 0.0028120981510109814, 
    0.002999997558106351, 0.0031439173268276305, 0.0032430709694196468, 
    0.0032984018030664838, 0.0033121799341807056, 0.0032875334137407882, 
    0.0032279903576082321, 0.0031371202767607707, 0.0030183089958361639, 
    0.0028746962746523459, 0.0027092717118539721, 0.0025250817343638421, 
    0.0023254624439174561, 0.0021142079826467477, 0.0018956325049969056, 
    0.0016744982656053437, 0.0014558461910337034, 0.0012447735960295695, 
    0.0010461910318952973, 0.00086458124516256474, 0.00070374108342853114, 
    0.00056655223589487753, 0.00045480744434693164, 0.00036916641570234286, 
    0.00030924539308667788, 0.0002738381748512087, 0.00026120063099636058, 
    0.00026931950988505737, 0.0002960625574223543, 0.00033919957693243042, 
    0.00039630077572376873, 0.00046459421214328919, 0.0005408719233584566, 
    0.00062153003342235399, 0.00070279072829150351, 0.00078107340224577409, 
    0.00085344714071113319, 0.00091804829663797035, 0.00097432794938541434, 
    0.0010230193492626648, 0.0010658051550297008, 0.0011046944799214453, 
    0.001141229628067778, 0.0011756890290437238, 0.0012064883949920145, 
    0.0012299397580320059, 0.0012404618481995616, 0.0012312139452798777, 
    0.0011950727818355079, 0.001125752901628147, 0.0010188647937211621, 
    0.00087271920673642138, 0.00068875509246691194, 0.00047153852223039426, 
    0.00022837578704058053, -3.1367331140329973e-05, -0.00029715152925028428, 
    -0.00055817875173910531, -0.00080427416445263749, -0.0010266157678278907, 
    -0.001218258526308818, -0.0013744258023871039, -0.001492583693587514, 
    -0.0015723442050313678, -0.001615243572148488, -0.001624422036911373, 
    -0.0016042365631830507, -0.0015597944179255418, -0.0014964727225650421, 
    -0.0014194895082438278, -0.0013335932241594661, -0.0012428790536649691, 
    -0.0011507632132339812, -0.001060018303549163, -0.00097284638887078234, 
    -0.00089092308029218973, -0.0008153763764106954, -0.00074672491990271372, 
    -0.00068481454102398923, -0.0006287933714865801, -0.00057717501071610322, 
    -0.00052805669119352456, -0.00047947683936240087, 
    -0.00042990479782532593, -0.00037873400725030949, 
    -0.00032664436985459526, -0.00027569342009838905, 
    -0.00022906684327266382, -0.00019048732429925795, 
    -0.00016340204599123116, -0.00015014136761621678, -0.000151222942891812, 
    -0.00016500663179555515, -0.00018772736044412084, 
    -0.00021395098762297361, -0.00023731128021924053, 
    -0.00025138455345364755, -0.00025051487108991197, 
    -0.00023045615242135454, -0.00018872497598967225, 
    -0.00012465605961626945, -3.9202879583734415e-05, 6.5441684804731705e-05, 
    0.00018627201583252439, 0.00031986741625010892, 0.00046269557618472325, 
    0.00061129876622641362, 0.00076238836108009781, 0.00091288284739846374, 
    0.0010599436884525205, 0.0012010240485637064, 0.0013339450786317435, 
    0.0014569668655723608, 0.0015688138959252572, 0.0016686201063909659, 
    0.001755798861282219, 0.0018298394792300029, 0.0018901090866492356, 
    0.0019356596342135395, 0.0019650919680402569, 0.0019764684601001553, 
    0.0019672891380886799, 0.0019345530108513321, 0.0018749153720548984, 
    0.0017849816063879222, 0.0016617173931969841, 0.0015029475961525819, 
    0.0013078964937643491, 0.0010776703890947501, 0.00081558431524668277, 
    0.00052728565800583727, 0.00022062117258598289, -9.4773988620949247e-05, 
    -0.000408089545971909, -0.00070811534207687772, -0.00098404512565728342, 
    -0.001226221840553239, -0.001426732883772697, -0.0015798071137447744, 
    -0.0016819888721153111, -0.0017321055146932267, -0.0017310626089826425, 
    -0.0016815357398092734, -0.0015876258776313708, -0.0014545220787097011, 
    -0.0012882200276901701, -0.0010952955270467912, -0.00088272106175425248, 
    -0.00065770746041232794, -0.00042750804887482368, 
    -0.00019917853598081073, 2.0693291503661284e-05, 0.00022627592482720902, 
    0.00041276933059654765, 0.00057662964446782974, 0.00071572068062816232, 
    0.00082938540647947343, 0.00091839168286217507, 0.00098476561304665171, 
    0.0010315047823847609, 0.0010622537816240242, 0.0010809972512077269, 
    0.0010918324232596646, 0.001098831686563695, 0.0011059894785068363, 
    0.0011172049805334059, 0.0011362511703131716, 0.0011667166000160272, 
    0.0012118934421191066, 0.0012746241695141313, 0.0013571362472627759, 
    0.0014608901906407992, 0.001586487688096661, 0.0017336368829176186, 
    0.0019011749266469853, 0.0020871123099567173, 0.0022886842209371154, 
    0.0025023752905610347, 0.0027239292823666703, 0.002948354158884353, 
    0.0031699714264517443, 0.0033825216336379558, 0.0035793742661623445, 
    0.0037538598269724389, 0.0038996933673968504, 0.0040114779604178722, 
    0.0040852142357151369, 0.0041187427977239363, 0.0041120500560222744, 
    0.004067364107393172, 0.0039890165542012289, 0.0038830659411073073, 
    0.0037567413331298411, 0.0036177794133071882, 0.0034737390650591993, 
    0.0033313773911229955, 0.0031961158306027279, 0.0030716493390294916, 
    0.0029597277832483539, 0.0028601065041868922, 0.0027707038018077871, 
    0.0026879101470071182, 0.0026070501147622983, 0.0025229385121327249, 
    0.0024305038094225725, 0.0023254023655245684, 0.0022046015193477133, 
    0.002066861332333067, 0.0019130986758016818, 0.0017465749694629451, 
    0.0015729095981367232, 0.0013998682232487442, 0.0012369602574671757, 
    0.0010948390817505842, 0.00098453586970468862, 0.00091658866707643519, 
    0.00090015075819207852, 0.00094217740652859496, 0.0010467616586210865, 
    0.0012147318374256643, 0.0014435224790408567, 0.0017273432243102855, 
    0.0020576017985940403, 0.0024234953017216888, 0.0028126712316992163, 
    0.0032118656801885938, 0.0036074399490996583, 0.0039858006496291702, 
    0.0043337054057388767, 0.0046385665429310701, 0.0048887693026418077, 
    0.0050741033946250591, 0.005186273120561833, 0.0052194908876791301, 
    0.0051710766754513538, 0.0050419818866835678, 0.0048371289245817978, 
    0.0045654449376092273, 0.0042395382009399454, 0.003874971132878084, 
    0.0034891687438141908, 0.0031000753028796366, 0.0027247287012842139, 
    0.0023779707807907425, 0.0020714847203696638, 0.001813327385752242, 
    0.0016079962207287838, 0.0014569908768727738, 0.0013596982358374003, 
    0.0013143837490104892, 0.0013190403353393948, 0.0013719270084434814, 
    0.0014717231321769611, 0.0016173055445535098, 0.0018072707645892887, 
    0.0020393461473624513, 0.0023098234403589029, 0.0026131778451279333, 
    0.0029419190096058589, 0.0032867493738571256, 0.0036369719594441024, 
    0.0039810885293387957, 0.0043075217745378244, 0.004605317098095283, 
    0.0048647399432308683, 0.0050776720535846542, 0.0052377695236532108, 
    0.0053403955236905765, 0.0053823943050826566, 0.005361812085025076, 
    0.0052776882806075242, 0.0051299418825243755, 0.0049194085296810491, 
    0.0046479906502787226, 0.0043189079075785291, 0.0039370132395948228, 
    0.0035090900136598097, 0.0030441196872104566, 0.0025534055902970963, 
    0.00205047722502059, 0.0015507384373720334, 0.0010708087019450484, 
    0.00062764196667637628, 0.00023748282943382275, -8.5195784858087958e-05, 
    -0.00032866087643373888, -0.00048468289052628607, 
    -0.00054903543448817809, -0.00052168285028192699, 
    -0.00040668560836509452, -0.0002118270861270927, 5.1994004156268297e-05, 
    0.00037154064152599125, 0.00073211823949012687, 0.0011184489163256232, 
    0.0015154457118546781, 0.0019087970907978981, 0.0022853611273665041, 
    0.0026334073118026023, 0.0029428048085289003, 0.0032052146690165939, 
    0.0034143593594266131, 0.0035663600546430078, 0.0036600925893897551, 
    0.0036974561757343407, 0.003683422330435887, 0.0036257231841259662, 
    0.0035341921692393268, 0.0034198279574347251, 0.0032937447939756534, 
    0.0031661677065545285, 0.0030455980275373986, 0.002938205595351415, 
    0.0028474781539072061, 0.0027741884630641989, 0.0027166749667943539, 
    0.0026714057950545694, 0.0026337446408404674, 0.0025987913220493816, 
    0.0025621670610602373, 0.0025206298278113524, 0.0024724112537684098, 
    0.0024172253925660281, 0.00235601149836525, 0.0022905267784584971, 
    0.0022229160443614144, 0.0021553757445152972, 0.002089920258952617, 
    0.0020282440451370111, 0.0019716036040041711, 0.0019206660674916836, 
    0.0018753102983749233, 0.0018343706969605768, 0.0017953904989560848, 
    0.001754503485521937, 0.0017066251223669094, 0.0016460518543313233, 
    0.001567411041046391, 0.0014667871330629779, 0.0013427053642190326, 
    0.0011967327453670899, 0.0010335505717196112, 0.00086048492552031881, 
    0.00068662041496927995, 0.00052164284369040498, 0.00037461077194867831, 
    0.00025287687055582011, 0.0001612737422700586, 0.00010170424322218863, 
    7.3147514627259558e-05, 7.2010130308314659e-05, 9.2719019739573099e-05, 
    0.00012840578213273716, 0.0001716038603533819, 0.00021483743870890254, 
    0.0002511153563903435, 0.00027427919110966688, 0.00027924464981120864, 
    0.00026213865291279986, 0.00022037921622362585, 0.00015269670186729924, 
    5.9108485412957785e-05, -5.9141266107214994e-05, -0.00019974091461512467, 
    -0.00035954124553267352, -0.00053487466793554505, 
    -0.00072190122621379178, -0.00091691633559176124, -0.001116539632738894, 
    -0.001317780421861179, -0.0015179704482086902, -0.0017145895286900296, 
    -0.0019050654842738134, -0.0020866177627035312, -0.0022561480862270779, 
    -0.0024102847762025948, -0.0025455875015905063, -0.0026589124176374015, 
    -0.0027478779643255518, -0.0028113162382493234, -0.0028495787444824108, 
    -0.0028646094894858405, -0.0028597625149534974, -0.0028393601945956625, 
    -0.0028081324262278842, -0.0027706190885406182, -0.0027306193232290443, 
    -0.0026907957642236524, -0.0026524334231039044, -0.0026153598838924682, 
    -0.0025780301384011185, -0.0025377431509636698, -0.0024910080927406783, 
    -0.0024339885741486798, -0.0023630525447159104, -0.0022753281585622324, 
    -0.0021692455972140839, -0.0020449088094819765, -0.0019042497687501248, 
    -0.0017508484627269741, -0.0015893855809956726, -0.001424847029937313, 
    -0.0012616376351219554, -0.0011028602772351092, -0.00094997597614248546, 
    -0.00080297166621876048, -0.00066097047007330166, 
    -0.00052308691651100627, -0.00038920715701909887, 
    -0.00026047493657903033, -0.00013932123919169003, 
    -2.9046880423730034e-05, 6.6906514886043374e-05, 0.00014580501360798688, 
    0.00020637772521753053, 0.00024928878892012353, 0.00027722691760225312, 
    0.0002945771662637162, 0.00030673174578692232, 0.00031915638328618666, 
    0.00033640694837812454, 0.00036127716502212798, 0.0003942444345229656, 
    0.00043333834779618564, 0.00047443226441529944, 0.00051193273822473437, 
    0.00053970827914756278, 0.00055212304779723369, 0.00054495541034118916, 
    0.00051610044638879574, 0.00046589574467948119, 0.00039705527758943625, 
    0.00031423989179393412, 0.00022332120279351382, 0.00013048422405557221, 
    4.1297435992313332e-05, -4.012457797977542e-05, -0.00011173215069992226, 
    -0.00017387382780567682, -0.00022927655693149874, 
    -0.00028265515315516518, -0.00034001758091100454, 
    -0.00040773798278580703, -0.00049153124510754073, 
    -0.00059549937768923892, -0.00072139082734929035, -0.0008681658817532318, 
    -0.0010319244918134479, -0.0012062184121199499, -0.0013827115062391591, 
    -0.0015521102272856059, -0.001705308949766948, -0.0018345674190777313, 
    -0.0019345680217160036, -0.0020031987533819348, -0.0020419237310467337, 
    -0.002055640479342992, -0.0020520979410955749, -0.0020409191790321446, 
    -0.0020324153327210396, -0.002036332808282533, -0.0020607701581345111, 
    -0.0021113343191567851, -0.0021906486692022885, -0.0022982242777095097, 
    -0.0024306089627225331, -0.002581755756575117, -0.0027434929481769525, 
    -0.0029060427438956202, -0.0030585414234976221, -0.0031895930816473544, 
    -0.0032878343051805448, -0.0033425610764506132, -0.0033443891474075498, 
    -0.0032859179205259829, -0.0031623203105296148, -0.002971798683419514, 
    -0.0027158480064698605, -0.0023992705146612539, -0.0020299718043769043, 
    -0.0016185429357700718, -0.001177702497842513, -0.00072161796155981249, 
    -0.0002652018371877569, 0.00017664564842454964, 0.00058979053829264958, 
    0.00096161365549391809, 0.0012817393295529592, 0.0015427002592290793, 
    0.0017404591503580042, 0.0018747678632678685, 0.0019492640009533949, 
    0.0019712799839240311, 0.0019513047044369448, 0.0019021659903689855, 
    0.0018379619631171897, 0.0017728877631597803, 0.0017200667530134063, 
    0.0016905286360987997, 0.0016924094984725935, 0.0017304389726452507, 
    0.0018057248365795893, 0.0019158369492579229, 0.0020551828396211834, 
    0.0022156189254399494, 0.0023872981865109243, 0.0025596161320642057, 
    0.002722212249902105, 0.0028658738552582341, 0.0029832835186037825, 
    0.0030695323507480394, 0.0031223908892047719, 0.0031423438987793428, 
    0.003132415838152909, 0.0030978422373203703, 0.0030455921937954621, 
    0.0029837535361300063, 0.002920778284863609, 0.0028645828613121341, 
    0.0028215688927444725, 0.0027956449069771582, 0.0027874228564930938, 
    0.0027937452115739153, 0.0028076747144125938, 0.0028190381288791914, 
    0.0028155039504803277, 0.0027840918115102451, 0.0027128827830025255, 
    0.0025926830632881049, 0.0024183433798333947, 0.0021895703806559881, 
    0.0019111160372736354, 0.0015923440175129541, 0.0012463301122499675, 
    0.00088861620732209412, 0.00053584924788518051, 0.00020446231853953696, 
    -9.0463653789593255e-05, -0.00033603615089040212, -0.0005220867546020737, 
    -0.00064139828702901064, -0.00068970694655245252, 
    -0.00066548921981430457, -0.00056968692826619646, 
    -0.00040537841161032739, -0.00017747666072623759, 0.00010755368664060053, 
    0.00044194363863132565, 0.0008168348581199681, 0.0012225391323498142, 
    0.0016487935042230465, 0.0020850431366363836, 0.0025207270411843406, 
    0.0029455546882562879, 0.003349758169622056, 0.0037243441711232879, 
    0.0040613367266392232, 0.0043540311508028784, 0.0045972170591149948, 
    0.0047873635408868858, 0.0049226813665161637, 0.005003030255238447, 
    0.0050296675537883353, 0.005004839792806158, 0.0049313131199509516, 
    0.0048119498715402352, 0.0046494000139882538, 0.0044460213546818235, 
    0.0042040076444974607, 0.0039257162462938908, 0.0036141268865740577, 
    0.0032733370291380668, 0.0029089433141435113, 0.0025281512823564223, 
    0.0021395108155785793, 0.0017522721043472973, 0.0013755048859469703, 
    0.0010171859166061346, 0.0006834476872264086, 0.00037811909855015046, 
    0.00010261779406821163, -0.00014384915005948175, -0.0003638001905557731, 
    -0.00056077763296284429, -0.00073857050329147959, 
    -0.00090049516167218396, -0.0010489564920747963, -0.0011853358931175598, 
    -0.0013102172128719911, -0.0014238598757250428, -0.00152677627804411, 
    -0.001620225351383368, -0.0017064882388689723, -0.001788812083723521, 
    -0.0018710099505953193, -0.0019567432244252422, -0.0020486353037339495, 
    -0.0021474120779032806, -0.0022513067018093136, -0.002355891151615665, 
    -0.0024543946182442487, -0.0025384887347327414, -0.0025993873854928133, 
    -0.0026290639120136795, -0.002621408438809739, -0.0025731774605986784, 
    -0.002484625834054459, -0.0023597932145219035, -0.0022063818568449399, 
    -0.0020352670867371555, -0.001859643418635214, -0.0016939425946025264, 
    -0.0015525768722583172, -0.0014486676688819239, -0.0013928988763180468, 
    -0.0013926131723067049, -0.0014512607089526377, -0.0015681860375126237, 
    -0.0017387908517530366, -0.001954974471350822, -0.0022057776607879477, 
    -0.0024781508301334881, -0.0027577865731216143, -0.0030299734587575055, 
    -0.0032804421954147024, -0.003496147576503128, -0.0036659137616302574, 
    -0.0037808590888870745, -0.0038346170410520678, -0.0038234000926531996, 
    -0.0037460157347664366, -0.0036038789749372473, -0.0034009874432986815, 
    -0.0031438482153572688, -0.0028412237654612603, -0.0025037148805559903, 
    -0.0021431625277446419, -0.0017719413212394551, -0.0014021818533810086, 
    -0.0010450468448974918, -0.00071008187779332131, -0.00040481271848636312, 
    -0.0001345909616960327, 9.7233581103998968e-05, 0.00028890039298035418, 
    0.00043964020836671276, 0.00054911409830248655, 0.00061697163323329047, 
    0.00064270338861475756, 0.00062573885778769724, 0.00056576638405106557, 
    0.00046318014318215157, 0.00031951475929781843, 0.00013781189581452594, 
    -7.7166534342468831e-05, -0.00031887823437119474, 
    -0.00057911006285356532, -0.00084821776847055017, -0.0011154495062421039, 
    -0.0013693494301270559, -0.0015982056227695266, -0.0017905177460129317, 
    -0.0019355216024052871, -0.0020236899728076256, -0.0020472263212729319, 
    -0.0020005229780686142, -0.0018805775451039787, -0.0016873577798525734, 
    -0.0014240968644647926, -0.0010975533329436618, -0.00071813574926102471, 
    -0.00029984225768580589, 0.00014010471060328691, 0.00058197435457087838, 
    0.0010046214752082491, 0.0013868820803086821, 0.0017091768206714778, 
    0.0019551010463913494, 0.0021128483073584487, 0.0021762255483620155, 
    0.0021451728026503965, 0.0020256774607279628, 0.0018291489335521885, 
    0.0015712977570937782, 0.001270732500584727, 0.00094733143072205897, 
    0.0006206477192909933, 0.00030843726402676101, 2.5446355910483092e-05, 
    -0.00021745570885504207, -0.00041373287831290037, 
    -0.00056115975694597073, -0.00066133182772776581, 
    -0.00071871009459521372, -0.00073946510153916479, 
    -0.00073030750490978946, -0.00069748679518616885, 
    -0.00064612774552137567, -0.00057988545971187147, 
    -0.00050094464484580319, -0.0004102561940541637, -0.00030794587695224309, 
    -0.00019377737119856002, -6.7557150439242434e-05, 7.0553780223966923e-05, 
    0.00021984531330386233, 0.00037898085009062702, 0.00054597248553197491, 
    0.00071822710102832274, 0.00089260344855618965, 0.0010655214411040815, 
    0.0012331411795284957, 0.0013916299776819533, 0.001537499241664122, 
    0.0016679968384290015, 0.0017814533410300201, 0.0018775405919953412, 
    0.0019573493265082399, 0.0020232492296566522, 0.0020784938618613894, 
    0.0021266215556780309, 0.002170678042758709, 0.0022123733741155555, 
    0.0022512881805960396, 0.0022843361075381621, 0.002305588872611656, 
    0.00230655350357197, 0.0022769314357354692, 0.0022057224960420662, 
    0.0020825340323420032, 0.0018989200020599062, 0.0016495403518291668, 
    0.00133296985525967, 0.00095211958751923917, 0.00051413558419558046, 
    2.9874370891398206e-05, -0.00048704398804367546, -0.0010214118937685076, 
    -0.0015577052806235794, -0.0020812859131095246, -0.0025793556408178885, 
    -0.0030416478062689433, -0.0034608040861308781, -0.003832482500436071, 
    -0.0041552336151293749, -0.0044302225088033798, -0.0046608385494716683, 
    -0.0048522381898425514, -0.0050108995821217354, -0.0051441177496099498, 
    -0.0052595161087884241, -0.0053644780520668766, -0.00546560806047357, 
    -0.0055682172518701726, -0.0056759286552017021, -0.0057904885017328687, 
    -0.0059117541547483955, -0.0060378510641421511, -0.006165414400203551, 
    -0.0062898684615506637, -0.0064057508063613371, -0.006507026408277659, 
    -0.0065874390083336589, -0.0066409343208741964, -0.0066620592352462206, 
    -0.0066463990883664208, -0.006590953337782879, -0.0064944450042677153, 
    -0.0063574956858345162, -0.0061826456517641371, -0.0059742678429222651, 
    -0.0057383126553675846, -0.0054819611699044131, -0.0052131535993007148, 
    -0.0049399844813269346, -0.0046699553738688152, -0.0044091618671506143, 
    -0.0041615606672023584, -0.0039283996849655348, -0.0037079779680832575, 
    -0.0034957756864636767, -0.0032849541584301432, -0.0030671708094849727, 
    -0.0028335739328775563, -0.0025757551177719345, -0.0022865713486446633, 
    -0.0019607090526936673, -0.0015950029230866367, -0.0011885353045757987, 
    -0.00074262193735423932, -0.00026076185908044906, 0.00025140306392469196, 
    0.00078617745466098171, 0.0013340294485054197, 0.0018839230867047604, 
    0.0024237765275485256, 0.0029408660381752935, 0.0034221696639039323, 
    0.0038547130377097364, 0.0042259838397478034, 0.0045245638494097289, 
    0.0047409230436884064, 0.004868325087300414, 0.0049036892902717868, 
    0.0048482526922608137, 0.0047078724505998587, 0.0044928079087478891, 
    0.0042170553533551845, 0.003897231301311328, 0.003551235653611289, 
    0.0031968460967834503, 0.0028504321499576543, 0.0025259011247180715, 
    0.0022339561854145306, 0.0019817000351817888, 0.0017725685733062482, 
    0.001606636998162246, 0.0014811252582980746, 0.0013910717342113697, 
    0.0013300190154215939, 0.0012906320739319837, 0.0012651903341144026, 
    0.0012460617933770487, 0.0012261734349213777, 0.0011995903542095223, 
    0.001162154886936273, 0.0011120857702905478, 0.0010503952260823173, 
    0.00098094343299674151, 0.0009100603676254112, 0.00084570366509089995, 
    0.00079627512550536428, 0.00076932564082671608, 0.00077041245862475953, 
    0.0008023691957112811, 0.00086522037463768772, 0.00095671397328299271, 
    0.0010732948445354587, 0.0012112635822100729, 0.00136773485678975, 
    0.0015411631812842835, 0.0017312484062276235, 0.0019382995240874714, 
    0.0021621286629555547, 0.0024008462425012984, 0.0026497786203368741, 
    0.0029008165541214897, 0.0031423430209579725, 0.0033598319879707137, 
    0.0035370165743213015, 0.0036574625425703678, 0.0037062944474343224, 
    0.0036717141400525446, 0.0035460953055781608, 0.0033264898697400527, 
    0.0030145484944569443, 0.0026159211583394477, 0.002139363812075495, 
    0.0015958088066650208, 0.00099752919288611944, 0.00035755130703641187, 
    -0.00031076808133239547, -0.00099402576570946171, -0.0016790404364175292, 
    -0.0023531155997983909, -0.0030043392807792327, -0.003621872249010939, 
    -0.0041961813148666, -0.0047192009388096409, -0.0051844323583519949, 
    -0.0055870278399894578, -0.0059238477161854576, -0.0061934637183098367, 
    -0.0063960281994354792, -0.006532945026114843, -0.0066064746281598447, 
    -0.0066195071533151368, -0.0065755789231135096, -0.0064791752879499627, 
    -0.0063359980812946982, -0.0061529606149179619, -0.0059378392566979462, 
    -0.0056985813667988936, -0.0054424541759685117, -0.0051752350280799501, 
    -0.0049005463297489942, -0.0046194426993292495, -0.0043303385072276587, 
    -0.0040292531751870741, -0.0037104603435156856, -0.0033674300452967119, 
    -0.0029939147235808978, -0.0025850170214267113, -0.0021380317735455899, 
    -0.0016529429030785331, -0.0011325130645122104, -0.0005820116745328777, 
    -8.6480297035568775e-06, 0.00057908511603205648, 0.0011720430899455334, 
    0.0017609462470190621, 0.0023366816359187146, 0.0028903893684073716, 
    0.0034134840036456177, 0.0038976406081980297, 0.0043348911794198744, 
    0.004717746410199496, 0.0050392604097100622, 0.0052929846014994333, 
    0.0054726951123152592, 0.0055720505388002425, 0.0055843021043191637, 
    0.0055022729389032389, 0.005318743407887112, 0.0050273434118276493, 
    0.004623811035884883, 0.0041074815264291169, 0.0034826777230061515, 
    0.0027597357771320602, 0.0019553400341267685, 0.0010921018709857929, 
    0.00019730844806968952, -0.00069893075881847003, -0.001565913383828611, 
    -0.0023745722616214807, -0.0030994338413033967, -0.0037201115310511795, 
    -0.0042222415605492822, -0.0045978294363215825, -0.004845060447118253, 
    -0.0049676882667886802, -0.0049741248532973849, -0.004876292019136667, 
    -0.0046884188288731513, -0.0044259094234540631, -0.0041044250738567298, 
    -0.0037392379020246822, -0.0033448524163399301, -0.0029346806315748934, 
    -0.0025207152258193951, -0.0021131350410012917, -0.0017198719259052038, 
    -0.001346167259181957, -0.00099425472121326573, -0.00066325491094057238, 
    -0.00034938762297805244, -4.647347650830032e-05, 0.00025324646417279395, 
    0.00055807345964239215, 0.00087573320768025609, 0.0012123195749142866, 
    0.0015714588509473154, 0.0019537525846933931, 0.0023566473512692874, 
    0.0027747181507904255, 0.0032003211704061453, 0.003624488458156288, 
    0.0040379110729721083, 0.0044318621085851877, 0.0047989407895129505, 
    0.0051336496043819548, 0.0054327876343137479, 0.0056957397999537586, 
    0.0059246317591215916, 0.0061242782644224314, 0.0063017908594072986, 
    0.0064657921986326413, 0.0066252703656353518, 0.0067882476087945216, 
    0.0069604876939149771, 0.0071444147124055044, 0.0073384211861886629, 
    0.0075366654244553993, 0.0077294281871146354, 0.0079039837999642804, 
    0.0080459074632561953, 0.0081405752739512529, 0.0081745968973930168, 
    0.0081369952234566657, 0.0080199314466886194, 0.0078189596269783983, 
    0.0075329092100427158, 0.0071634676575217642, 0.0067146494802316622, 
    0.0061921356984371845, 0.0056025693983702534, 0.0049529214687172116, 
    0.004250025186696196, 0.0035003975205209546, 0.0027104339599176904, 
    0.0018868787839305869, 0.0010375724730016524, 0.00017220468714545091, 
    -0.00069707534770810419, -0.0015554110370470733, -0.0023854335047460932, 
    -0.0031680363280903604, -0.0038836726531870005, -0.0045140329004647716, 
    -0.0050438906312981775, -0.0054628135654897977, -0.0057664589692508813, 
    -0.0059573147784869347, -0.0060447029508243844, -0.0060440925581587042, 
    -0.0059757201044343417, -0.0058626911980785307, -0.0057287753863719173, 
    -0.0055960446287828397, -0.0054827262306750852, -0.0054014936176536481, 
    -0.0053583021315215329, -0.0053518749898345055, -0.005373856523158544, 
    -0.0054097849811763519, -0.0054408707713040584, -0.0054465041310663292, 
    -0.0054069977644947533, -0.0053060366574631179, -0.0051324527087913416, 
    -0.0048813348835282464, -0.0045543876164404759, -0.0041596867187115739, 
    -0.0037107289081234236, -0.0032249122763053461, -0.0027214484003097259, 
    -0.0022192016639827799, -0.001734766931124546, -0.0012811910255260169, 
    -0.00086744104697856236, -0.00049856569649103257, 
    -0.00017627347374650235, 0.00010035040977545174, 0.00033431631145316732, 
    0.00053034025585316897, 0.00069455885954234112, 0.00083427805341066406, 
    0.00095754155266570423, 0.0010725310910230765, 0.0011868579404384172, 
    0.0013067346851674481, 0.0014363161328067799, 0.0015771259402489739, 
    0.0017277806226944788, 0.0018841264346367336, 0.002039806151531964, 
    0.0021871984706038259, 0.0023185875413852101, 0.0024273873138047864, 
    0.0025092339432409329, 0.002562641213240506, 0.0025892216774268235, 
    0.0025933820156974772, 0.0025816248040821102, 0.0025615311921657305, 
    0.0025405290250747133, 0.0025247184644896607, 0.0025177522323952851, 
    0.0025200996439559511, 0.0025286446007835874, 0.0025367859251723742, 
    0.002535118236668106, 0.0025124904478157368, 0.0024573853746493765, 
    0.0023592813852858206, 0.0022099418541494066, 0.0020043239170844602, 
    0.0017411398077309625, 0.0014229651783449117, 0.0010560297560637351, 
    0.00064970940196405107, 0.00021588381480610187, -0.00023176517972144203, 
    -0.0006784222862432159, -0.0011088126794146251, -0.0015078559658832122, 
    -0.0018613163140389082, -0.002156498991534945, -0.0023827750958896844, 
    -0.0025320832013254061, -0.0025991987082089143, -0.0025818193793552932, 
    -0.0024805221000626545, -0.0022985785763202865, -0.002041704031178559, 
    -0.0017176391902449955, -0.0013356910428602225, -0.00090615002251430616, 
    -0.00043962443079839799, 5.3604397304883177e-05, 0.00056419686151264127, 
    0.0010842403914975655, 0.0016076062791451481, 0.0021301598755997602, 
    0.002649767509562171, 0.0031662399863138795, 0.0036810249744504524, 
    0.0041967706644842426, 0.0047166898901494225, 0.0052437840374849731, 
    0.0057799712600440827, 0.006325195178131203, 0.0068765962849716552, 
    0.0074279273290758481, 0.0079694720576030872, 0.008488509591171256, 
    0.0089703756722528064, 0.0093999652392235018, 0.0097632485439331194, 
    0.010048731664535954, 0.010248417941227037, 0.01035832130531829, 
    0.010378531956642512, 0.010313072617317396, 0.010169564166729313, 
    0.0099588646994737181, 0.0096946007034280964, 0.0093925538804212096, 
    0.0090697685222573751, 0.0087435214613368773, 0.0084301888415272332, 
    0.0081440931183173245, 0.0078965595808758136, 0.0076952459044940733, 
    0.0075437602529714945, 0.00744156084852215, 0.0073843124810357612, 
    0.0073644504406076804, 0.0073719387752778451, 0.0073951501566018422, 
    0.0074216250308145803, 0.0074388595960385067, 0.0074348980668540064, 
    0.0073988062543570935, 0.0073210904567336584, 0.0071939401396311116, 
    0.0070113753933435004, 0.0067692172179795425, 0.0064650598472599597, 
    0.0060983537841648268, 0.0056706983794465784, 0.005186394635912547, 
    0.0046530929183450486, 0.0040821643126709699, 0.0034884926260221518, 
    0.002889336578817439, 0.0023023027523941661, 0.0017427683004869292, 
    0.0012214810757044106, 0.00074289123728568608, 0.00030480746467476225, 
    -0.00010076096138522369, -0.00048581657309889714, -0.000864034432304634, 
    -0.0012482669192920893, -0.0016480709045781825, -0.0020677761674814227, 
    -0.0025051702791258632, -0.0029512950821341407, -0.0033913320860808728, 
    -0.0038064721533939035, -0.0041763385786298254, -0.0044815099933075767, 
    -0.0047055414306401509, -0.004836258622080758, -0.0048661434932194391, 
    -0.0047919593107630162, -0.0046139834706684854, -0.0043349300073557391, 
    -0.0039592305578870692, -0.0034924297421315203, -0.0029410968626742409, 
    -0.002313199476299994, -0.0016186909942348714, -0.0008701464776913121, 
    -8.3203999285579695e-05, 0.00072344170974631078, 0.0015287846494624452, 
    0.0023108000352810893, 0.0030482216921158072, 0.0037225246672411469, 
    0.0043197600974076902, 0.004831914720082417, 0.005257590752046102, 
    0.0056018747374247009, 0.0058752875981685892, 0.0060921751482777443, 
    0.0062684537185959174, 0.0064192532458463292, 0.0065568084042365573, 
    0.0066889557207340201, 0.0068184518346864932, 0.0069432126578091559, 
    0.007057383209499609, 0.0071530714101475101, 0.0072221769640849432, 
    0.0072579843606209171, 0.0072560392031130166, 0.0072140615427462055, 
    0.0071310106069094499, 0.0070058807288048549, 0.006836719754120031, 
    0.0066203827203306408, 0.0063529685426289223, 0.0060309372643387324, 
    0.0056521277094320451, 0.0052167222716941108, 0.0047278203132321579, 
    0.0041917834998625742, 0.0036182765139416697, 0.0030199400133774854, 
    0.0024116353746061279, 0.0018094134803394997, 0.0012293682727041117, 
    0.00068657670226662045, 0.00019436052052367573, -0.00023600684236314915, 
    -0.00059528539373057449, -0.0008760674514394092, -0.001072325921391602, 
    -0.0011790476871938887, -0.0011919761513723088, -0.0011073518948725276, 
    -0.00092201449840372852, -0.00063330599294659042, 
    -0.00023899083382072537, 0.00026293159962163766, 0.00087414930296160769, 
    0.0015953076992642329, 0.0024247998445129123, 0.0033567970136302492, 
    0.0043793013149468303, 0.0054727227991697922, 0.0066093060421021522, 
    0.0077533235824919187, 0.0088625292719712225, 0.0098900661913959576, 
    0.010786941972467042, 0.011505047680696641, 0.012000798828127773, 
    0.012238801228702242, 0.012195905927244375, 0.01186475564074636, 
    0.011256395424837012, 0.01040106477585068, 0.0093467674798353977, 
    0.0081556067049400882, 0.0068982928332925837, 0.0056477278013616853, 
    0.0044729782411666906, 0.0034343629012012211, 0.0025807287182549065, 
    0.0019485553963085357, 0.0015627989328158304, 0.0014386465867646209, 
    0.0015835846620598578, 0.0019991495415915038, 0.0026819340294479094, 
    0.0036231068231912509, 0.0048066963802159517, 0.0062068856474747037, 
    0.0077856568236537166, 0.009492370424343647, 0.01126650103998493, 
    0.013042999404732554, 0.014758910468444363, 0.016359273377124069, 
    0.017800932751599399, 0.019053357783951577, 0.02009657747732542, 
    0.020917005710701816, 0.021501995563683322, 0.021835182763768543, 
    0.021893738038999657, 0.021649090172139191, 0.021071664294351096, 
    0.020138521681106893, 0.018841429694195066, 0.017192443498935967, 
    0.015224466556432243, 0.012987067550608364, 0.010538977935231099, 
    0.0079407419966116451, 0.0052490259327010874, 0.0025141632855024401, 
    -0.00021969086221250303, -0.0029119864744555865, -0.0055236562997533906, 
    -0.0080152170581571768, -0.010347940995935851, -0.012486858149555925, 
    -0.01440659709459245, -0.016097298987762399, -0.01756770445007513, 
    -0.018843064273219971, -0.019956271049674075, -0.020936314815587852, 
    -0.021798434731904331, -0.022539570481072795, -0.023139668703859216, 
    -0.023566573989704142, -0.023782015514595051, -0.023747006856519343, 
    -0.023424851064161541, -0.022784442231859235, -0.021803484564848694, 
    -0.020473093536831587, -0.018803147816235787, -0.016827240393992155, 
    -0.014605520830518772, -0.012221360462140516, -0.0097743015734581724, 
    -0.0073668526612160768, -0.0050910055274819496, -0.0030159577140190397, 
    -0.0011811145528957527, 0.00040689508985898917, 0.0017726392253173975, 
    0.0029664052318488713,
  // Fqt-F(9, 0-1999)
    1, 0.98893242323054786, 0.95654649626830779, 0.90518486840591794, 
    0.83840625841353089, 0.76053732734872936, 0.67617215782278217, 
    0.5897045462402597, 0.50495955355189759, 0.42496077174530078, 
    0.35183810885683181, 0.286855561658862, 0.23052381639150124, 
    0.18275875601141331, 0.14305184470531154, 0.11062784053642744, 
    0.084575827775116394, 0.063948753773166278, 0.047832722063701462, 
    0.035390713208733299, 0.025886477557880257, 0.018693865710151865, 
    0.013295979400047042, 0.0092774652108557985, 0.0063124774614186467, 
    0.0041503713295463875, 0.0026007640370849629, 0.0015194081748312466, 
    0.00079591356195117177, 0.00034394959802728071, 9.4140660228180317e-05, 
    -1.0597999730973279e-05, -1.7763223281116821e-05, 3.3369016889773419e-05, 
    0.00011114585588517178, 0.00019126358766605379, 0.00025654103331819618, 
    0.00029658646412719669, 0.00030731624745847821, 0.00029029547856186715, 
    0.00025189000881910197, 0.0002021983564615055, 0.00015375124446030295, 
    0.00011998256407912486, 0.0001134912018754446, 0.00014426105046372355, 
    0.00021803295017921811, 0.00033514131898175931, 0.0004900612981449256, 
    0.00067180342716395504, 0.00086511338150077122, 0.0010523213241013737, 
    0.0012155335556392351, 0.0013388372527067605, 0.001410166286348304, 
    0.0014225648113844755, 0.0013746706840282951, 0.001270394824430716, 
    0.0011179409359016908, 0.00092835853402457771, 0.00071391162118351523, 
    0.00048652003381922265, 0.00025650988574602734, 3.1818085593003902e-05, 
    -0.00018224852691419395, -0.00038273682697327301, 
    -0.00056835724635373539, -0.0007385957023936068, -0.00089283886308728021, 
    -0.0010297301153225809, -0.0011468943263948728, -0.0012410473037059923, 
    -0.001308447791102414, -0.0013455370244662074, -0.001349623438736547, 
    -0.0013194527210985188, -0.0012555660617370194, -0.0011604181015385385, 
    -0.0010382450968035436, -0.00089474184589527007, -0.00073662005191261766, 
    -0.00057113565707566478, -0.00040566785517900125, 
    -0.00024738431406170927, -0.00010299873700874679, 2.142016371327267e-05, 
    0.00012066289269128987, 0.0001906360051101244, 0.00022870555173834707, 
    0.0002340517021204, 0.00020798388763526701, 0.00015407290448478074, 
    7.8048055221897146e-05, -1.2622863613943273e-05, -0.00010941787902534947, 
    -0.00020365557029021036, -0.00028741592428638545, 
    -0.00035438915307991461, -0.00040051408569149506, 
    -0.00042432222968657172, -0.00042698501651631984, 
    -0.00041203141661943523, -0.0003848067642933387, -0.00035173613698454064, 
    -0.00031950054701203025, -0.00029425603208261771, -0.0002810066477791929, 
    -0.00028321454349993403, -0.00030267759907859132, 
    -0.00033967368899416611, -0.00039328391912390364, 
    -0.00046180488579774815, -0.00054313113803647621, 
    -0.00063501912801329562, -0.00073516433135391399, 
    -0.00084108515509113307, -0.00094987257815439745, -0.0010578757932854803, 
    -0.0011604650969985189, -0.0012519693602794056, -0.0013258780275075749, 
    -0.0013753184045253051, -0.0013937665097467917, -0.0013758792145752174, 
    -0.0013183305403478927, -0.0012205096105323894, -0.001084990554148889, 
    -0.00091769171877871525, -0.00072769918745306029, 
    -0.00052673856850712485, -0.0003283398210218933, -0.00014678815546673526, 
    4.0516440087258834e-06, 0.00011188625291497217, 0.00016700251082748261, 
    0.00016303429002488247, 9.7404506977215923e-05, -2.8580039533189264e-05, 
    -0.00020995059591758953, -0.00043856031181244983, 
    -0.00070373878826538133, -0.00099302258843989347, -0.0012928967601798114, 
    -0.0015894745095528793, -0.0018691015266182019, -0.0021188466566239251, 
    -0.0023269351231795729, -0.00248313634921576, -0.0025791448450720399, 
    -0.0026089694229634161, -0.0025693119848441189, -0.0024598720778885043, 
    -0.0022835008993393482, -0.0020461520676363608, -0.0017565809588871101, 
    -0.0014258295927382298, -0.0010665111396537157, -0.0006920135023846507, 
    -0.00031567966581418896, 4.9936823471148195e-05, 0.00039371343522525256, 
    0.00070645285382601455, 0.00098126287867960553, 0.0012138026666861452, 
    0.0014023835564982868, 0.0015479241807418336, 0.0016536791307481468, 
    0.0017247220140305128, 0.0017671461558138436, 0.0017870609723700489, 
    0.001789501486205638, 0.0017774467574405155, 0.001751110594554068, 
    0.0017076930005108641, 0.0016416876187261994, 0.0015457035241925607, 
    0.0014116576514275046, 0.0012320535106446664, 0.0010011379970614671, 
    0.00071572740045800008, 0.00037565204026677047, -1.6152425003460529e-05, 
    -0.00045382098373275461, -0.00092890197759566326, -0.0014307932152131041, 
    -0.0019471916711095785, -0.002464580293481281, -0.0029687187623257906, 
    -0.0034451799902558136, -0.0038799362409801131, -0.0042600034240851143, 
    -0.0045740949315130645, -0.0048132859534555025, -0.0049715857465655721, 
    -0.0050463987303317652, -0.0050387839723940314, -0.0049534706596578775, 
    -0.0047986014253016632, -0.0045851834480451596, -0.0043262795401007434, 
    -0.0040360288115492814, -0.0037286104702424269, -0.0034172744926144684, 
    -0.0031135673713238651, -0.0028268116349064172, -0.0025639103123319558, 
    -0.0023294573907709937, -0.0021261061705674027, -0.0019550884377643996, 
    -0.0018167908090414957, -0.0017112532369451862, -0.001638516786041766, 
    -0.0015987499846768125, -0.0015921430511340086, -0.0016185824655022705, 
    -0.0016771477543640698, -0.0017655314632115679, -0.0018795015466440122, 
    -0.0020125435945946317, -0.0021558096249093958, -0.0022984757141284967, 
    -0.0024284813352043284, -0.0025335962572700503, -0.0026026434858439631, 
    -0.0026267080288727138, -0.0026001315412863091, -0.0025211681388737322, 
    -0.0023922123331039883, -0.0022196103896907965, -0.0020131045987498292, 
    -0.00178500761077011, -0.0015492361593066261, -0.0013202820334942407, 
    -0.0011121894389261742, -0.00093758295441360984, -0.00080678707210724064, 
    -0.00072707748864567396, -0.00070210423767691173, 
    -0.00073155579335348843, -0.00081110270205340799, -0.0009326849774525304, 
    -0.0010851370625516211, -0.0012551294231784606, -0.0014283302972826486, 
    -0.0015906577132292108, -0.0017295091403150531, -0.0018348376146749587, 
    -0.0019000113191301776, -0.0019223785931482323, -0.0019035335882153571, 
    -0.0018492156213552574, -0.0017688322183225386, -0.0016745871255927204, 
    -0.0015802635849813003, -0.0014997302238305347, -0.001445350140140769, 
    -0.0014264549022536383, -0.0014481046678020914, -0.0015103111042684937, 
    -0.0016078589896108258, -0.001730767723898696, -0.0018653457760658613, 
    -0.0019957231731836376, -0.0021056421264345265, -0.0021802588579122439, 
    -0.0022077342920024268, -0.0021803895063842813, -0.0020953329364577842, 
    -0.0019545603472291744, -0.0017645901770334958, -0.0015357530749765635, 
    -0.0012812625975781302, -0.0010161519102502722, -0.00075614939471594842, 
    -0.00051652527805152028, -0.00031094573326801816, 
    -0.00015037887811169236, -4.2110896870231133e-05, 1.1015404208582528e-05, 
    1.1030314319616309e-05, -3.5202887865607769e-05, -0.00011658182341080678, 
    -0.00021893633185740528, -0.00032669431680198741, 
    -0.00042485283040295785, -0.00050098976184349755, 
    -0.00054696073164779094, -0.00055999304538832423, 
    -0.00054292779509312503, -0.00050353366943169922, 
    -0.00045297475774660215, -0.00040372958558063181, 
    -0.00036736349783797896, -0.00035263532371689955, 
    -0.00036434115647871889, -0.00040312501314669147, 
    -0.00046625380298583459, -0.0005490917309223072, -0.00064681449442820162, 
    -0.00075585899552821963, -0.00087470098796752676, -0.0010037626409448812, 
    -0.0011445462176410412, -0.0012983330143965027, -0.0014649126437466704, 
    -0.0016417874081083356, -0.0018240788308710463, -0.0020051653409088903, 
    -0.0021777569374102084, -0.0023350632247673636, -0.0024716760650963518, 
    -0.0025839416598196384, -0.0026698346088481757, -0.0027284904930486059, 
    -0.0027596554727156285, -0.0027632688644103711, -0.0027392589111871943, 
    -0.0026875331278004224, -0.0026080314640591486, -0.0025007498943579601, 
    -0.0023656881165947312, -0.0022027526495891746, -0.002011705464196351, 
    -0.0017922433562235049, -0.0015442609590893431, -0.001268301394454235, 
    -0.00096612498521430452, -0.00064130543624168319, 
    -0.00029970822435228749, 5.0264360036504467e-05, 0.00039778666833084749, 
    0.00073015614639173492, 0.0010338007085315172, 0.0012956473691601879, 
    0.0015047077318446353, 0.0016536229068723376, 0.0017398882461227745, 
    0.0017665263649069797, 0.0017419841192301572, 0.0016792548643958887, 
    0.0015943104690042131, 0.0015041010769948728, 0.001424460494919308, 
    0.0013682651353009801, 0.0013441415481213407, 0.0013559152030570253, 
    0.0014028223448757399, 0.0014803900809062685, 0.0015817399089643263, 
    0.0016990300847985822, 0.001824701568504866, 0.001952310316232221, 
    0.0020768015925530623, 0.0021942972922171346, 0.0023015447342882465, 
    0.002395269605121477, 0.0024716320213997302, 0.0025259205224974035, 
    0.0025525876610413825, 0.0025456497486135909, 0.0024994005144930429, 
    0.0024092686542096097, 0.0022726575329851256, 0.0020895406690672994, 
    0.0018627661407860947, 0.0015980068146174715, 0.0013034481685634672, 
    0.00098925956809514464, 0.00066694554648977005, 0.0003486241852268321, 
    4.6288615927573905e-05, -0.00022892141347206774, -0.00046740671835465171, 
    -0.00066172508118789457, -0.00080711410873487044, 
    -0.00090186582231103118, -0.00094753210482703253, 
    -0.00094890208802342042, -0.00091369222438929644, 
    -0.00085192614987765003, -0.00077500588834279716, 
    -0.00069454251003134922, -0.00062111326536679783, 
    -0.00056308110580593628, -0.00052566201012647223, 
    -0.00051035112735016549, -0.00051480033841444549, 
    -0.00053317542543700538, -0.0005569724163478571, -0.00057620459861467441, 
    -0.00058082458864016902, -0.00056215949824144529, -0.0005141644114562366, 
    -0.0004343295072468712, -0.00032421359843636893, -0.00018956904696942241, 
    -4.0127000325868487e-05, 0.00011099584772823255, 0.00024822727934612832, 
    0.00035482219856815457, 0.00041442817127923439, 0.00041279707861228759, 
    0.00033951215824814428, 0.00018947043944053009, -3.6060086355266854e-05, 
    -0.00032901848609274834, -0.00067487002452985205, -0.0010536785521119713, 
    -0.0014418329643035319, -0.0018142324317394808, -0.0021466696626491798, 
    -0.0024180866190735241, -0.002612446271854022, -0.002719987541066921, 
    -0.0027377191434410477, -0.0026691764614324522, -0.0025235044359129943, 
    -0.0023141026482076509, -0.0020570191274979555, -0.0017693173861675034, 
    -0.0014675811368391189, -0.0011666712004036277, -0.0008788569600235753, 
    -0.00061334013230908695, -0.00037617440400978587, 
    -0.00017049877571999835, 3.0515307607703579e-06, 0.00014585802007251533, 
    0.00026085278384761464, 0.00035211750400886035, 0.00042451617647882743, 
    0.0004833100299718331, 0.00053371019279462625, 0.00058034104392740951, 
    0.00062668580614259309, 0.00067462791530073225, 0.0007241715963281324, 
    0.00077345120165765952, 0.00081902241098987373, 0.00085640618032579324, 
    0.00088077673549321104, 0.00088770928747014879, 0.00087383244315483288, 
    0.00083729485005324766, 0.00077794379684122832, 0.0006972028598261125, 
    0.00059774471336798631, 0.00048306395455927179, 0.00035704056312121799, 
    0.00022354182571324795, 8.607103252229601e-05, -5.2499884647665357e-05, 
    -0.00019005745916449634, -0.00032519514608268395, -0.0004569981236030022, 
    -0.00058468990094191862, -0.00070724090598307874, 
    -0.00082303411443663123, -0.00092968160099460816, -0.0010240775366515964, 
    -0.00110271558015601, -0.0011622339706592781, -0.0012000736722586932, 
    -0.001215102995354693, -0.0012080526399389628, -0.0011816298889078996, 
    -0.0011402779612743631, -0.0010895831852475528, -0.0010354652049902188, 
    -0.00098329847322908967, -0.00093713647988840872, 
    -0.00089918408039765362, -0.00086962187842782343, 
    -0.00084681442178308121, -0.0008278264186190017, -0.0008091342213301418, 
    -0.00078733032806384317, -0.00075965478559108233, 
    -0.00072420534472270634, -0.00067980461734946083, 
    -0.00062561587049020861, -0.00056064506301315559, 
    -0.00048336147868465395, -0.00039158610567906899, 
    -0.00028273959601481731, -0.00015445151917759084, 
    -5.4078045364601554e-06, 0.00016376757535251606, 0.00034983307274349848, 
    0.00054663180745195741, 0.00074534289929153129, 0.0009352836474414277, 
    0.0011051338384706216, 0.0012443761766107063, 0.0013446948601051111, 
    0.001401072924979801, 0.001412413607859179, 0.0013816168228281119, 
    0.0013151197175467143, 0.0012220396170486425, 0.0011130776529000058, 
    0.00099940672377311435, 0.0008916491970481135, 0.00079910273515147419, 
    0.0007292220755932353, 0.00068738813851301653, 0.00067692369770212747, 
    0.00069930178471017221, 0.00075448419050325058, 0.00084130650177984901, 
    0.00095782578524882033, 0.0011015745630790327, 0.0012696715220504469, 
    0.0014587875719329379, 0.0016650162482769429, 0.0018837073811416635, 
    0.0021093405750289246, 0.0023355108462550511, 0.0025551050578622851, 
    0.0027606530328628115, 0.0029448376335907871, 0.0031010555890690255, 
    0.0032239565941921235, 0.0033098798019367912, 0.0033571259881588836, 
    0.0033660542777105324, 0.0033389971200603226, 0.003279964297673489, 
    0.0031941306224871849, 0.0030871314904680272, 0.002964308320437317, 
    0.0028300167493103463, 0.0026871755878098516, 0.0025370858271958306, 
    0.0023795687524123445, 0.0022133542444705517, 0.0020366496139330665, 
    0.0018477904848022537, 0.0016458305179868949, 0.0014309669597149565, 
    0.0012047263024985303, 0.00096988755554581368, 0.00073022118206582864, 
    0.00049008048750625449, 0.00025392312359585098, 2.5773362318518136e-05, 
    -0.00019132201849963177, -0.00039580696578899724, 
    -0.00058799923964441777, -0.00077024420616419141, 
    -0.00094674751234220551, -0.0011230455029648605, -0.0013050988929104669, 
    -0.0014981398296721323, -0.0017054131511093043, -0.0019270798229648533, 
    -0.0021594995481647116, -0.0023950592633383509, -0.0026226172274620963, 
    -0.0028285212435525489, -0.002998022997286862, -0.0031168932453983994, 
    -0.0031730229599587576, -0.0031578049821742202, -0.0030671037718644624, 
    -0.0029016591498411946, -0.0026668865569336366, -0.0023721508214042293, 
    -0.0020296622060402402, -0.0016532468773334224, -0.0012571763948858459, 
    -0.00085521871522446303, -0.0004599836282980635, -8.2550428914918801e-05, 
    0.00026768599757899037, 0.00058302363876337846, 0.00085740913501162108, 
    0.0010864154123226609, 0.0012672489156487702, 0.001398769305384016, 
    0.0014814886774613002, 0.0015174976197868798, 0.0015102813735606681, 
    0.0014644196650423634, 0.0013851668043905804, 0.0012780043269110726, 
    0.0011482103094054099, 0.0010005373857866449, 0.00083901738744388823, 
    0.00066692914934850028, 0.00048686223692985563, 0.00030086786347892705, 
    0.00011067234868143998, -8.2082561550758507e-05, -0.00027559759094668475, 
    -0.00046771211041670465, -0.0006557598686963848, -0.00083649224854247478, 
    -0.0010060787910920162, -0.001160136875445424, -0.0012938496215347739, 
    -0.0014021446010867591, -0.0014799865599013618, -0.001522779281904254, 
    -0.0015268934137430369, -0.0014902393283014188, -0.0014128013526519927, 
    -0.0012970001144952314, -0.0011477161792613319, -0.00097192499328542362, 
    -0.00077795656796205456, -0.00057451492381426546, 
    -0.00036969515404709937, -0.00017020589929454919, 1.9015876435511127e-05, 
    0.0001947744580635439, 0.00035524369487578499, 0.00049940975481712474, 
    0.00062652585929559123, 0.00073571515269570597, 0.00082579500323252389, 
    0.00089532014072105266, 0.00094278117111490736, 0.00096689102928265312, 
    0.00096685177308318223, 0.00094256394236276041, 0.00089471082602904871, 
    0.00082470376807373827, 0.00073450690496259564, 0.00062642961957075079, 
    0.00050295419792307453, 0.00036667645007715244, 0.00022039501085017961, 
    6.7297734554947348e-05, -8.8823381708339646e-05, -0.00024341163211436768, 
    -0.0003910980298490078, -0.0005258260874899123, -0.00064114843558886047, 
    -0.00073066151229254504, -0.00078854358103789158, 
    -0.00081008849407655022, -0.00079216347265234491, 
    -0.00073354161892131588, -0.0006350620008157325, -0.00049960278312623186, 
    -0.00033185864107790548, -0.00013795654836090817, 7.5025695897754942e-05, 
    0.00029956186305843516, 0.0005281128137435868, 0.00075340937741369429, 
    0.00096854233706681627, 0.0011668634806827416, 0.0013417427151487921, 
    0.0014862834501803465, 0.0015931266519897008, 0.0016544788508277776, 
    0.0016624423373965184, 0.0016096451822235054, 0.0014901506239767184, 
    0.0013005161230918148, 0.0010408327358791423, 0.00071555741319861087, 
    0.00033391317199461942, -9.0280716903154716e-05, -0.00053942751410489048, 
    -0.00099353915517354707, -0.0014319815040899271, -0.0018353145732004645, 
    -0.0021869174129150863, -0.0024741886586735181, -0.0026892078401330793, 
    -0.0028288422863373564, -0.0028943854028820261, -0.002890791730760059, 
    -0.0028257110254734387, -0.002708432492601586, -0.0025488716253943308, 
    -0.002356693146701133, -0.0021406404507959016, -0.0019080816906518023, 
    -0.0016647850748487982, -0.0014148915956771462, -0.0011610268529269909, 
    -0.0009045531512078351, -0.00064591578574926876, -0.00038511528830035061, 
    -0.00012225683906037766, 0.00014185376536225724, 0.00040519637282375855, 
    0.00066425318939416882, 0.00091401975126790744, 0.0011482632501619557, 
    0.0013598922293400675, 0.0015413166104069156, 0.0016847459324868573, 
    0.0017824696787121, 0.0018271806223537934, 0.0018124015149923092, 
    0.0017330465327825817, 0.0015860846332147948, 0.001371256640574043, 
    0.001091700393308043, 0.00075430915559416569, 0.000369656138976091, 
    -4.8609122017758332e-05, -0.00048485554599052657, 
    -0.00092290798973104771, -0.0013475642714645892, -0.001745945133849383, 
    -0.0021084742220481602, -0.0024293085217979987, -0.0027062118731910551, 
    -0.0029398985606257913, -0.003133017020193377, -0.0032889804478220424, 
    -0.0034108941262561347, -0.0035008157667830307, -0.0035594822054657222, 
    -0.0035865804692920356, -0.0035814704885460034, -0.0035441830729183547, 
    -0.0034764523559346018, -0.0033825005783595045, -0.0032693561037984535, 
    -0.0031465974402078321, -0.0030255193213416642, -0.0029178787634922066, 
    -0.0028344559108800828, -0.0027837196911711906, -0.0027708575408348511, 
    -0.0027973364299824729, -0.0028609979878743193, -0.0029566116814840624, 
    -0.0030766981651971208, -0.0032124274694454967, -0.0033544395086221191, 
    -0.0034934852363947256, -0.0036208731698574893, -0.0037287220839782561, 
    -0.0038100834411324536, -0.0038589819968947912, -0.0038704328281666308, 
    -0.0038405286648235623, -0.0037666584870160412, -0.0036478569963089512, 
    -0.0034852022331755546, -0.0032820840089092368, -0.0030441453746030815, 
    -0.0027787595065959011, -0.0024940300281628669, -0.0021975023278062158, 
    -0.0018948135636591569, -0.0015886505454093482, -0.0012782525417800443, 
    -0.00095962947649446957, -0.00062647397204428372, 
    -0.00027164862749512627, 0.00011105990781584951, 0.00052521143928579061, 
    0.00097036765046564497, 0.001441395675229204, 0.0019285650339746225, 
    0.0024184009199370859, 0.0028950764642936195, 0.0033420436434968186, 
    0.0037435950212348222, 0.0040861115684918065, 0.004358885948979061, 
    0.0045545205918948927, 0.0046690104752111217, 0.0047016249975904536, 
    0.0046547483855953848, 0.0045337540842179799, 0.0043469145680001845, 
    0.0041052905655784861, 0.0038224700449965275, 0.0035140349884648443, 
    0.0031966990737470123, 0.0028871377288314758, 0.0026006719138698502, 
    0.0023500066373250616, 0.002144268788301294, 0.001988513121541018, 
    0.001883751289595991, 0.0018274654463927898, 0.0018144208897387928, 
    0.0018376120558271959, 0.0018891304004153889, 0.0019608521297972401, 
    0.0020449002418012137, 0.0021339176421427642, 0.0022212517029530573, 
    0.0023010999854519614, 0.0023686791243673513, 0.0024204081947731635, 
    0.0024540197550813724, 0.0024685449219185181, 0.0024640978010590522, 
    0.0024415006879630308, 0.0024018249860742807, 0.0023459748783184469, 
    0.0022744666383846695, 0.0021874506615064291, 0.0020849598221655366, 
    0.0019673133187971671, 0.0018355321942941565, 0.0016916477836870041, 
    0.0015388330835420841, 0.0013813069455474456, 0.0012240143285809396, 
    0.0010721362910639308, 0.00093051010503963937, 0.00080306281022354462, 
    0.00069233557779619888, 0.00059922802683285835, 0.0005229651668329857, 
    0.00046129708711153267, 0.00041089880171251325, 0.00036788630131696855, 
    0.00032836315021252756, 0.00028891491816640134, 0.00024697028779587296, 
    0.00020096853491068711, 0.00015029053379446208, 9.4957287924930445e-05, 
    3.5162521398591071e-05, -2.9272522125521204e-05, -9.9400769763107128e-05, 
    -0.00017747238432217892, -0.0002670179412154698, -0.0003726450737740941, 
    -0.00049962324313216721, -0.00065328413828582882, 
    -0.00083833591668398388, -0.0010581623129400331, -0.001314151547204261, 
    -0.0016051039678595452, -0.0019267971281010355, -0.0022718267618796451, 
    -0.0026298587515828061, -0.0029883357421827462, -0.0033336359623734181, 
    -0.0036525276800079241, -0.003933689105089077, -0.004169071147277055, 
    -0.0043548577268156625, -0.0044918722553977872, -0.0045853346126273108, 
    -0.0046439627148216686, -0.0046785490904451693, -0.0047002001310608868, 
    -0.0047185168782058395, -0.0047400241954244837, -0.0047670941702791427, 
    -0.0047975229859364612, -0.0048248350133108598, -0.0048392051515645318, 
    -0.0048288407616312208, -0.0047815544787564689, -0.0046862879281533362, 
    -0.0045343433267678061, -0.004320190114853387, -0.0040417659465011345, 
    -0.003700338411891331, -0.0033000063720639893, -0.0028470095072133973, 
    -0.0023490306766521724, -0.0018146300998737601, -0.0012528742137121944, 
    -0.0006731681906060286, -8.5247463589858009e-05, 0.00050079018851764234, 
    0.0010744898822518116, 0.0016251716237235718, 0.0021422469707564834, 
    0.0026156985617673215, 0.0030366414910964522, 0.0033978716101857173, 
    0.0036943098607146027, 0.0039233396808433102, 0.0040850053399920077, 
    0.0041820946446115143, 0.0042200369923118429, 0.00420660517505295, 
    0.0041513860041104333, 0.0040650230828515356, 0.0039583137611498703, 
    0.0038412622069115368, 0.0037221667512177363, 0.003606891038813567, 
    0.0034983425368093637, 0.0033962413883658793, 0.00329713124670646, 
    0.0031946762978645933, 0.0030802279105622554, 0.0029436831457484423, 
    0.0027745999887912941, 0.0025634744510512632, 0.0023030536106718059, 
    0.0019894618889216187, 0.0016229618613326656, 0.0012081992831800004, 
    0.00075388573384929799, 0.00027197178723882521, -0.00022357159516287476, 
    -0.00071816596269591842, -0.0011980109481608365, -0.0016511937889560095, 
    -0.0020683617928549097, -0.0024428440726835992, -0.0027702733886874509, 
    -0.0030478565894391327, -0.0032735666699223714, -0.003445506388775737, 
    -0.0035616427876344046, -0.0036199595992656586, -0.0036189455099343896, 
    -0.0035582771105476174, -0.003439453157306501, -0.0032661708898035794, 
    -0.003044292401481883, -0.0027813671339983353, -0.0024858483325492179, 
    -0.0021662838898901162, -0.0018307672151881855, -0.0014868379692527375, 
    -0.0011418477500879836, -0.00080356002585094414, -0.0004806664128750868, 
    -0.00018285523392703735, 7.9724389675307251e-05, 0.0002976155298379129, 
    0.00046353885572551225, 0.00057387828390743651, 0.00062970786403299377, 
    0.00063708388341825986, 0.00060642298115411999, 0.00055107848301664609, 
    0.00048541818685640735, 0.00042276871344796668, 0.00037366474383288527, 
    0.00034469308334273888, 0.0003380782005354214, 0.0003520358822586695, 
    0.00038171101829700033, 0.0004205052981145503, 0.00046151388059721801, 
    0.00049881073347407068, 0.00052834867366180049, 0.00054830950619534787, 
    0.00055891483992432333, 0.0005618249027988301, 0.00055934633809760943, 
    0.00055369340244773308, 0.00054641740386213698, 0.00053807895939593574, 
    0.00052812770179466143, 0.00051494402834628716, 0.00049602810746466317, 
    0.00046827488527640608, 0.00042833118406884594, 0.0003730299248291289, 
    0.00029988778754359738, 0.00020764079463073254, 9.6751962028737769e-05, 
    -3.0205626745405032e-05, -0.00016840610525799786, 
    -0.00031092116704969409, -0.00044915063914112273, 
    -0.00057342544845591793, -0.00067369987136831197, 
    -0.00074025521309400489, -0.00076435671296582971, 
    -0.00073886225739127807, -0.00065877990830732959, 
    -0.00052172960357166158, -0.00032822975557737376, 
    -8.1766723362828285e-05, 0.00021139839780926921, 0.00054265147897691532, 
    0.00090158765354133512, 0.0012765854300509137, 0.001655253840002561, 
    0.0020247202768190454, 0.0023717876698479976, 0.0026831602005442266, 
    0.0029458772446926702, 0.0031480933962505105, 0.0032801824560300626, 
    0.0033359815471225344, 0.0033139791852206234, 0.0032181542378995898, 
    0.003058180860119985, 0.0028488300104661749, 0.0026085118281159851, 
    0.002357155264308275, 0.0021137337877698719, 0.0018938482390459918, 
    0.0017077562159579021, 0.0015591576759360552, 0.00144494329816808, 
    0.0013559991678671487, 0.0012789595875648974, 0.0011986729952416695, 
    0.001100964344209555, 0.00097521029468724445, 0.00081624440477827995, 
    0.00062530645846596154, 0.00040992368607650233, 0.00018282780105983434, 
    -3.9854042204801884e-05, -0.00024081854333251687, 
    -0.00040391396240950202, -0.00051630133474647451, 
    -0.00057017930564892553, -0.00056378564294356213, 
    -0.00050149297692590809, -0.00039296364333677315, -0.0002515346802721886, 
    -9.2175305679471377e-05, 7.052543012323032e-05, 0.00022403312348558677, 
    0.00035896090193760633, 0.0004695596342653845, 0.00055367114049678667, 
    0.00061225363342543471, 0.00064863493874670834, 0.00066765468185179004, 
    0.00067484888722967257, 0.00067578767592697602, 0.00067566852745613816, 
    0.00067919206583903974, 0.00069067095106352351, 0.00071428354255177772, 
    0.00075437097944184943, 0.0008156153919860621, 0.0009030185198187976, 
    0.0010215695793396767, 0.0011756869568000615, 0.0013685130659383843, 
    0.0016012350652899014, 0.0018725856743158195, 0.002178567771668821, 
    0.0025124345245038709, 0.0028648726014039766, 0.0032243788123788222, 
    0.0035778399723049321, 0.0039113048926075721, 0.0042108611597546928, 
    0.0044635248706449407, 0.0046579693126968715, 0.0047850089748255357, 
    0.0048378512912906312, 0.0048122305468245082, 0.0047065905269412303, 
    0.0045223658659161283, 0.0042642610903456373, 0.0039403303848890769, 
    0.0035616865393073684, 0.0031417321530609809, 0.0026949770484537765, 
    0.0022356504027602518, 0.001776385205920307, 0.0013272344397993129, 
    0.0008952186487052329, 0.00048450250446839619, 9.7059843299102322e-05, 
    -0.00026638284202147486, -0.00060543127491697289, 
    -0.00091942174063423387, -0.0012072779007136338, -0.0014678174146483566, 
    -0.001700340814136765, -0.0019052301180493099, -0.0020843022761540706, 
    -0.0022407377156362122, -0.0023785472923753214, -0.0025016625668554966, 
    -0.0026128467490086713, -0.0027126805603789302, -0.0027988507816079757, 
    -0.0028659331549328016, -0.0029057155998709746, -0.0029080648858757835, 
    -0.0028621582657885579, -0.0027579017514658688, -0.0025873465845390833, 
    -0.0023458916335003838, -0.0020331795118447476, -0.0016535327872129848, 
    -0.0012158913196675355, -0.00073322834141632581, -0.00022154170098770816, 
    0.00030142923662701061, 0.0008175626453772076, 0.0013096066422851949, 
    0.0017621581609972875, 0.0021622677119803447, 0.002499695597447376, 
    0.002766881827271249, 0.0029587549402023848, 0.0030725319754754594, 
    0.003107581851328191, 0.0030654229871650137, 0.0029497680057136723, 
    0.0027666075980086278, 0.0025241409826113788, 0.0022325207990556892, 
    0.0019033367407705636, 0.001548861889263869, 0.0011811696860149457, 
    0.00081124954607488778, 0.000448304903206473, 9.9344984348285136e-05, 
    -0.00023081688775185763, -0.00053917867716000328, 
    -0.00082381718788396329, -0.0010830111048436347, -0.0013144201225734529, 
    -0.0015145354014149657, -0.0016785717010828851, -0.0018008816931367796, 
    -0.0018758436350034202, -0.0018990426602500459, -0.0018684837068325892, 
    -0.0017856026903322077, -0.0016558776616991792, -0.0014888928017472978, 
    -0.001297811835595032, -0.0010982715534231322, -0.00090686241804035746, 
    -0.00073936300048723529, -0.0006089838376225642, -0.00052484443745382013, 
    -0.00049090170941274163, -0.00050546462991057505, 
    -0.00056139704538479525, -0.00064694709771229608, -0.0007471181790423742, 
    -0.00084537489912571363, -0.00092546378622430144, 
    -0.00097309740990308004, -0.00097731794096370811, 
    -0.00093136878383621156, -0.00083302885646586165, 
    -0.00068443965567230064, -0.00049157075318033211, -0.0002634850212244303, 
    -1.1549162503264514e-05, 0.00025135780489523641, 0.00051159626839021306, 
    0.00075552570703814532, 0.0009702954918425074, 0.0011446481880776661, 
    0.0012696776774223731, 0.0013394550958900867, 0.0013513933669150819, 
    0.0013062903158415371, 0.0012080239916052397, 0.001062955813369861, 
    0.00087910142260953761, 0.00066519825294610979, 0.00042984331280921534, 
    0.00018078545127472563, -7.5457345231177324e-05, -0.00033365161070417562, 
    -0.00058960106936824881, -0.00083973030819664638, -0.0010806633891998834, 
    -0.0013089546954222089, -0.0015209907031765539, -0.0017131209034227895, 
    -0.0018819376151743097, -0.0020245824179824911, -0.0021389717182958359, 
    -0.0022238835900274413, -0.0022788828510972147, -0.002304137162881398, 
    -0.0023002085878199635, -0.0022679063425372877, -0.0022082165679987763, 
    -0.0021222623859067096, -0.0020112785143086868, -0.0018765062908240725, 
    -0.0017190585809492348, -0.0015398185440948183, -0.0013394761208554836, 
    -0.0011188157786083766, -0.00087919041467613519, -0.00062310635049415237, 
    -0.00035468556619345105, -7.9864816879285806e-05, 0.00019379747953146749, 
    0.00045765239142982905, 0.00070279860538262806, 0.00092100226892904177, 
    0.0011055720447207397, 0.0012520363418988593, 0.0013585080620447942, 
    0.0014257387430210394, 0.0014568838023343903, 0.0014571372847741139, 
    0.0014332682869422312, 0.0013931348137047298, 0.0013450899796332739, 
    0.0012972619959958982, 0.001256671724537561, 0.0012282411062653569, 
    0.0012138733292625617, 0.0012118681341925144, 0.0012169005478514286, 
    0.0012206937915341402, 0.0012133202062193193, 0.0011848723501973503, 
    0.0011271841967684672, 0.0010351762918113547, 0.00090764605559062262, 
    0.0007473398070584927, 0.00056036931308702453, 0.00035511770142525941, 
    0.00014084987383163679, -7.3750857236250114e-05, -0.00028185925843071658, 
    -0.00047936762446018828, -0.00066510888330328954, 
    -0.00084039048881068149, -0.0010079157098530148, -0.0011703430615814137, 
    -0.0013288214758380846, -0.0014818682338793418, -0.0016248275348626699, 
    -0.0017500666402558351, -0.0018478231744103301, -0.0019075803267746114, 
    -0.0019196494750732536, -0.0018767229217615132, -0.0017751119639968806, 
    -0.0016155311311731261, -0.0014033691542023204, -0.0011484282143638632, 
    -0.00086420395759573472, -0.00056684085069487553, 
    -0.00027388899429421724, -3.0152039706622978e-06, 0.00022924513686168354, 
    0.00040858717678574964, 0.00052396483184761447, 0.00056846029151067531, 
    0.0005399442841572883, 0.00044132356779021348, 0.00028018662908005506, 
    6.7756212041219903e-05, -0.00018286196012147731, -0.00045885667888856347, 
    -0.00074988567879574232, -0.0010496693489313845, -0.0013565092988686721, 
    -0.0016725732727661704, -0.0020021156726123431, -0.0023491487412066955, 
    -0.0027150818126708254, -0.0030968145616331231, -0.0034855712696961689, 
    -0.0038666256889056151, -0.0042200585257370742, -0.0045224392899152225, 
    -0.0047492653819837744, -0.0048778431110738521, -0.0048901572511902231, 
    -0.0047753660369537427, -0.0045315651259375317, -0.0041665305960525492, 
    -0.003697369758510401, -0.0031490549507664544, -0.0025520382019135592, 
    -0.001939234488329548, -0.0013428063552969353, -0.00079120605728410435, 
    -0.00030688867075227366, 9.4966327107771898e-05, 0.00040664623050540235, 
    0.00062707162987661082, 0.000760259882542814, 0.00081343093096059016, 
    0.00079518420165331535, 0.00071407860163612215, 0.00057780930813553465, 
    0.00039308638477879954, 0.00016611253654497831, -9.6518421237943479e-05, 
    -0.000386795004743427, -0.00069442941208202062, -0.0010064511211118348, 
    -0.0013074072793541349, -0.001580230478452147, -0.0018076315586024706, 
    -0.0019738161704596796, -0.0020662049303837365, -0.002076871428446635, 
    -0.0020034603159237406, -0.0018494870247084173, -0.0016239490254297512, 
    -0.0013403407472858358, -0.0010151956263456719, -0.00066635950258072069, 
    -0.00031128213704888599, 3.4358092362807248e-05, 0.00035743727886025417, 
    0.00064747039387124338, 0.00089618357252701283, 0.0010969296880334746, 
    0.0012443405174624952, 0.001334340187982046, 0.0013643916825004905, 
    0.0013337676144887303, 0.0012436578600651727, 0.0010970215252724188, 
    0.0008982621387763031, 0.0006527678959720464, 0.00036638616648409128, 
    4.4956013196733495e-05, -0.00030602159709026174, -0.00068145985814066674, 
    -0.0010765042452802278, -0.0014860030481213158, -0.0019037931622110111, 
    -0.0023219114068903685, -0.0027300059089628943, -0.003115156977489153, 
    -0.0034623055767281042, -0.0037553457821125364, -0.0039787764842409302, 
    -0.004119603707994645, -0.0041691448734731381, -0.0041243028736555739, 
    -0.0039880975587306775, -0.0037693195527673381, -0.0034814230978503584, 
    -0.0031408421065050617, -0.00276503751302955, -0.0023706445863278082, 
    -0.0019719906264960407, -0.0015801777743526179, -0.0012028288705349332, 
    -0.00084444557807096532, -0.00050724922345650534, 
    -0.00019227356741622649, 9.956508609250365e-05, 0.00036668343882473065, 
    0.00060648387805078659, 0.00081548247625815745, 0.00098981846337280362, 
    0.0011259741210851899, 0.0012215492421849177, 0.0012759612966093722, 
    0.0012910047322922135, 0.0012712021419705338, 0.0012239006754659117, 
    0.0011591207238393938, 0.001089054364220938, 0.0010272235286511047, 
    0.00098730538755417642, 0.00098169100606434892, 0.0010199148527304926, 
    0.0011072294122117714, 0.0012435261441522216, 0.0014228939742071118, 
    0.0016338418583976429, 0.0018602648255466017, 0.0020829933730577483, 
    0.0022817758037165462, 0.0024374577507607297, 0.0025341010318504983, 
    0.0025607893775230831, 0.0025128556167450357, 0.0023923909069299074, 
    0.0022079601199690071, 0.0019736292832975523, 0.0017074573850622164, 
    0.0014296529075493117, 0.0011606355936310318, 0.00091917539382637369, 
    0.00072084055536623904, 0.00057686364803735896, 0.00049349740083854407, 
    0.00047181529351450642, 0.00050794572470692369, 0.00059352849377878204, 
    0.00071638785200575411, 0.00086138492225784949, 0.0010115043262261306, 
    0.0011492488309572499, 0.0012582799433529697, 0.0013252172307847594, 
    0.0013413653025504927, 0.0013039385206914729, 0.0012165205466171287, 
    0.0010885606415164018, 0.00093395462851390918, 0.00076901744680169979, 
    0.00061027372127588672, 0.00047251528520080152, 0.00036739496576079875, 
    0.00030271190083472989, 0.00028240917020518167, 0.00030710807508984938, 
    0.00037511124525736148, 0.00048354733618217511, 0.00062946160185234237, 
    0.00081057568620460996, 0.0010254955547562179, 0.0012733033157490215, 
    0.0015526018183529377, 0.001860322320629895, 0.0021906260426979465, 
    0.0025343667128597401, 0.0028792681802434746, 0.0032108522884050795, 
    0.0035138863358380986, 0.003773997747285639, 0.0039791291151600166, 
    0.0041205651450281185, 0.0041934007099732034, 0.00419646197116888, 
    0.0041318073231923682, 0.0040040255885400366, 0.0038194875541721794, 
    0.0035856973200696519, 0.0033107770312021815, 0.0030030932999964574, 
    0.0026709606522373522, 0.0023224395188128424, 0.0019651817063838185, 
    0.0016062766710213726, 0.0012521188872844438, 0.00090828557703135444, 
    0.00057947264099918487, 0.00026947690075904287, -1.8725409328688763e-05, 
    -0.00028285043894920946, -0.00052113815473290854, -0.0007321550686569476, 
    -0.00091458853215452892, -0.0010670111295365576, -0.0011877310501057685, 
    -0.0012748201339046589, -0.0013263643389891616, -0.0013409627018505198, 
    -0.0013184135603176695, -0.0012604097798191746, -0.0011711622958423338, 
    -0.0010576534910825444, -0.00092946930974930481, -0.0007980803102000764, 
    -0.0006756660610590169, -0.0005735538933367728, -0.00050057633219257789, 
    -0.00046153396266465077, -0.00045608133437090829, 
    -0.00047823611461649798, -0.00051675041653498929, 
    -0.00055636126095442572, -0.00057974558720239803, 
    -0.00056981938500503832, -0.00051187873889075696, 
    -0.00039509584467614504, -0.00021328663213536058, 3.4963766995284827e-05, 
    0.00034647797056550436, 0.00071373704118697092, 0.0011250920106571135, 
    0.0015652886926304016, 0.0020164940273460471, 0.0024599070102779728, 
    0.0028776862590861505, 0.0032546551961804928, 0.0035794505356264855, 
    0.0038448880934024913, 0.0040475953975088498, 0.0041872187254764562, 
    0.0042653966391186064, 0.0042847322774556065, 0.0042479029233809425, 
    0.0041569739476453515, 0.0040130196270735091, 0.0038160418332512354, 
    0.0035652188684634463, 0.0032594007034060539, 0.0028978711464100726, 
    0.0024811889635826985, 0.0020119911335931642, 0.001495690720142727, 
    0.00094085143789480324, 0.00035912429383600614, -0.00023532600977150582, 
    -0.00082686053858654874, -0.0013997545811774478, -0.0019396141634409774, 
    -0.0024344404019083937, -0.0028750924172902975, -0.0032551045497932253, 
    -0.0035700248012502998, -0.0038165930534071568, -0.0039921573064557233, 
    -0.0040944945740372827, -0.0041220319240065457, -0.004074346434918814, 
    -0.003952759101200836, -0.0037608749167309945, -0.0035049612857817177, 
    -0.0031940207127979293, -0.0028394161568947415, -0.0024540254332567871, 
    -0.0020509699134787047, -0.0016422220387888472, -0.0012374178284572167, 
    -0.00084324474544094014, -0.00046366781288018614, 
    -0.00010101579092114013, 0.00024234789874750406, 0.00056225298361841898, 
    0.00085145437592425003, 0.0010993793172874476, 0.0012930634157435937, 
    0.0014190694170347399, 0.0014658803782977813, 0.0014260605745814265, 
    0.001297713162278692, 0.0010848656146605355, 0.0007969024321311973, 
    0.00044731439892274226, 5.2150563178284437e-05, -0.00037152627466755395, 
    -0.00080690292537554406, -0.0012383349754567588, -0.0016519216547715686, 
    -0.0020357833275551135, -0.0023800376586546649, -0.002676634565928909, 
    -0.0029190836873623457, -0.0031023077425790324, -0.0032226364086924402, 
    -0.0032780606139151481, -0.0032686371653441143, -0.0031970311605705507, 
    -0.0030689706690714517, -0.0028935273148502604, -0.0026830027139163369, 
    -0.0024524930182049159, -0.0022190157018587356, -0.0020003042739916437, 
    -0.0018134341621333372, -0.0016734093072484032, -0.0015919762609046513, 
    -0.0015767294657330299, -0.0016306195616688879, -0.0017519573636465384, 
    -0.0019349642522148549, -0.002170777488793468, -0.0024486125840990931, 
    -0.0027567882382577317, -0.0030833224626778824, -0.0034161321606507593, 
    -0.0037429005134731927, -0.0040509918610143738, -0.0043275455856887184, 
    -0.004559997930226367, -0.0047369283406087231, -0.0048491142894725118, 
    -0.0048905456321248642, -0.0048590705731639686, -0.0047565328301694496, 
    -0.004588305336255807, -0.0043623896992770507, -0.004088240593619381, 
    -0.0037756089387649501, -0.0034335600646051376, -0.0030697779264014209, 
    -0.0026902751668427989, -0.0022994652257629037, -0.0019006315506163716, 
    -0.0014967238868131259, -0.0010913808409089855, -0.00069003542704392125, 
    -0.00030082330134941718, 6.4963774365567675e-05, 0.00039318963505629277, 
    0.0006680990235671875, 0.00087432366287663334, 0.00099933230508152679, 
    0.0010357823317410069, 0.00098318743148909245, 0.00084847574939123918, 
    0.00064531114480057483, 0.00039224457359603832, 0.00011014987503688099, 
    -0.00018051042154434299, -0.00046214649277808069, 
    -0.00072168359425806841, -0.0009513432481188846, -0.0011485385689076226, 
    -0.0013151761707870767, -0.0014566432314758676, -0.0015806958173898572, 
    -0.0016964807597641489, -0.0018136404777801592, -0.0019415612415590641, 
    -0.0020887176943875244, -0.0022620560269048461, -0.0024664771874652381, 
    -0.0027044619565663084, -0.0029759554405637363, -0.0032784634516543074, 
    -0.0036073602936845684, -0.003956355747819734, -0.0043179920603664901, 
    -0.0046842030883365538, -0.0050468592755549459, -0.00539823264297957, 
    -0.0057312579947286545, -0.0060395119660459438, -0.0063170549902842061, 
    -0.0065582247888110136, -0.0067577646363720543, -0.0069113435789329601, 
    -0.0070164861734676029, -0.0070736741148230628, -0.0070872475037156626, 
    -0.0070657817935470737, -0.0070217882158214676, -0.006970611580052001, 
    -0.0069288528280298505, -0.0069125318137136594, -0.0069353398454851207, 
    -0.0070072763753072755, -0.0071336873920634777, -0.0073147156021533075, 
    -0.0075451269061256893, -0.0078143270489834191, -0.008106726036498247, 
    -0.0084024820646963847, -0.0086788962108824749, -0.0089124640119553084, 
    -0.009081316688711101, -0.0091674695731747604, -0.0091583286205606015, 
    -0.0090472364500955322, -0.0088330825649715321, -0.0085192661965144169, 
    -0.0081122690055081027, -0.0076202400768470308, -0.0070518507184730234, 
    -0.0064157104659833836, -0.005720465931401077, -0.0049754324305983167, 
    -0.0041915141932172334, -0.0033819505945925283, -0.0025626711371137252, 
    -0.0017519497103133368, -0.00096945576895910888, -0.00023479515258180395, 
    0.00043418224358809097, 0.0010230701954112237, 0.0015222620437521637, 
    0.0019277188650984644, 0.0022410214634158419, 0.0024686786205474834, 
    0.0026207548023559619, 0.0027090979157790946, 0.0027454970252029842, 
    0.0027401574964907166, 0.0027005843524692255, 0.0026312602924587207, 
    0.0025339459459335226, 0.0024085254094407763, 0.0022541415740659084, 
    0.0020702312229979748, 0.0018573553543460707, 0.0016176677898689803, 
    0.0013549891373341421, 0.0010746393754001069, 0.00078296387910494652, 
    0.00048663374574356243, 0.00019174016491631788, -9.7289629821021477e-05, 
    -0.00037869927369197298, -0.00065393051672173619, 
    -0.00092743739817950969, -0.0012054903726886799, -0.0014943187294034026, 
    -0.0017979427861659599, -0.0021162489092838169, -0.0024435849596384819, 
    -0.0027680827201380653, -0.0030719766314860021, -0.0033330378047196261, 
    -0.0035270632732463118, -0.0036310210017768646, -0.003626039932914599, 
    -0.0034997325084431714, -0.0032474393839279571, -0.0028724156585520719, 
    -0.0023850326646015826, -0.0018012788151708086, -0.0011408957384943753, 
    -0.00042552762191802167, 0.00032285008292066921, 0.0010830218725328979, 
    0.0018350801041050609, 0.0025604844503018735, 0.0032419878751630275, 
    0.0038634799666966736, 0.0044100370155737423, 0.0048681894756527162, 
    0.0052262649211940069, 0.0054748729486838723, 0.0056073919383149758, 
    0.0056204059699746624, 0.005514240546019792, 0.005293572948977243, 
    0.0049681362022330573, 0.0045533059310134795, 0.0040703116011888661, 
    0.0035456750199356823, 0.0030098367138334811, 0.002494925916612609, 
    0.0020320166817960252, 0.0016483186076660349, 0.0013647684644823067, 
    0.0011943977795169317, 0.0011416684170343038, 0.0012028332020260113, 
    0.0013672248496170935, 0.0016193220689686809, 0.0019412115186090858, 
    0.0023150332388773304, 0.0027249881325686356, 0.0031584805040611257, 
    0.0036062981611492792, 0.0040618294956252582, 0.0045197259483114836, 
    0.0049744355038284192, 0.0054189782985010378, 0.005844210823313269, 
    0.0062387678654075443, 0.0065895229827480067, 0.0068825745505557579, 
    0.0071045325890884432, 0.0072439331960175123, 0.0072925320517621805, 
    0.0072463178837787892, 0.0071060329026631343, 0.0068771304361516968, 
    0.0065692179158246908, 0.0061949304370786671, 0.0057685846170976033, 
    0.0053046366551389376, 0.0048163387726694101, 0.0043147575238160624, 
    0.0038083806805735533, 0.0033033091073871469, 0.0028040227889529982, 
    0.0023145046454062551, 0.0018394229704385425, 0.0013849727056872243, 
    0.00095904716501590619, 0.00057061847879677659, 0.00022846987621685013, 
    -6.0359533766643687e-05, -0.0002920794704917012, -0.00046713149347138146, 
    -0.00059045435785127598, -0.00067092540262832451, 
    -0.00071993750740619424, -0.00074943938522258145, 
    -0.00076974609317725321, -0.0007874794020241928, -0.00080424578882163961, 
    -0.00081628816997906801, -0.00081533360138601164, 
    -0.00079045899150438008, -0.00073057843778814835, 
    -0.00062699396993558297, -0.00047532573507643052, 
    -0.00027639891480738237, -3.5955387041102893e-05, 0.00023680238630969077, 
    0.00053126395747171565, 0.00083761449838215432, 0.0011485464058372591, 
    0.0014600025189964072, 0.0017707863193345355, 0.0020812904552194671, 
    0.0023917762548215735, 0.0027009670383238617, 0.0030051972825876606, 
    0.0032984790578104053, 0.0035735206735083725, 0.00382326939961866, 
    0.004042592172991682, 0.0042299245415563123, 0.0043882876680543369, 
    0.004525701342575252, 0.0046547814089262325, 0.0047914896367946122, 
    0.0049530002883165676, 0.0051549596341641645, 0.0054084791152417769, 
    0.0057176086430450277, 0.0060777801373939934, 0.0064758569714869199, 
    0.0068916837640206705, 0.0073007571997101839, 0.0076771999642906204, 
    0.0079964686038345046, 0.0082373976606105806, 0.008383516183696026, 
    0.0084241351735998022, 0.0083555028735333957, 0.0081821798931824112, 
    0.0079180986614518344, 0.0075868856003107124, 0.0072209631332117181, 
    0.0068591567578337245, 0.006543013355707665, 0.0063120038230669254, 
    0.0061986465217506066, 0.0062242039794479023, 0.0063953828364749221, 
    0.0067026319656874724, 0.0071198675807288628, 0.0076059082848078802, 
    0.0081076594518979771, 0.0085651919090684956, 0.0089181491257041869, 
    0.0091124486553255963, 0.0091062795894880453, 0.008874425324872301, 
    0.0084105237107272093, 0.007727134891401052, 0.0068539438928074898, 
    0.0058344905087198131, 0.004721806870153126, 0.0035734585510094645, 
    0.0024463954320918541, 0.0013923445067601258, 0.00045390802236581969, 
    -0.00033816432469310179, -0.00096642021737464797, -0.0014268408575730737, 
    -0.0017275938453514433, -0.0018868348292518172, -0.0019294754360155617, 
    -0.0018836137859877086, -0.0017769942767106785, -0.0016338408060610492, 
    -0.0014726448528761906, -0.0013050239076878966, -0.0011355420034258211, 
    -0.00096246909748367031, -0.00077901686356234229, 
    -0.00057496373260611233, -0.00033831780904078617, 
    -5.7083686842700914e-05, 0.00027886467457374005, 0.00067606666019827421, 
    0.0011358038811666391, 0.0016530194602221711, 0.0022161342213773833, 
    0.0028078787004782542, 0.0034070975864337084, 0.003991183272573153, 
    0.0045386639145459052, 0.0050316033568497632, 0.005457467685552179, 
    0.0058101767288289315, 0.0060904342745404993, 0.0063051902412012938, 
    0.0064665610135918082, 0.0065904532787047099, 0.0066949401016581219, 
    0.0067987958320849763, 0.0069195277781893471, 0.0070712911776500834, 
    0.0072625004379256401, 0.0074941188289336727, 0.0077590388386624071, 
    0.0080428456738108438, 0.0083257574357967629, 0.0085848542674306534, 
    0.0087959227548908055, 0.0089347663217112794, 0.0089778622977218312, 
    0.0089032137171197734, 0.0086918186240846091, 0.0083299737332015872, 
    0.0078122460207961618, 0.007144337481121415, 0.0063451647614091002, 
    0.0054474348917961327, 0.0044962358298620544, 0.0035457804860169776, 
    0.0026542951212667064, 0.0018780643360654244, 0.0012650733360971269, 
    0.00084968311586042624, 0.00064920378583598472, 0.00066294560452058058, 
    0.00087389862559869743, 0.0012520402419860417, 0.0017584616801736693, 
    0.0023491981960928479, 0.002978394467789771, 0.0036008776416147489, 
    0.0041742407693408489, 0.0046609398750090533, 0.0050302923945279455, 
    0.0052606241817891395, 0.0053412238444911376, 0.0052740874045771081, 
    0.0050744702011301509, 0.0047701995030114252, 0.0043989611814954834, 
    0.0040035289829942425, 0.0036257436375770986, 0.0033002685179182316, 
    0.0030499208337806559, 0.0028836218182389877, 0.0027975635484742208, 
    0.0027781277799910371, 0.0028055974090631852, 0.0028568168944728169, 
    0.0029073036312541245, 0.0029330002471710682, 0.0029133913312135717, 
    0.0028362390623259837, 0.002702520307212988, 0.0025301986166890692, 
    0.0023542777019803169, 0.0022219690765857567, 0.0021837648589175759, 
    0.0022826245802152387, 0.002544375918166595, 0.0029717581310340102, 
    0.0035430361396967336, 0.0042149268411106749, 0.0049288650545637053, 
    0.005619342813074267, 0.0062225263062661955, 0.0066835084853909205, 
    0.0069616917477509426, 0.0070327265843371269, 0.0068878777320621528, 
    0.0065310928417218628, 0.0059758615533791514, 0.0052431681536461959, 
    0.0043610681429446145, 0.0033654546071763564, 0.0022991039909770394, 
    0.0012087843540256867, 0.00013980597111866964, -0.00087054289985239873, 
    -0.0017985485634466739, -0.0026374173047940034, -0.0033980597069676447, 
    -0.0041067975795807702, -0.0048002740935826037, -0.0055187688575955652, 
    -0.0062988281098652213, -0.0071668039518171306, -0.0081370718854259852, 
    -0.0092133369191941625, -0.010393653996624751, -0.011674965121869812, 
    -0.013052941823617242, -0.014518218487901802, -0.016049860987275451, 
    -0.017609873917982195, -0.019138950597556405, -0.020555947684977267, 
    -0.021762643426323589, -0.0226529240155653, -0.023125095248749519, 
    -0.023095073904620657, -0.022505190131911355, -0.021330630316602185, 
    -0.019581183063821912, -0.017300910551862985, -0.014565988157510652, 
    -0.011480795688368279, -0.0081735333777772923, -0.0047916150776234458, 
    -0.0014928339832148826, 0.0015629124213077826, 0.0042274391168724028, 
    0.0063783644455004795, 0.0079309219486246897, 0.0088419351918969363 ;

 frequency = 0, 0.12499999406281886, 0.24999998812563773, 
    0.37499998218845659, 0.49999997625127546, 0.62499997031409438, 
    0.74999996437691319, 0.87499995843973211, 0.99999995250255092, 
    1.1249999465653697, 1.2499999406281888, 1.3749999346910076, 
    1.4999999287538264, 1.6249999228166454, 1.7499999168794642, 
    1.874999910942283, 1.9999999050051018, 2.1249998990679209, 
    2.2499998931307394, 2.3749998871935585, 2.4999998812563775, 
    2.6249998753191961, 2.7499998693820151, 2.8749998634448342, 
    2.9999998575076527, 3.1249998515704718, 3.2499998456332908, 
    3.3749998396961094, 3.4999998337589284, 3.624999827821747, 
    3.749999821884566, 3.8749998159473851, 3.9999998100102037, 
    4.1249998040730222, 4.2499997981358417, 4.3749997921986603, 
    4.4999997862614789, 4.6249997803242984, 4.749999774387117, 
    4.8749997684499355, 4.999999762512755, 5.1249997565755736, 
    5.2499997506383922, 5.3749997447012117, 5.4999997387640303, 
    5.6249997328268488, 5.7499997268896683, 5.8749997209524869, 
    5.9999997150153055, 6.124999709078125, 6.2499997031409436, 
    6.3749996972037621, 6.4999996912665816, 6.6249996853294002, 
    6.7499996793922188, 6.8749996734550374, 6.9999996675178568, 
    7.1249996615806754, 7.249999655643494, 7.3749996497063135, 
    7.4999996437691321, 7.6249996378319507, 7.7499996318947701, 
    7.8749996259575887, 7.9999996200204073, 8.1249996140832259, 
    8.2499996081460445, 8.3749996022088649, 8.4999995962716834, 
    8.624999590334502, 8.7499995843973206, 8.8749995784601392, 
    8.9999995725229578, 9.1249995665857782, 9.2499995606485967, 
    9.3749995547114153, 9.4999995487742339, 9.6249995428370525, 
    9.7499995368998711, 9.8749995309626915, 9.99999952502551, 
    10.124999519088329, 10.249999513151147, 10.374999507213966, 
    10.499999501276784, 10.624999495339603, 10.749999489402423, 
    10.874999483465242, 10.999999477528061, 11.124999471590879, 
    11.249999465653698, 11.374999459716516, 11.499999453779337, 
    11.624999447842155, 11.749999441904974, 11.874999435967792, 
    11.999999430030611, 12.12499942409343, 12.24999941815625, 
    12.374999412219069, 12.499999406281887, 12.624999400344706, 
    12.749999394407524, 12.874999388470343, 12.999999382533163, 
    13.124999376595982, 13.2499993706588, 13.374999364721619, 
    13.499999358784438, 13.624999352847256, 13.749999346910075, 
    13.874999340972895, 13.999999335035714, 14.124999329098532, 
    14.249999323161351, 14.374999317224169, 14.499999311286988, 
    14.624999305349808, 14.749999299412627, 14.874999293475446, 
    14.999999287538264, 15.124999281601083, 15.249999275663901, 
    15.374999269726722, 15.49999926378954, 15.624999257852359, 
    15.749999251915177, 15.874999245977996, 15.999999240040815, 
    16.124999234103633, 16.249999228166452, 16.37499922222927, 
    16.499999216292089, 16.624999210354911, 16.74999920441773, 
    16.874999198480548, 16.999999192543367, 17.124999186606185, 
    17.249999180669004, 17.374999174731823, 17.499999168794641, 
    17.62499916285746, 17.749999156920278, 17.874999150983097, 
    17.999999145045916, 18.124999139108738, 18.249999133171556, 
    18.374999127234375, 18.499999121297193, 18.624999115360012, 
    18.749999109422831, 18.874999103485649, 18.999999097548468, 
    19.124999091611286, 19.249999085674105, 19.374999079736924, 
    19.499999073799742, 19.624999067862561, 19.749999061925383, 
    19.874999055988201, 19.99999905005102, 20.124999044113839, 
    20.249999038176657, 20.374999032239476, 20.499999026302294, 
    20.624999020365113, 20.749999014427932, 20.87499900849075, 
    20.999999002553569, 21.124998996616387, 21.249998990679206, 
    21.374998984742028, 21.499998978804847, 21.624998972867665, 
    21.749998966930484, 21.874998960993302, 21.999998955056121, 
    22.12499894911894, 22.249998943181758, 22.374998937244577, 
    22.499998931307395, 22.624998925370214, 22.749998919433033, 
    22.874998913495855, 22.999998907558673, 23.124998901621492, 
    23.24999889568431, 23.374998889747129, 23.499998883809948, 
    23.624998877872766, 23.749998871935585, 23.874998865998403, 
    23.999998860061222, 24.124998854124041, 24.249998848186859, 
    24.374998842249678, 24.4999988363125, 24.624998830375318, 
    24.749998824438137, 24.874998818500956, 24.999998812563774, 
    25.124998806626593, 25.249998800689411, 25.37499879475223, 
    25.499998788815049, 25.624998782877867, 25.749998776940686, 
    25.874998771003504, 25.999998765066326, 26.124998759129145, 
    26.249998753191964, 26.374998747254782, 26.499998741317601, 
    26.624998735380419, 26.749998729443238, 26.874998723506057, 
    26.999998717568875, 27.124998711631694, 27.249998705694512, 
    27.374998699757331, 27.499998693820149, 27.624998687882972, 
    27.74999868194579, 27.874998676008609, 27.999998670071427, 
    28.124998664134246, 28.249998658197065, 28.374998652259883, 
    28.499998646322702, 28.62499864038552, 28.749998634448339, 
    28.874998628511158, 28.999998622573976, 29.124998616636795, 
    29.249998610699617, 29.374998604762435, 29.499998598825254, 
    29.624998592888073, 29.749998586950891, 29.87499858101371, 
    29.999998575076528, 30.124998569139347, 30.249998563202166, 
    30.374998557264984, 30.499998551327803, 30.624998545390621, 
    30.749998539453443, 30.874998533516262, 30.999998527579081, 
    31.124998521641899, 31.249998515704718, 31.374998509767536, 
    31.499998503830355, 31.624998497893174, 31.749998491955992, 
    31.874998486018811, 31.999998480081629, 32.124998474144448, 
    32.249998468207266, 32.374998462270085, 32.499998456332904, 
    32.624998450395722, 32.749998444458541, 32.874998438521359, 
    32.999998432584178, 33.124998426647004, 33.249998420709822, 
    33.374998414772641, 33.499998408835459, 33.624998402898278, 
    33.749998396961097, 33.874998391023915, 33.999998385086734, 
    34.124998379149552, 34.249998373212371, 34.37499836727519, 
    34.499998361338008, 34.624998355400827, 34.749998349463645, 
    34.874998343526464, 34.999998337589282, 35.124998331652101, 
    35.24999832571492, 35.374998319777738, 35.499998313840557, 
    35.624998307903375, 35.749998301966194, 35.874998296029013, 
    35.999998290091831, 36.12499828415465, 36.249998278217475, 
    36.374998272280294, 36.499998266343113, 36.624998260405931, 
    36.74999825446875, 36.874998248531568, 36.999998242594387, 
    37.124998236657206, 37.249998230720024, 37.374998224782843, 
    37.499998218845661, 37.62499821290848, 37.749998206971298, 
    37.874998201034117, 37.999998195096936, 38.124998189159754, 
    38.249998183222573, 38.374998177285391, 38.49999817134821, 
    38.624998165411029, 38.749998159473847, 38.874998153536666, 
    38.999998147599484, 39.124998141662303, 39.249998135725122, 
    39.374998129787947, 39.499998123850766, 39.624998117913584, 
    39.749998111976403, 39.874998106039222, 39.99999810010204, 
    40.124998094164859, 40.249998088227677, 40.374998082290496, 
    40.499998076353315, 40.624998070416133, 40.749998064478952, 
    40.87499805854177, 40.999998052604589, 41.124998046667407, 
    41.249998040730226, 41.374998034793045, 41.499998028855863, 
    41.624998022918682, 41.7499980169815, 41.874998011044319, 
    41.999998005107138, 42.124997999169956, 42.249997993232775, 
    42.374997987295593, 42.499997981358412, 42.624997975421238, 
    42.749997969484056, 42.874997963546875, 42.999997957609693, 
    43.124997951672512, 43.249997945735331, 43.374997939798149, 
    43.499997933860968, 43.624997927923786, 43.749997921986605, 
    43.874997916049423, 43.999997910112242, 44.124997904175061, 
    44.249997898237879, 44.374997892300698, 44.499997886363516, 
    44.624997880426335, 44.749997874489154, 44.874997868551972, 
    44.999997862614791, 45.124997856677609, 45.249997850740428, 
    45.374997844803246, 45.499997838866065, 45.624997832928884, 
    45.749997826991709, 45.874997821054528, 45.999997815117347, 
    46.124997809180165, 46.249997803242984, 46.374997797305802, 
    46.499997791368621, 46.624997785431439, 46.749997779494258, 
    46.874997773557077, 46.999997767619895, 47.124997761682714, 
    47.249997755745532, 47.374997749808351, 47.49999774387117, 
    47.624997737933988, 47.749997731996807, 47.874997726059625, 
    47.999997720122444, 48.124997714185263, 48.249997708248081, 
    48.3749977023109, 48.499997696373718, 48.624997690436537, 
    48.749997684499355, 48.874997678562181, 48.999997672625, 
    49.124997666687818, 49.249997660750637, 49.374997654813455, 
    49.499997648876274, 49.624997642939093, 49.749997637001911, 
    49.87499763106473, 49.999997625127548, 50.124997619190367, 
    50.249997613253186, 50.374997607316004, 50.499997601378823, 
    50.624997595441641, 50.74999758950446, 50.874997583567279, 
    50.999997577630097, 51.124997571692916, 51.249997565755734, 
    51.374997559818553, 51.499997553881371, 51.62499754794419, 
    51.749997542007009, 51.874997536069827, 51.999997530132653, 
    52.124997524195471, 52.24999751825829, 52.374997512321109, 
    52.499997506383927, 52.624997500446746, 52.749997494509564, 
    52.874997488572383, 52.999997482635202, 53.12499747669802, 
    53.249997470760839, 53.374997464823657, 53.499997458886476, 
    53.624997452949295, 53.749997447012113, 53.874997441074932, 
    53.99999743513775, 54.124997429200569, 54.249997423263387, 
    54.374997417326206, 54.499997411389025, 54.624997405451843, 
    54.749997399514662, 54.87499739357748, 54.999997387640299, 
    55.124997381703125, 55.249997375765943, 55.374997369828762, 
    55.49999736389158, 55.624997357954399, 55.749997352017218, 
    55.874997346080036, 55.999997340142855, 56.124997334205673, 
    56.249997328268492, 56.374997322331311, 56.499997316394129, 
    56.624997310456948, 56.749997304519766, 56.874997298582585, 
    56.999997292645403, 57.124997286708222, 57.249997280771041, 
    57.374997274833859, 57.499997268896678, 57.624997262959496, 
    57.749997257022315, 57.874997251085134, 57.999997245147952, 
    58.124997239210771, 58.249997233273589, 58.374997227336415, 
    58.499997221399234, 58.624997215462052, 58.749997209524871, 
    58.874997203587689, 58.999997197650508, 59.124997191713327, 
    59.249997185776145, 59.374997179838964, 59.499997173901782, 
    59.624997167964601, 59.74999716202742, 59.874997156090238, 
    59.999997150153057, 60.124997144215875, 60.249997138278694, 
    60.374997132341512, 60.499997126404331, 60.62499712046715, 
    60.749997114529968, 60.874997108592787, 60.999997102655605, 
    61.124997096718424, 61.249997090781243, 61.374997084844061, 
    61.499997078906887, 61.624997072969705, 61.749997067032524, 
    61.874997061095343, 61.999997055158161, 62.12499704922098, 
    62.249997043283798, 62.374997037346617, 62.499997031409436, 
    62.624997025472254, 62.749997019535073, 62.874997013597891, 
    62.99999700766071, 63.124997001723528, 63.249996995786347, 
    63.374996989849166, 63.499996983911984, 63.624996977974803, 
    63.749996972037621, 63.87499696610044, 63.999996960163259, 
    64.124996954226077, 64.249996948288896, 64.374996942351714, 
    64.499996936414533, 64.624996930477351, 64.74999692454017, 
    64.874996918602989, 64.999996912665807, 65.124996906728626, 
    65.249996900791444, 65.374996894854263, 65.499996888917082, 
    65.6249968829799, 65.749996877042719, 65.874996871105537, 
    65.999996865168356, 66.124996859231175, 66.249996853294007, 
    66.374996847356826, 66.499996841419645, 66.624996835482463, 
    66.749996829545282, 66.8749968236081, 66.999996817670919, 
    67.124996811733737, 67.249996805796556, 67.374996799859375, 
    67.499996793922193, 67.624996787985012, 67.74999678204783, 
    67.874996776110649, 67.999996770173468, 68.124996764236286, 
    68.249996758299105, 68.374996752361923, 68.499996746424742, 
    68.62499674048756, 68.749996734550379, 68.874996728613198, 
    68.999996722676016, 69.124996716738835, 69.249996710801653, 
    69.374996704864472, 69.499996698927291, 69.624996692990109, 
    69.749996687052928, 69.874996681115746, 69.999996675178565, 
    70.124996669241384, 70.249996663304202, 70.374996657367021, 
    70.499996651429839, 70.624996645492658, 70.749996639555476, 
    70.874996633618295, 70.999996627681114, 71.124996621743932, 
    71.249996615806751, 71.374996609869569, 71.499996603932388, 
    71.624996597995207, 71.749996592058025, 71.874996586120844, 
    71.999996580183662, 72.124996574246481, 72.2499965683093, 
    72.374996562372118, 72.499996556434951, 72.624996550497769, 
    72.749996544560588, 72.874996538623407, 72.999996532686225, 
    73.124996526749044, 73.249996520811862, 73.374996514874681, 
    73.4999965089375, 73.624996503000318, 73.749996497063137, 
    73.874996491125955, 73.999996485188774, 74.124996479251593, 
    74.249996473314411, 74.37499646737723, 74.499996461440048, 
    74.624996455502867, 74.749996449565685, 74.874996443628504, 
    74.999996437691323, 75.124996431754141, 75.24999642581696, 
    75.374996419879778, 75.499996413942597, 75.624996408005416, 
    75.749996402068234, 75.874996396131053, 75.999996390193871, 
    76.12499638425669, 76.249996378319508, 76.374996372382327, 
    76.499996366445146, 76.624996360507964, 76.749996354570783, 
    76.874996348633601, 76.99999634269642, 77.124996336759239, 
    77.249996330822057, 77.374996324884876, 77.499996318947694, 
    77.624996313010513, 77.749996307073332, 77.87499630113615, 
    77.999996295198969, 78.124996289261787, 78.249996283324606, 
    78.374996277387424, 78.499996271450243, 78.624996265513062, 
    78.749996259575894, 78.874996253638713, 78.999996247701532, 
    79.12499624176435, 79.249996235827169, 79.374996229889987, 
    79.499996223952806, 79.624996218015625, 79.749996212078443, 
    79.874996206141262, 79.99999620020408, 80.124996194266899, 
    80.249996188329717, 80.374996182392536, 80.499996176455355, 
    80.624996170518173, 80.749996164580992, 80.87499615864381, 
    80.999996152706629, 81.124996146769448, 81.249996140832266, 
    81.374996134895085, 81.499996128957903, 81.624996123020722, 
    81.749996117083541, 81.874996111146359, 81.999996105209178, 
    82.124996099271996, 82.249996093334815, 82.374996087397633, 
    82.499996081460452, 82.624996075523271, 82.749996069586089, 
    82.874996063648908, 82.999996057711726, 83.124996051774545, 
    83.249996045837364, 83.374996039900182, 83.499996033963001, 
    83.624996028025819, 83.749996022088638, 83.874996016151457, 
    83.999996010214275, 84.124996004277094, 84.249995998339912, 
    84.374995992402731, 84.499995986465549, 84.624995980528368, 
    84.749995974591187, 84.874995968654005, 84.999995962716824, 
    85.124995956779657, 85.249995950842475, 85.374995944905294, 
    85.499995938968112, 85.624995933030931, 85.74999592709375, 
    85.874995921156568, 85.999995915219387, 86.124995909282205, 
    86.249995903345024, 86.374995897407842, 86.499995891470661, 
    86.62499588553348, 86.749995879596298, 86.874995873659117, 
    86.999995867721935, 87.124995861784754, 87.249995855847573, 
    87.374995849910391, 87.49999584397321, 87.624995838036028, 
    87.749995832098847, 87.874995826161665, 87.999995820224484, 
    88.124995814287303, 88.249995808350121, 88.37499580241294, 
    88.499995796475758, 88.624995790538577, 88.749995784601396, 
    88.874995778664214, 88.999995772727033, 89.124995766789851, 
    89.24999576085267, 89.374995754915489, 89.499995748978307, 
    89.624995743041126, 89.749995737103944, 89.874995731166763, 
    89.999995725229581, 90.1249957192924, 90.249995713355219, 
    90.374995707418037, 90.499995701480856, 90.624995695543674, 
    90.749995689606493, 90.874995683669312, 90.99999567773213, 
    91.124995671794949, 91.249995665857767, 91.3749956599206, 
    91.499995653983419, 91.624995648046237, 91.749995642109056, 
    91.874995636171874, 91.999995630234693, 92.124995624297512, 
    92.24999561836033, 92.374995612423149, 92.499995606485967, 
    92.624995600548786, 92.749995594611605, 92.874995588674423, 
    92.999995582737242, 93.12499557680006, 93.249995570862879, 
    93.374995564925698, 93.499995558988516, 93.624995553051335, 
    93.749995547114153, 93.874995541176972, 93.99999553523979, 
    94.124995529302609, 94.249995523365428, 94.374995517428246, 
    94.499995511491065, 94.624995505553883, 94.749995499616702, 
    94.874995493679521, 94.999995487742339, 95.124995481805158, 
    95.249995475867976, 95.374995469930795, 95.499995463993613, 
    95.624995458056432, 95.749995452119251, 95.874995446182069, 
    95.999995440244888, 96.124995434307706, 96.249995428370525, 
    96.374995422433344, 96.499995416496162, 96.624995410558981, 
    96.749995404621799, 96.874995398684618, 96.999995392747437, 
    97.124995386810255, 97.249995380873074, 97.374995374935892, 
    97.499995368998711, 97.624995363061529, 97.749995357124362, 
    97.874995351187181, 97.999995345249999, 98.124995339312818, 
    98.249995333375637, 98.374995327438455, 98.499995321501274, 
    98.624995315564092, 98.749995309626911, 98.87499530368973, 
    98.999995297752548, 99.124995291815367, 99.249995285878185, 
    99.374995279941004, 99.499995274003822, 99.624995268066641, 
    99.74999526212946, 99.874995256192278, 99.999995250255097, 
    100.12499524431792, 100.24999523838073, 100.37499523244355, 
    100.49999522650637, 100.62499522056919, 100.74999521463201, 
    100.87499520869483, 100.99999520275765, 101.12499519682046, 
    101.24999519088328, 101.3749951849461, 101.49999517900892, 
    101.62499517307174, 101.74999516713456, 101.87499516119738, 
    101.99999515526019, 102.12499514932301, 102.24999514338583, 
    102.37499513744865, 102.49999513151147, 102.62499512557429, 
    102.74999511963711, 102.87499511369992, 102.99999510776274, 
    103.12499510182556, 103.24999509588838, 103.3749950899512, 
    103.49999508401402, 103.62499507807684, 103.74999507213965, 
    103.87499506620247, 103.99999506026531, 104.12499505432812, 
    104.24999504839094, 104.37499504245376, 104.49999503651658, 
    104.6249950305794, 104.74999502464222, 104.87499501870504, 
    104.99999501276785, 105.12499500683067, 105.24999500089349, 
    105.37499499495631, 105.49999498901913, 105.62499498308195, 
    105.74999497714477, 105.87499497120758, 105.9999949652704, 
    106.12499495933322, 106.24999495339604, 106.37499494745886, 
    106.49999494152168, 106.6249949355845, 106.74999492964731, 
    106.87499492371013, 106.99999491777295, 107.12499491183577, 
    107.24999490589859, 107.37499489996141, 107.49999489402423, 
    107.62499488808704, 107.74999488214986, 107.87499487621268, 
    107.9999948702755, 108.12499486433832, 108.24999485840114, 
    108.37499485246396, 108.49999484652677, 108.62499484058959, 
    108.74999483465241, 108.87499482871523, 108.99999482277805, 
    109.12499481684087, 109.24999481090369, 109.37499480496651, 
    109.49999479902932, 109.62499479309214, 109.74999478715496, 
    109.87499478121778, 109.9999947752806, 110.12499476934342, 
    110.24999476340625, 110.37499475746907, 110.49999475153189, 
    110.62499474559471, 110.74999473965752, 110.87499473372034, 
    110.99999472778316, 111.12499472184598, 111.2499947159088, 
    111.37499470997162, 111.49999470403444, 111.62499469809725, 
    111.74999469216007, 111.87499468622289, 111.99999468028571, 
    112.12499467434853, 112.24999466841135, 112.37499466247417, 
    112.49999465653698, 112.6249946505998, 112.74999464466262, 
    112.87499463872544, 112.99999463278826, 113.12499462685108, 
    113.2499946209139, 113.37499461497671, 113.49999460903953, 
    113.62499460310235, 113.74999459716517, 113.87499459122799, 
    113.99999458529081, 114.12499457935363, 114.24999457341644, 
    114.37499456747926, 114.49999456154208, 114.6249945556049, 
    114.74999454966772, 114.87499454373054, 114.99999453779336, 
    115.12499453185617, 115.24999452591899, 115.37499451998181, 
    115.49999451404463, 115.62499450810745, 115.74999450217027, 
    115.87499449623309, 115.9999944902959, 116.12499448435872, 
    116.24999447842154, 116.37499447248436, 116.49999446654718, 
    116.62499446061001, 116.74999445467283, 116.87499444873565, 
    116.99999444279847, 117.12499443686129, 117.2499944309241, 
    117.37499442498692, 117.49999441904974, 117.62499441311256, 
    117.74999440717538, 117.8749944012382, 117.99999439530102, 
    118.12499438936383, 118.24999438342665, 118.37499437748947, 
    118.49999437155229, 118.62499436561511, 118.74999435967793, 
    118.87499435374075, 118.99999434780356, 119.12499434186638, 
    119.2499943359292, 119.37499432999202, 119.49999432405484, 
    119.62499431811766, 119.74999431218048, 119.87499430624329, 
    119.99999430030611, 120.12499429436893, 120.24999428843175, 
    120.37499428249457, 120.49999427655739, 120.62499427062021, 
    120.74999426468302, 120.87499425874584, 120.99999425280866, 
    121.12499424687148, 121.2499942409343, 121.37499423499712, 
    121.49999422905994, 121.62499422312275, 121.74999421718557, 
    121.87499421124839, 121.99999420531121, 122.12499419937403, 
    122.24999419343685, 122.37499418749967, 122.49999418156249, 
    122.6249941756253, 122.74999416968812, 122.87499416375096, 
    122.99999415781377, 123.12499415187659, 123.24999414593941, 
    123.37499414000223, 123.49999413406505, 123.62499412812787, 
    123.74999412219069, 123.8749941162535, 123.99999411031632, 
    124.12499410437914, 124.24999409844196, 124.37499409250478, 
    124.4999940865676, 124.62499408063042, 124.74999407469323, 
    124.87499406875605, 124.99999406281887, 125.12499405688169, 
    125.24999405094451, 125.37499404500733, 125.49999403907015, 
    125.62499403313296, 125.74999402719578, 125.8749940212586, 
    125.99999401532142, 126.12499400938424, 126.24999400344706, 
    126.37499399750988, 126.49999399157269, 126.62499398563551, 
    126.74999397969833, 126.87499397376115, 126.99999396782397, 
    127.12499396188679, 127.24999395594961, 127.37499395001242, 
    127.49999394407524, 127.62499393813806, 127.74999393220088, 
    127.8749939262637, 127.99999392032652, 128.12499391438934, 
    128.24999390845215, 128.37499390251497, 128.49999389657779, 
    128.62499389064061, 128.74999388470343, 128.87499387876625, 
    128.99999387282907, 129.12499386689188, 129.2499938609547, 
    129.37499385501752, 129.49999384908034, 129.62499384314316, 
    129.74999383720598, 129.8749938312688, 129.99999382533161, 
    130.12499381939443, 130.24999381345725, 130.37499380752007, 
    130.49999380158289, 130.62499379564571, 130.74999378970853, 
    130.87499378377134, 130.99999377783416, 131.12499377189698, 
    131.2499937659598, 131.37499376002262, 131.49999375408544, 
    131.62499374814826, 131.74999374221107, 131.87499373627389, 
    131.99999373033671, 132.12499372439953, 132.24999371846235, 
    132.3749937125252, 132.49999370658801, 132.62499370065083, 
    132.74999369471365, 132.87499368877647, 132.99999368283929, 
    133.12499367690211, 133.24999367096493, 133.37499366502774, 
    133.49999365909056, 133.62499365315338, 133.7499936472162, 
    133.87499364127902, 133.99999363534184, 134.12499362940466, 
    134.24999362346747, 134.37499361753029, 134.49999361159311, 
    134.62499360565593, 134.74999359971875, 134.87499359378157, 
    134.99999358784439, 135.1249935819072, 135.24999357597002, 
    135.37499357003284, 135.49999356409566, 135.62499355815848, 
    135.7499935522213, 135.87499354628412, 135.99999354034694, 
    136.12499353440975, 136.24999352847257, 136.37499352253539, 
    136.49999351659821, 136.62499351066103, 136.74999350472385, 
    136.87499349878667, 136.99999349284948, 137.1249934869123, 
    137.24999348097512, 137.37499347503794, 137.49999346910076, 
    137.62499346316358, 137.7499934572264, 137.87499345128921, 
    137.99999344535203, 138.12499343941485, 138.24999343347767, 
    138.37499342754049, 138.49999342160331, 138.62499341566613, 
    138.74999340972894, 138.87499340379176, 138.99999339785458, 
    139.1249933919174, 139.24999338598022, 139.37499338004304, 
    139.49999337410586, 139.62499336816867, 139.74999336223149, 
    139.87499335629431, 139.99999335035713, 140.12499334441995, 
    140.24999333848277, 140.37499333254559, 140.4999933266084, 
    140.62499332067122, 140.74999331473404, 140.87499330879686, 
    140.99999330285968, 141.1249932969225, 141.24999329098532, 
    141.37499328504813, 141.49999327911095, 141.62499327317377, 
    141.74999326723659, 141.87499326129941, 141.99999325536223, 
    142.12499324942505, 142.24999324348786, 142.37499323755068, 
    142.4999932316135, 142.62499322567632, 142.74999321973914, 
    142.87499321380196, 142.99999320786478, 143.12499320192759, 
    143.24999319599041, 143.37499319005323, 143.49999318411605, 
    143.62499317817887, 143.74999317224169, 143.87499316630451, 
    143.99999316036732, 144.12499315443014, 144.24999314849296, 
    144.37499314255578, 144.4999931366186, 144.62499313068142, 
    144.74999312474424, 144.87499311880705, 144.9999931128699, 
    145.12499310693272, 145.24999310099554, 145.37499309505836, 
    145.49999308912118, 145.62499308318399, 145.74999307724681, 
    145.87499307130963, 145.99999306537245, 146.12499305943527, 
    146.24999305349809, 146.37499304756091, 146.49999304162372, 
    146.62499303568654, 146.74999302974936, 146.87499302381218, 
    146.999993017875, 147.12499301193782, 147.24999300600064, 
    147.37499300006345, 147.49999299412627, 147.62499298818909, 
    147.74999298225191, 147.87499297631473, 147.99999297037755, 
    148.12499296444037, 148.24999295850319, 148.374992952566, 
    148.49999294662882, 148.62499294069164, 148.74999293475446, 
    148.87499292881728, 148.9999929228801, 149.12499291694292, 
    149.24999291100573, 149.37499290506855, 149.49999289913137, 
    149.62499289319419, 149.74999288725701, 149.87499288131983, 
    149.99999287538265, 150.12499286944546, 150.24999286350828, 
    150.3749928575711, 150.49999285163392, 150.62499284569674, 
    150.74999283975956, 150.87499283382238, 150.99999282788519, 
    151.12499282194801, 151.24999281601083, 151.37499281007365, 
    151.49999280413647, 151.62499279819929, 151.74999279226211, 
    151.87499278632492, 151.99999278038774, 152.12499277445056, 
    152.24999276851338, 152.3749927625762, 152.49999275663902, 
    152.62499275070184, 152.74999274476465, 152.87499273882747, 
    152.99999273289029, 153.12499272695311, 153.24999272101593, 
    153.37499271507875, 153.49999270914157, 153.62499270320438, 
    153.7499926972672, 153.87499269133002, 153.99999268539284, 
    154.12499267945566, 154.24999267351848, 154.3749926675813, 
    154.49999266164411, 154.62499265570693, 154.74999264976975, 
    154.87499264383257, 154.99999263789539, 155.12499263195821, 
    155.24999262602103, 155.37499262008384, 155.49999261414666, 
    155.62499260820948, 155.7499926022723, 155.87499259633512, 
    155.99999259039794, 156.12499258446076, 156.24999257852357, 
    156.37499257258639, 156.49999256664921, 156.62499256071203, 
    156.74999255477485, 156.87499254883767, 156.99999254290049, 
    157.1249925369633, 157.24999253102612, 157.37499252508894, 
    157.49999251915179, 157.62499251321461, 157.74999250727743, 
    157.87499250134024, 157.99999249540306, 158.12499248946588, 
    158.2499924835287, 158.37499247759152, 158.49999247165434, 
    158.62499246571716, 158.74999245977997, 158.87499245384279, 
    158.99999244790561, 159.12499244196843, 159.24999243603125, 
    159.37499243009407, 159.49999242415689, 159.6249924182197, 
    159.74999241228252, 159.87499240634534, 159.99999240040816, 
    160.12499239447098, 160.2499923885338, 160.37499238259662, 
    160.49999237665943, 160.62499237072225, 160.74999236478507, 
    160.87499235884789, 160.99999235291071, 161.12499234697353, 
    161.24999234103635, 161.37499233509917, 161.49999232916198, 
    161.6249923232248, 161.74999231728762, 161.87499231135044, 
    161.99999230541326, 162.12499229947608, 162.2499922935389, 
    162.37499228760171, 162.49999228166453, 162.62499227572735, 
    162.74999226979017, 162.87499226385299, 162.99999225791581, 
    163.12499225197863, 163.24999224604144, 163.37499224010426, 
    163.49999223416708, 163.6249922282299, 163.74999222229272, 
    163.87499221635554, 163.99999221041836, 164.12499220448117, 
    164.24999219854399, 164.37499219260681, 164.49999218666963, 
    164.62499218073245, 164.74999217479527, 164.87499216885809, 
    164.9999921629209, 165.12499215698372, 165.24999215104654, 
    165.37499214510936, 165.49999213917218, 165.624992133235, 
    165.74999212729782, 165.87499212136063, 165.99999211542345, 
    166.12499210948627, 166.24999210354909, 166.37499209761191, 
    166.49999209167473, 166.62499208573755, 166.74999207980036, 
    166.87499207386318, 166.999992067926, 167.12499206198882, 
    167.24999205605164, 167.37499205011446, 167.49999204417728, 
    167.62499203824009, 167.74999203230291, 167.87499202636573, 
    167.99999202042855, 168.12499201449137, 168.24999200855419, 
    168.37499200261701, 168.49999199667982, 168.62499199074264, 
    168.74999198480546, 168.87499197886828, 168.9999919729311, 
    169.12499196699392, 169.24999196105674, 169.37499195511955, 
    169.49999194918237, 169.62499194324519, 169.74999193730801, 
    169.87499193137083, 169.99999192543365, 170.12499191949649, 
    170.24999191355931, 170.37499190762213, 170.49999190168495, 
    170.62499189574777, 170.74999188981059, 170.87499188387341, 
    170.99999187793622, 171.12499187199904, 171.24999186606186, 
    171.37499186012468, 171.4999918541875, 171.62499184825032, 
    171.74999184231314, 171.87499183637595, 171.99999183043877, 
    172.12499182450159, 172.24999181856441, 172.37499181262723, 
    172.49999180669005, 172.62499180075287, 172.74999179481568, 
    172.8749917888785, 172.99999178294132, 173.12499177700414, 
    173.24999177106696, 173.37499176512978, 173.4999917591926, 
    173.62499175325542, 173.74999174731823, 173.87499174138105, 
    173.99999173544387, 174.12499172950669, 174.24999172356951, 
    174.37499171763233, 174.49999171169515, 174.62499170575796, 
    174.74999169982078, 174.8749916938836, 174.99999168794642, 
    175.12499168200924, 175.24999167607206, 175.37499167013488, 
    175.49999166419769, 175.62499165826051, 175.74999165232333, 
    175.87499164638615, 175.99999164044897, 176.12499163451179, 
    176.24999162857461, 176.37499162263742, 176.49999161670024, 
    176.62499161076306, 176.74999160482588, 176.8749915988887, 
    176.99999159295152, 177.12499158701434, 177.24999158107715, 
    177.37499157513997, 177.49999156920279, 177.62499156326561, 
    177.74999155732843, 177.87499155139125, 177.99999154545407, 
    178.12499153951688, 178.2499915335797, 178.37499152764252, 
    178.49999152170534, 178.62499151576816, 178.74999150983098, 
    178.8749915038938, 178.99999149795661, 179.12499149201943, 
    179.24999148608225, 179.37499148014507, 179.49999147420789, 
    179.62499146827071, 179.74999146233353, 179.87499145639634, 
    179.99999145045916, 180.12499144452198, 180.2499914385848, 
    180.37499143264762, 180.49999142671044, 180.62499142077326, 
    180.74999141483607, 180.87499140889889, 180.99999140296171, 
    181.12499139702453, 181.24999139108735, 181.37499138515017, 
    181.49999137921299, 181.6249913732758, 181.74999136733862, 
    181.87499136140144, 181.99999135546426, 182.12499134952708, 
    182.2499913435899, 182.37499133765272, 182.49999133171553, 
    182.62499132577835, 182.7499913198412, 182.87499131390402, 
    182.99999130796684, 183.12499130202966, 183.24999129609247, 
    183.37499129015529, 183.49999128421811, 183.62499127828093, 
    183.74999127234375, 183.87499126640657, 183.99999126046939, 
    184.1249912545322, 184.24999124859502, 184.37499124265784, 
    184.49999123672066, 184.62499123078348, 184.7499912248463, 
    184.87499121890912, 184.99999121297193, 185.12499120703475, 
    185.24999120109757, 185.37499119516039, 185.49999118922321, 
    185.62499118328603, 185.74999117734885, 185.87499117141166, 
    185.99999116547448, 186.1249911595373, 186.24999115360012, 
    186.37499114766294, 186.49999114172576, 186.62499113578858, 
    186.7499911298514, 186.87499112391421, 186.99999111797703, 
    187.12499111203985, 187.24999110610267, 187.37499110016549, 
    187.49999109422831, 187.62499108829113, 187.74999108235394, 
    187.87499107641676, 187.99999107047958, 188.1249910645424, 
    188.24999105860522, 188.37499105266804, 188.49999104673086, 
    188.62499104079367, 188.74999103485649, 188.87499102891931, 
    188.99999102298213, 189.12499101704495, 189.24999101110777, 
    189.37499100517059, 189.4999909992334, 189.62499099329622, 
    189.74999098735904, 189.87499098142186, 189.99999097548468, 
    190.1249909695475, 190.24999096361032, 190.37499095767313, 
    190.49999095173595, 190.62499094579877, 190.74999093986159, 
    190.87499093392441, 190.99999092798723, 191.12499092205005, 
    191.24999091611286, 191.37499091017568, 191.4999909042385, 
    191.62499089830132, 191.74999089236414, 191.87499088642696, 
    191.99999088048978, 192.12499087455259, 192.24999086861541, 
    192.37499086267823, 192.49999085674105, 192.62499085080387, 
    192.74999084486669, 192.87499083892951, 192.99999083299232, 
    193.12499082705514, 193.24999082111796, 193.37499081518078, 
    193.4999908092436, 193.62499080330642, 193.74999079736924, 
    193.87499079143205, 193.99999078549487, 194.12499077955769, 
    194.24999077362051, 194.37499076768333, 194.49999076174615, 
    194.62499075580897, 194.74999074987178, 194.8749907439346, 
    194.99999073799742, 195.12499073206024, 195.24999072612306, 
    195.37499072018591, 195.49999071424872, 195.62499070831154, 
    195.74999070237436, 195.87499069643718, 195.9999906905, 
    196.12499068456282, 196.24999067862564, 196.37499067268845, 
    196.49999066675127, 196.62499066081409, 196.74999065487691, 
    196.87499064893973, 196.99999064300255, 197.12499063706537, 
    197.24999063112818, 197.374990625191, 197.49999061925382, 
    197.62499061331664, 197.74999060737946, 197.87499060144228, 
    197.9999905955051, 198.12499058956791, 198.24999058363073, 
    198.37499057769355, 198.49999057175637, 198.62499056581919, 
    198.74999055988201, 198.87499055394483, 198.99999054800764, 
    199.12499054207046, 199.24999053613328, 199.3749905301961, 
    199.49999052425892, 199.62499051832174, 199.74999051238456, 
    199.87499050644738, 199.99999050051019, 200.12499049457301, 
    200.24999048863583, 200.37499048269865, 200.49999047676147, 
    200.62499047082429, 200.74999046488711, 200.87499045894992, 
    200.99999045301274, 201.12499044707556, 201.24999044113838, 
    201.3749904352012, 201.49999042926402, 201.62499042332684, 
    201.74999041738965, 201.87499041145247, 201.99999040551529, 
    202.12499039957811, 202.24999039364093, 202.37499038770375, 
    202.49999038176657, 202.62499037582938, 202.7499903698922, 
    202.87499036395502, 202.99999035801784, 203.12499035208066, 
    203.24999034614348, 203.3749903402063, 203.49999033426911, 
    203.62499032833193, 203.74999032239475, 203.87499031645757, 
    203.99999031052039, 204.12499030458321, 204.24999029864603, 
    204.37499029270884, 204.49999028677166, 204.62499028083448, 
    204.7499902748973, 204.87499026896012, 204.99999026302294, 
    205.12499025708576, 205.24999025114857, 205.37499024521139, 
    205.49999023927421, 205.62499023333703, 205.74999022739985, 
    205.87499022146267, 205.99999021552549, 206.1249902095883, 
    206.24999020365112, 206.37499019771394, 206.49999019177676, 
    206.62499018583958, 206.7499901799024, 206.87499017396522, 
    206.99999016802803, 207.12499016209085, 207.24999015615367, 
    207.37499015021649, 207.49999014427931, 207.62499013834213, 
    207.74999013240495, 207.87499012646779, 207.99999012053061, 
    208.12499011459343, 208.24999010865625, 208.37499010271907, 
    208.49999009678189, 208.6249900908447, 208.74999008490752, 
    208.87499007897034, 208.99999007303316, 209.12499006709598, 
    209.2499900611588, 209.37499005522162, 209.49999004928443, 
    209.62499004334725, 209.74999003741007, 209.87499003147289, 
    209.99999002553571, 210.12499001959853, 210.24999001366135, 
    210.37499000772416, 210.49999000178698, 210.6249899958498, 
    210.74998998991262, 210.87498998397544, 210.99998997803826, 
    211.12498997210108, 211.24998996616389, 211.37498996022671, 
    211.49998995428953, 211.62498994835235, 211.74998994241517, 
    211.87498993647799, 211.99998993054081, 212.12498992460363, 
    212.24998991866644, 212.37498991272926, 212.49998990679208, 
    212.6249899008549, 212.74998989491772, 212.87498988898054, 
    212.99998988304336, 213.12498987710617, 213.24998987116899, 
    213.37498986523181, 213.49998985929463, 213.62498985335745, 
    213.74998984742027, 213.87498984148309, 213.9999898355459, 
    214.12498982960872, 214.24998982367154, 214.37498981773436, 
    214.49998981179718, 214.62498980586, 214.74998979992282, 
    214.87498979398563, 214.99998978804845, 215.12498978211127, 
    215.24998977617409, 215.37498977023691, 215.49998976429973, 
    215.62498975836255, 215.74998975242536, 215.87498974648818, 
    215.999989740551, 216.12498973461382, 216.24998972867664, 
    216.37498972273946, 216.49998971680228, 216.62498971086509, 
    216.74998970492791, 216.87498969899073, 216.99998969305355, 
    217.12498968711637, 217.24998968117919, 217.37498967524201, 
    217.49998966930482, 217.62498966336764, 217.74998965743046, 
    217.87498965149328, 217.9999896455561, 218.12498963961892, 
    218.24998963368174, 218.37498962774455, 218.49998962180737, 
    218.62498961587019, 218.74998960993301, 218.87498960399583, 
    218.99998959805865, 219.12498959212147, 219.24998958618428, 
    219.3749895802471, 219.49998957430992, 219.62498956837274, 
    219.74998956243556, 219.87498955649838, 219.9999895505612, 
    220.12498954462401, 220.24998953868683, 220.37498953274965, 
    220.4999895268125, 220.62498952087532, 220.74998951493814, 
    220.87498950900095, 220.99998950306377, 221.12498949712659, 
    221.24998949118941, 221.37498948525223, 221.49998947931505, 
    221.62498947337787, 221.74998946744068, 221.8749894615035, 
    221.99998945556632, 222.12498944962914, 222.24998944369196, 
    222.37498943775478, 222.4999894318176, 222.62498942588041, 
    222.74998941994323, 222.87498941400605, 222.99998940806887, 
    223.12498940213169, 223.24998939619451, 223.37498939025733, 
    223.49998938432014, 223.62498937838296, 223.74998937244578, 
    223.8749893665086, 223.99998936057142, 224.12498935463424, 
    224.24998934869706, 224.37498934275987, 224.49998933682269, 
    224.62498933088551, 224.74998932494833, 224.87498931901115, 
    224.99998931307397, 225.12498930713679, 225.24998930119961, 
    225.37498929526242, 225.49998928932524, 225.62498928338806, 
    225.74998927745088, 225.8749892715137, 225.99998926557652, 
    226.12498925963934, 226.24998925370215, 226.37498924776497, 
    226.49998924182779, 226.62498923589061, 226.74998922995343, 
    226.87498922401625, 226.99998921807907, 227.12498921214188, 
    227.2499892062047, 227.37498920026752, 227.49998919433034, 
    227.62498918839316, 227.74998918245598, 227.8749891765188, 
    227.99998917058161, 228.12498916464443, 228.24998915870725, 
    228.37498915277007, 228.49998914683289, 228.62498914089571, 
    228.74998913495853, 228.87498912902134, 228.99998912308416, 
    229.12498911714698, 229.2499891112098, 229.37498910527262, 
    229.49998909933544, 229.62498909339826, 229.74998908746107, 
    229.87498908152389, 229.99998907558671, 230.12498906964953, 
    230.24998906371235, 230.37498905777517, 230.49998905183799, 
    230.6249890459008, 230.74998903996362, 230.87498903402644, 
    230.99998902808926, 231.12498902215208, 231.2499890162149, 
    231.37498901027772, 231.49998900434053, 231.62498899840335, 
    231.74998899246617, 231.87498898652899, 231.99998898059181, 
    232.12498897465463, 232.24998896871745, 232.37498896278026, 
    232.49998895684308, 232.6249889509059, 232.74998894496872, 
    232.87498893903154, 232.99998893309436, 233.1249889271572, 
    233.24998892122002, 233.37498891528284, 233.49998890934566, 
    233.62498890340848, 233.7499888974713, 233.87498889153412, 
    233.99998888559693, 234.12498887965975, 234.24998887372257, 
    234.37498886778539, 234.49998886184821, 234.62498885591103, 
    234.74998884997385, 234.87498884403666, 234.99998883809948, 
    235.1249888321623, 235.24998882622512, 235.37498882028794, 
    235.49998881435076, 235.62498880841358, 235.74998880247639, 
    235.87498879653921, 235.99998879060203, 236.12498878466485, 
    236.24998877872767, 236.37498877279049, 236.49998876685331, 
    236.62498876091612, 236.74998875497894, 236.87498874904176, 
    236.99998874310458, 237.1249887371674, 237.24998873123022, 
    237.37498872529304, 237.49998871935585, 237.62498871341867, 
    237.74998870748149, 237.87498870154431, 237.99998869560713, 
    238.12498868966995, 238.24998868373277, 238.37498867779559, 
    238.4999886718584, 238.62498866592122, 238.74998865998404, 
    238.87498865404686, 238.99998864810968, 239.1249886421725, 
    239.24998863623532, 239.37498863029813, 239.49998862436095, 
    239.62498861842377, 239.74998861248659, 239.87498860654941, 
    239.99998860061223, 240.12498859467505, 240.24998858873786, 
    240.37498858280068, 240.4999885768635, 240.62498857092632, 
    240.74998856498914, 240.87498855905196, 240.99998855311478, 
    241.12498854717759, 241.24998854124041, 241.37498853530323, 
    241.49998852936605, 241.62498852342887, 241.74998851749169, 
    241.87498851155451, 241.99998850561732, 242.12498849968014, 
    242.24998849374296, 242.37498848780578, 242.4999884818686, 
    242.62498847593142, 242.74998846999424, 242.87498846405705, 
    242.99998845811987, 243.12498845218269, 243.24998844624551, 
    243.37498844030833, 243.49998843437115, 243.62498842843397, 
    243.74998842249678, 243.8749884165596, 243.99998841062242, 
    244.12498840468524, 244.24998839874806, 244.37498839281088, 
    244.4999883868737, 244.62498838093651, 244.74998837499933, 
    244.87498836906215, 244.99998836312497, 245.12498835718779, 
    245.24998835125061, 245.37498834531343, 245.49998833937624, 
    245.62498833343906, 245.74998832750191, 245.87498832156473, 
    245.99998831562755, 246.12498830969037, 246.24998830375318, 
    246.374988297816, 246.49998829187882, 246.62498828594164, 
    246.74998828000446, 246.87498827406728, 246.9999882681301, 
    247.12498826219291, 247.24998825625573, 247.37498825031855, 
    247.49998824438137, 247.62498823844419, 247.74998823250701, 
    247.87498822656983, 247.99998822063264, 248.12498821469546, 
    248.24998820875828, 248.3749882028211, 248.49998819688392, 
    248.62498819094674, 248.74998818500956, 248.87498817907237, 
    248.99998817313519, 249.12498816719801, 249.24998816126083, 
    249.37498815532365, 249.49998814938647, 249.62498814344929, 
    249.7499881375121, 249.87498813157492 ;

 angular_frequency = 0, 0.78539812609303905, 1.5707962521860781, 
    2.3561943782791168, 3.1415925043721562, 3.9269906304651951, 
    4.7123887565582336, 5.4977868826512735, 6.2831850087443124, 
    7.0685831348373505, 7.8539812609303903, 8.6393793870234301, 
    9.4247775131164673, 10.210175639209508, 10.995573765302547, 
    11.780971891395586, 12.566370017488625, 13.351768143581664, 
    14.137166269674701, 14.922564395767742, 15.707962521860781, 
    16.493360647953818, 17.27875877404686, 18.064156900139899, 
    18.849555026232935, 19.634953152325977, 20.420351278419016, 
    21.205749404512055, 21.991147530605094, 22.776545656698129, 
    23.561943782791172, 24.347341908884211, 25.13274003497725, 
    25.918138161070285, 26.703536287163328, 27.488934413256366, 
    28.274332539349402, 29.059730665442444, 29.845128791535483, 
    30.630526917628519, 31.415925043721561, 32.2013231698146, 
    32.986721295907635, 33.772119422000678, 34.55751754809372, 
    35.342915674186756, 36.128313800279798, 36.913711926372834, 
    37.699110052465869, 38.484508178558912, 39.269906304651954, 
    40.055304430744989, 40.840702556838032, 41.626100682931067, 
    42.41149880902411, 43.196896935117145, 43.982295061210188, 
    44.767693187303223, 45.553091313396258, 46.338489439489301, 
    47.123887565582343, 47.909285691675379, 48.694683817768421, 
    49.480081943861457, 50.265480069954499, 51.050878196047535, 
    51.83627632214057, 52.62167444823362, 53.407072574326655, 
    54.19247070041969, 54.977868826512733, 55.763266952605768, 
    56.548665078698804, 57.334063204791853, 58.119461330884889, 
    58.904859456977931, 59.690257583070967, 60.475655709164002, 
    61.261053835257037, 62.046451961350087, 62.831850087443122, 
    63.617248213536165, 64.4026463396292, 65.188044465722243, 
    65.973442591815271, 66.758840717908313, 67.544238844001356, 
    68.329636970094398, 69.115035096187441, 69.900433222280469, 
    70.685831348373512, 71.47122947446654, 72.256627600559597, 
    73.042025726652639, 73.827423852745667, 74.61282197883871, 
    75.398220104931738, 76.183618231024781, 76.969016357117823, 
    77.754414483210866, 78.539812609303908, 79.325210735396936, 
    80.110608861489979, 80.896006987583021, 81.681405113676064, 
    82.466803239769106, 83.252201365862135, 84.037599491955177, 
    84.82299761804822, 85.608395744141248, 86.39379387023429, 
    87.179191996327333, 87.964590122420375, 88.749988248513418, 
    89.535386374606446, 90.320784500699489, 91.106182626792517, 
    91.891580752885574, 92.676978878978602, 93.462377005071644, 
    94.247775131164687, 95.033173257257715, 95.818571383350758, 
    96.6039695094438, 97.389367635536843, 98.174765761629885, 
    98.960163887722914, 99.745562013815956, 100.530960139909, 
    101.31635826600203, 102.10175639209507, 102.8871545181881, 
    103.67255264428114, 104.4579507703742, 105.24334889646724, 
    106.02874702256028, 106.81414514865331, 107.59954327474635, 
    108.38494140083938, 109.17033952693242, 109.95573765302547, 
    110.74113577911849, 111.52653390521154, 112.31193203130458, 
    113.09733015739761, 113.88272828349066, 114.66812640958371, 
    115.45352453567675, 116.23892266176978, 117.02432078786282, 
    117.80971891395586, 118.59511704004889, 119.38051516614193, 
    120.16591329223496, 120.951311418328, 121.73670954442105, 
    122.52210767051407, 123.30750579660712, 124.09290392270017, 
    124.87830204879322, 125.66370017488624, 126.44909830097929, 
    127.23449642707233, 128.01989455316536, 128.8052926792584, 
    129.59069080535144, 130.37608893144449, 131.1614870575375, 
    131.94688518363054, 132.73228330972358, 133.51768143581663, 
    134.3030795619097, 135.08847768800271, 135.87387581409575, 
    136.6592739401888, 137.44467206628184, 138.23007019237488, 
    139.0154683184679, 139.80086644456094, 140.58626457065398, 
    141.37166269674702, 142.15706082284007, 142.94245894893308, 
    143.72785707502615, 144.51325520111919, 145.29865332721224, 
    146.08405145330528, 146.86944957939829, 147.65484770549133, 
    148.44024583158438, 149.22564395767742, 150.01104208377046, 
    150.79644020986348, 151.58183833595652, 152.36723646204956, 
    153.1526345881426, 153.93803271423565, 154.72343084032869, 
    155.50882896642173, 156.29422709251477, 157.07962521860782, 
    157.86502334470086, 158.65042147079387, 159.43581959688692, 
    160.22121772297996, 161.006615849073, 161.79201397516604, 
    162.57741210125906, 163.36281022735213, 164.14820835344517, 
    164.93360647953821, 165.71900460563123, 166.50440273172427, 
    167.28980085781731, 168.07519898391035, 168.8605971100034, 
    169.64599523609644, 170.43139336218945, 171.2167914882825, 
    172.00218961437554, 172.78758774046858, 173.57298586656162, 
    174.35838399265467, 175.14378211874771, 175.92918024484075, 
    176.71457837093379, 177.49997649702684, 178.28537462311985, 
    179.07077274921289, 179.85617087530593, 180.64156900139898, 
    181.42696712749202, 182.21236525358503, 182.99776337967808, 
    183.78316150577115, 184.56855963186419, 185.3539577579572, 
    186.13935588405025, 186.92475401014329, 187.71015213623633, 
    188.49555026232937, 189.28094838842242, 190.06634651451543, 
    190.85174464060847, 191.63714276670152, 192.42254089279456, 
    193.2079390188876, 193.99333714498064, 194.77873527107369, 
    195.56413339716673, 196.34953152325977, 197.13492964935278, 
    197.92032777544583, 198.70572590153887, 199.49112402763191, 
    200.27652215372495, 201.061920279818, 201.84731840591101, 
    202.63271653200405, 203.4181146580971, 204.20351278419014, 
    204.98891091028318, 205.7743090363762, 206.55970716246924, 
    207.34510528856228, 208.13050341465535, 208.91590154074839, 
    209.70129966684144, 210.48669779293448, 211.27209591902752, 
    212.05749404512056, 212.84289217121358, 213.62829029730662, 
    214.41368842339966, 215.1990865494927, 215.98448467558575, 
    216.76988280167876, 217.5552809277718, 218.34067905386485, 
    219.12607717995789, 219.91147530605093, 220.69687343214397, 
    221.48227155823699, 222.26766968433003, 223.05306781042307, 
    223.83846593651612, 224.62386406260916, 225.40926218870217, 
    226.19466031479521, 226.98005844088826, 227.76545656698133, 
    228.55085469307437, 229.33625281916741, 230.12165094526046, 
    230.9070490713535, 231.69244719744654, 232.47784532353955, 
    233.2632434496326, 234.04864157572564, 234.83403970181868, 
    235.61943782791172, 236.40483595400474, 237.19023408009778, 
    237.97563220619082, 238.76103033228387, 239.54642845837691, 
    240.33182658446992, 241.11722471056297, 241.90262283665601, 
    242.68802096274905, 243.47341908884209, 244.25881721493514, 
    245.04421534102815, 245.82961346712119, 246.61501159321423, 
    247.40040971930731, 248.18580784540035, 248.97120597149339, 
    249.75660409758643, 250.54200222367948, 251.32740034977249, 
    252.11279847586553, 252.89819660195857, 253.68359472805162, 
    254.46899285414466, 255.2543909802377, 256.03978910633072, 
    256.82518723242379, 257.6105853585168, 258.39598348460981, 
    259.18138161070289, 259.9667797367959, 260.75217786288897, 
    261.53757598898198, 262.322974115075, 263.10837224116807, 
    263.89377036726108, 264.67916849335415, 265.46456661944717, 
    266.24996474554018, 267.03536287163325, 267.82076099772632, 
    268.6061591238194, 269.39155724991241, 270.17695537600542, 
    270.96235350209849, 271.74775162819151, 272.53314975428458, 
    273.31854788037759, 274.10394600647061, 274.88934413256368, 
    275.67474225865669, 276.46014038474976, 277.24553851084278, 
    278.03093663693579, 278.81633476302886, 279.60173288912188, 
    280.38713101521495, 281.17252914130796, 281.95792726740098, 
    282.74332539349405, 283.52872351958706, 284.31412164568013, 
    285.09951977177315, 285.88491789786616, 286.67031602395923, 
    287.4557141500523, 288.24111227614532, 289.02651040223839, 
    289.8119085283314, 290.59730665442447, 291.38270478051749, 
    292.16810290661056, 292.95350103270357, 293.73889915879658, 
    294.52429728488966, 295.30969541098267, 296.09509353707574, 
    296.88049166316875, 297.66588978926177, 298.45128791535484, 
    299.23668604144785, 300.02208416754092, 300.80748229363394, 
    301.59288041972695, 302.37827854582002, 303.16367667191304, 
    303.94907479800611, 304.73447292409912, 305.51987105019214, 
    306.30526917628521, 307.09066730237828, 307.87606542847129, 
    308.66146355456436, 309.44686168065738, 310.23225980675045, 
    311.01765793284346, 311.80305605893653, 312.58845418502955, 
    313.37385231112256, 314.15925043721563, 314.94464856330865, 
    315.73004668940172, 316.51544481549473, 317.30084294158775, 
    318.08624106768082, 318.87163919377383, 319.6570373198669, 
    320.44243544595992, 321.22783357205293, 322.013231698146, 
    322.79862982423901, 323.58402795033209, 324.3694260764251, 
    325.15482420251811, 325.94022232861118, 326.72562045470426, 
    327.51101858079727, 328.29641670689034, 329.08181483298335, 
    329.86721295907643, 330.65261108516944, 331.43800921126245, 
    332.22340733735552, 333.00880546344854, 333.79420358954161, 
    334.57960171563462, 335.36499984172769, 336.15039796782071, 
    336.93579609391372, 337.72119422000679, 338.50659234609981, 
    339.29199047219288, 340.07738859828589, 340.86278672437891, 
    341.64818485047198, 342.43358297656499, 343.21898110265806, 
    344.00437922875108, 344.78977735484409, 345.57517548093716, 
    346.36057360703023, 347.14597173312325, 347.93136985921632, 
    348.71676798530933, 349.5021661114024, 350.28756423749542, 
    351.07296236358843, 351.8583604896815, 352.64375861577452, 
    353.42915674186759, 354.2145548679606, 354.99995299405367, 
    355.78535112014669, 356.5707492462397, 357.35614737233277, 
    358.14154549842578, 358.92694362451886, 359.71234175061187, 
    360.49773987670488, 361.28313800279795, 362.06853612889097, 
    362.85393425498404, 363.63933238107705, 364.42473050717007, 
    365.21012863326314, 365.99552675935615, 366.78092488544922, 
    367.56632301154229, 368.35172113763531, 369.13711926372838, 
    369.92251738982139, 370.70791551591441, 371.49331364200748, 
    372.27871176810049, 373.06410989419356, 373.84950802028658, 
    374.63490614637959, 375.42030427247266, 376.20570239856568, 
    376.99110052465875, 377.77649865075176, 378.56189677684483, 
    379.34729490293785, 380.13269302903086, 380.91809115512393, 
    381.70348928121695, 382.48888740731002, 383.27428553340303, 
    384.05968365949605, 384.84508178558912, 385.63047991168213, 
    386.4158780377752, 387.20127616386827, 387.98667428996129, 
    388.77207241605436, 389.55747054214737, 390.34286866824038, 
    391.12826679433346, 391.91366492042647, 392.69906304651954, 
    393.48446117261255, 394.26985929870557, 395.05525742479864, 
    395.84065555089165, 396.62605367698472, 397.41145180307774, 
    398.19684992917081, 398.98224805526382, 399.76764618135684, 
    400.55304430744991, 401.33844243354292, 402.12384055963599, 
    402.90923868572901, 403.69463681182202, 404.48003493791509, 
    405.26543306400811, 406.05083119010118, 406.83622931619419, 
    407.62162744228721, 408.40702556838028, 409.19242369447329, 
    409.97782182056636, 410.76321994665938, 411.54861807275239, 
    412.33401619884546, 413.11941432493848, 413.90481245103155, 
    414.69021057712456, 415.47560870321757, 416.2610068293107, 
    417.04640495540377, 417.83180308149679, 418.61720120758986, 
    419.40259933368287, 420.18799745977594, 420.97339558586896, 
    421.75879371196197, 422.54419183805504, 423.32958996414806, 
    424.11498809024113, 424.90038621633414, 425.68578434242716, 
    426.47118246852023, 427.25658059461324, 428.04197872070631, 
    428.82737684679932, 429.61277497289234, 430.39817309898541, 
    431.18357122507842, 431.96896935117149, 432.75436747726451, 
    433.53976560335752, 434.32516372945059, 435.11056185554361, 
    435.89595998163668, 436.68135810772969, 437.46675623382271, 
    438.25215435991578, 439.03755248600879, 439.82295061210186, 
    440.60834873819488, 441.39374686428795, 442.17914499038096, 
    442.96454311647398, 443.74994124256705, 444.53533936866006, 
    445.32073749475313, 446.10613562084615, 446.89153374693916, 
    447.67693187303223, 448.46232999912525, 449.24772812521832, 
    450.03312625131133, 450.81852437740434, 451.60392250349742, 
    452.38932062959043, 453.1747187556835, 453.96011688177651, 
    454.74551500786953, 455.53091313396266, 456.31631126005573, 
    457.10170938614874, 457.88710751224181, 458.67250563833483, 
    459.45790376442784, 460.24330189052091, 461.02870001661393, 
    461.814098142707, 462.59949626880001, 463.38489439489308, 
    464.1702925209861, 464.95569064707911, 465.74108877317218, 
    466.52648689926519, 467.31188502535827, 468.09728315145128, 
    468.88268127754429, 469.66807940363736, 470.45347752973038, 
    471.23887565582345, 472.02427378191646, 472.80967190800948, 
    473.59507003410255, 474.38046816019556, 475.16586628628863, 
    475.95126441238165, 476.73666253847466, 477.52206066456773, 
    478.30745879066075, 479.09285691675382, 479.87825504284683, 
    480.66365316893985, 481.44905129503292, 482.23444942112593, 
    483.019847547219, 483.80524567331202, 484.59064379940509, 
    485.3760419254981, 486.16144005159111, 486.94683817768419, 
    487.7322363037772, 488.51763442987027, 489.30303255596328, 
    490.0884306820563, 490.87382880814937, 491.65922693424238, 
    492.44462506033545, 493.23002318642847, 494.01542131252148, 
    494.80081943861461, 495.58621756470768, 496.3716156908007, 
    497.15701381689377, 497.94241194298678, 498.72781006907979, 
    499.51320819517287, 500.29860632126588, 501.08400444735895, 
    501.86940257345196, 502.65480069954498, 503.44019882563805, 
    504.22559695173106, 505.01099507782413, 505.79639320391715, 
    506.58179133001022, 507.36718945610323, 508.15258758219625, 
    508.93798570828932, 509.72338383438233, 510.5087819604754, 
    511.29418008656842, 512.07957821266143, 512.86497633875445, 
    513.65037446484757, 514.43577259094059, 515.2211707170336, 
    516.00656884312662, 516.79196696921963, 517.57736509531276, 
    518.36276322140577, 519.14816134749879, 519.9335594735918, 
    520.71895759968481, 521.50435572577794, 522.28975385187096, 
    523.07515197796397, 523.86055010405698, 524.64594823015, 
    525.43134635624313, 526.21674448233614, 527.00214260842915, 
    527.78754073452217, 528.57293886061518, 529.35833698670831, 
    530.14373511280132, 530.92913323889434, 531.71453136498735, 
    532.49992949108037, 533.28532761717349, 534.07072574326651, 
    534.85612386935964, 535.64152199545265, 536.42692012154566, 
    537.21231824763879, 537.99771637373181, 538.78311449982482, 
    539.56851262591783, 540.35391075201085, 541.13930887810398, 
    541.92470700419699, 542.71010513029, 543.49550325638302, 
    544.28090138247603, 545.06629950856916, 545.85169763466217, 
    546.63709576075519, 547.4224938868482, 548.20789201294122, 
    548.99329013903434, 549.77868826512736, 550.56408639122037, 
    551.34948451731339, 552.1348826434064, 552.92028076949953, 
    553.70567889559254, 554.49107702168556, 555.27647514777857, 
    556.06187327387158, 556.84727139996471, 557.63266952605773, 
    558.41806765215074, 559.20346577824375, 559.98886390433677, 
    560.7742620304299, 561.55966015652291, 562.34505828261592, 
    563.13045640870894, 563.91585453480195, 564.70125266089508, 
    565.48665078698809, 566.27204891308111, 567.05744703917412, 
    567.84284516526714, 568.62824329136026, 569.41364141745328, 
    570.19903954354629, 570.98443766963931, 571.76983579573232, 
    572.55523392182545, 573.34063204791846, 574.12603017401159, 
    574.9114283001046, 575.69682642619762, 576.48222455229063, 
    577.26762267838376, 578.05302080447677, 578.83841893056979, 
    579.6238170566628, 580.40921518275593, 581.19461330884894, 
    581.98001143494196, 582.76540956103497, 583.55080768712799, 
    584.33620581322111, 585.12160393931413, 585.90700206540714, 
    586.69240019150016, 587.47779831759317, 588.2631964436863, 
    589.04859456977931, 589.83399269587233, 590.61939082196534, 
    591.40478894805835, 592.19018707415148, 592.9755852002445, 
    593.76098332633751, 594.54638145243052, 595.33177957852354, 
    596.11717770461667, 596.90257583070968, 597.68797395680269, 
    598.47337208289571, 599.25877020898872, 600.04416833508185, 
    600.82956646117486, 601.61496458726788, 602.40036271336089, 
    603.18576083945391, 603.97115896554703, 604.75655709164005, 
    605.54195521773306, 606.32735334382608, 607.11275146991909, 
    607.89814959601222, 608.68354772210523, 609.46894584819825, 
    610.25434397429126, 611.03974210038427, 611.8251402264774, 
    612.61053835257042, 613.39593647866343, 614.18133460475656, 
    614.96673273084957, 615.75213085694259, 616.53752898303571, 
    617.32292710912873, 618.10832523522174, 618.89372336131476, 
    619.67912148740777, 620.4645196135009, 621.24991773959391, 
    622.03531586568693, 622.82071399177994, 623.60611211787307, 
    624.39151024396608, 625.1769083700591, 625.96230649615211, 
    626.74770462224512, 627.53310274833825, 628.31850087443127, 
    629.10389900052428, 629.88929712661729, 630.67469525271031, 
    631.46009337880344, 632.24549150489645, 633.03088963098946, 
    633.81628775708248, 634.60168588317549, 635.38708400926862, 
    636.17248213536163, 636.95788026145465, 637.74327838754766, 
    638.52867651364068, 639.3140746397338, 640.09947276582682, 
    640.88487089191983, 641.67026901801285, 642.45566714410586, 
    643.24106527019899, 644.026463396292, 644.81186152238502, 
    645.59725964847803, 646.38265777457104, 647.16805590066417, 
    647.95345402675719, 648.7388521528502, 649.52425027894321, 
    650.30964840503623, 651.09504653112936, 651.88044465722237, 
    652.66584278331538, 653.45124090940851, 654.23663903550153, 
    655.02203716159454, 655.80743528768767, 656.59283341378068, 
    657.3782315398737, 658.16362966596671, 658.94902779205972, 
    659.73442591815285, 660.51982404424587, 661.30522217033888, 
    662.09062029643189, 662.87601842252491, 663.66141654861804, 
    664.44681467471105, 665.23221280080406, 666.01761092689708, 
    666.80300905299021, 667.58840717908322, 668.37380530517623, 
    669.15920343126925, 669.94460155736226, 670.72999968345539, 
    671.5153978095484, 672.30079593564142, 673.08619406173443, 
    673.87159218782745, 674.65699031392057, 675.44238844001359, 
    676.2277865661066, 677.01318469219962, 677.79858281829263, 
    678.58398094438576, 679.36937907047877, 680.15477719657179, 
    680.9401753226648, 681.72557344875781, 682.51097157485094, 
    683.29636970094396, 684.08176782703697, 684.86716595312998, 
    685.652564079223, 686.43796220531613, 687.22336033140914, 
    688.00875845750215, 688.79415658359517, 689.57955470968818, 
    690.36495283578131, 691.15035096187432, 691.93574908796734, 
    692.72114721406047, 693.50654534015348, 694.29194346624649, 
    695.07734159233962, 695.86273971843264, 696.64813784452565, 
    697.43353597061866, 698.21893409671168, 699.00433222280481, 
    699.78973034889782, 700.57512847499083, 701.36052660108385, 
    702.14592472717686, 702.93132285326999, 703.716720979363, 
    704.50211910545602, 705.28751723154903, 706.07291535764205, 
    706.85831348373517, 707.64371160982819, 708.4291097359212, 
    709.21450786201422, 709.99990598810734, 710.78530411420036, 
    711.57070224029337, 712.35610036638639, 713.1414984924794, 
    713.92689661857253, 714.71229474466554, 715.49769287075856, 
    716.28309099685157, 717.06848912294458, 717.85388724903771, 
    718.63928537513073, 719.42468350122374, 720.21008162731675, 
    720.99547975340977, 721.7808778795029, 722.56627600559591, 
    723.35167413168892, 724.13707225778194, 724.92247038387495, 
    725.70786850996808, 726.49326663606109, 727.27866476215411, 
    728.06406288824712, 728.84946101434014, 729.63485914043326, 
    730.42025726652628, 731.20565539261929, 731.99105351871231, 
    732.77645164480543, 733.56184977089845, 734.34724789699158, 
    735.13264602308459, 735.9180441491776, 736.70344227527062, 
    737.48884040136363, 738.27423852745676, 739.05963665354977, 
    739.84503477964279, 740.6304329057358, 741.41583103182882, 
    742.20122915792194, 742.98662728401496, 743.77202541010797, 
    744.55742353620099, 745.342821662294, 746.12821978838713, 
    746.91361791448014, 747.69901604057316, 748.48441416666617, 
    749.26981229275918, 750.05521041885231, 750.84060854494533, 
    751.62600667103834, 752.41140479713135, 753.19680292322448, 
    753.9822010493175, 754.76759917541051, 755.55299730150352, 
    756.33839542759654, 757.12379355368967, 757.90919167978268, 
    758.69458980587569, 759.47998793196871, 760.26538605806172, 
    761.05078418415485, 761.83618231024786, 762.62158043634088, 
    763.40697856243389, 764.19237668852691, 764.97777481462003, 
    765.76317294071305, 766.54857106680606, 767.33396919289908, 
    768.11936731899209, 768.90476544508522, 769.69016357117823, 
    770.47556169727125, 771.26095982336426, 772.04635794945739, 
    772.8317560755504, 773.61715420164353, 774.40255232773654, 
    775.18795045382956, 775.97334857992257, 776.75874670601559, 
    777.54414483210871, 778.32954295820173, 779.11494108429474, 
    779.90033921038776, 780.68573733648077, 781.4711354625739, 
    782.25653358866691, 783.04193171475993, 783.82732984085294, 
    784.61272796694595, 785.39812609303908, 786.1835242191321, 
    786.96892234522511, 787.75432047131812, 788.53971859741114, 
    789.32511672350427, 790.11051484959728, 790.89591297569029, 
    791.68131110178331, 792.46670922787632, 793.25210735396945, 
    794.03750548006246, 794.82290360615548, 795.60830173224849, 
    796.39369985834162, 797.17909798443463, 797.96449611052765, 
    798.74989423662066, 799.53529236271368, 800.3206904888068, 
    801.10608861489982, 801.89148674099283, 802.67688486708585, 
    803.46228299317886, 804.24768111927199, 805.033079245365, 
    805.81847737145802, 806.60387549755103, 807.38927362364404, 
    808.17467174973717, 808.96006987583019, 809.7454680019232, 
    810.53086612801621, 811.31626425410923, 812.10166238020236, 
    812.88706050629537, 813.67245863238838, 814.4578567584814, 
    815.24325488457441, 816.02865301066754, 816.81405113676055, 
    817.59944926285357, 818.38484738894658, 819.1702455150396, 
    819.95564364113272, 820.74104176722574, 821.52643989331875, 
    822.31183801941177, 823.09723614550478, 823.88263427159791, 
    824.66803239769092, 825.45343052378394, 826.23882864987695, 
    827.02422677596996, 827.80962490206309, 828.59502302815611, 
    829.38042115424912, 830.16581928034213, 830.95121740643515, 
    831.73661553252839, 832.5220136586214, 833.30741178471453, 
    834.09280991080755, 834.87820803690056, 835.66360616299357, 
    836.44900428908659, 837.23440241517972, 838.01980054127273, 
    838.80519866736574, 839.59059679345876, 840.37599491955189, 
    841.1613930456449, 841.94679117173791, 842.73218929783093, 
    843.51758742392394, 844.30298555001707, 845.08838367611008, 
    845.8737818022031, 846.65917992829611, 847.44457805438913, 
    848.22997618048225, 849.01537430657527, 849.80077243266828, 
    850.5861705587613, 851.37156868485431, 852.15696681094744, 
    852.94236493704045, 853.72776306313347, 854.51316118922648, 
    855.29855931531949, 856.08395744141262, 856.86935556750564, 
    857.65475369359865, 858.44015181969166, 859.22554994578468, 
    860.01094807187781, 860.79634619797082, 861.58174432406383, 
    862.36714245015685, 863.15254057624986, 863.93793870234299, 
    864.723336828436, 865.50873495452902, 866.29413308062203, 
    867.07953120671505, 867.86492933280817, 868.65032745890119, 
    869.4357255849942, 870.22112371108722, 871.00652183718023, 
    871.79191996327336, 872.57731808936637, 873.36271621545939, 
    874.1481143415524, 874.93351246764541, 875.71891059373854, 
    876.50430871983156, 877.28970684592457, 878.07510497201758, 
    878.86050309811071, 879.64590122420373, 880.43129935029674, 
    881.21669747638975, 882.00209560248277, 882.7874937285759, 
    883.57289185466891, 884.35828998076192, 885.14368810685494, 
    885.92908623294795, 886.71448435904108, 887.49988248513409, 
    888.28528061122711, 889.07067873732012, 889.85607686341314, 
    890.64147498950626, 891.42687311559928, 892.21227124169229, 
    892.99766936778531, 893.78306749387832, 894.56846561997145, 
    895.35386374606446, 896.13926187215748, 896.92465999825049, 
    897.7100581243435, 898.49545625043663, 899.28085437652965, 
    900.06625250262266, 900.85165062871567, 901.63704875480869, 
    902.42244688090182, 903.20784500699483, 903.99324313308784, 
    904.77864125918086, 905.56403938527387, 906.349437511367, 
    907.13483563746001, 907.92023376355303, 908.70563188964604, 
    909.49103001573906, 910.27642814183218, 911.06182626792531, 
    911.84722439401844, 912.63262252011145, 913.41802064620447, 
    914.20341877229748, 914.9888168983905, 915.77421502448362, 
    916.55961315057664, 917.34501127666965, 918.13040940276267, 
    918.91580752885568, 919.70120565494881, 920.48660378104182, 
    921.27200190713484, 922.05740003322785, 922.84279815932086, 
    923.62819628541399, 924.41359441150701, 925.19899253760002, 
    925.98439066369303, 926.76978878978616, 927.55518691587918, 
    928.34058504197219, 929.1259831680652, 929.91138129415822, 
    930.69677942025135, 931.48217754634436, 932.26757567243737, 
    933.05297379853039, 933.8383719246234, 934.62377005071653, 
    935.40916817680954, 936.19456630290256, 936.97996442899557, 
    937.76536255508859, 938.55076068118171, 939.33615880727473, 
    940.12155693336774, 940.90695505946076, 941.69235318555377, 
    942.4777513116469, 943.26314943773991, 944.04854756383293, 
    944.83394568992594, 945.61934381601895, 946.40474194211208, 
    947.1901400682051, 947.97553819429811, 948.76093632039112, 
    949.54633444648414, 950.33173257257727, 951.11713069867028, 
    951.90252882476329, 952.68792695085631, 953.47332507694932, 
    954.25872320304245, 955.04412132913546, 955.82951945522848, 
    956.61491758132149, 957.40031570741451, 958.18571383350763, 
    958.97111195960065, 959.75651008569366, 960.54190821178668, 
    961.32730633787969, 962.11270446397282, 962.89810259006583, 
    963.68350071615885, 964.46889884225186, 965.25429696834499, 
    966.039695094438, 966.82509322053102, 967.61049134662403, 
    968.39588947271704, 969.18128759881017, 969.96668572490319, 
    970.7520838509962, 971.53748197708921, 972.32288010318223, 
    973.10827822927536, 973.89367635536837, 974.67907448146138, 
    975.4644726075544, 976.24987073364741, 977.03526885974054, 
    977.82066698583355, 978.60606511192657, 979.39146323801958, 
    980.1768613641126, 980.96225949020572, 981.74765761629874, 
    982.53305574239175, 983.31845386848477, 984.10385199457778, 
    984.88925012067091, 985.67464824676392, 986.46004637285694, 
    987.24544449894995, 988.03084262504296, 988.81624075113609, 
    989.60163887722922, 990.38703700332235, 991.17243512941536, 
    991.95783325550838, 992.74323138160139, 993.5286295076944, 
    994.31402763378753, 995.09942575988055, 995.88482388597356, 
    996.67022201206657, 997.45562013815959, 998.24101826425272, 
    999.02641639034573, 999.81181451643874, 1000.5972126425318, 
    1001.3826107686248, 1002.1680088947179, 1002.9534070208109, 
    1003.7388051469039, 1004.5242032729969, 1005.30960139909, 
    1006.0949995251831, 1006.8803976512761, 1007.6657957773691, 
    1008.4511939034621, 1009.2365920295553, 1010.0219901556483, 
    1010.8073882817413, 1011.5927864078343, 1012.3781845339273, 
    1013.1635826600204, 1013.9489807861135, 1014.7343789122065, 
    1015.5197770382995, 1016.3051751643925, 1017.0905732904856, 
    1017.8759714165786, 1018.6613695426717, 1019.4467676687647, 
    1020.2321657948577, 1021.0175639209508, 1021.8029620470438, 
    1022.5883601731368, 1023.3737582992298, 1024.1591564253229, 
    1024.9445545514159, 1025.7299526775089, 1026.5153508036019, 
    1027.3007489296951, 1028.0861470557882, 1028.8715451818812, 
    1029.6569433079742, 1030.4423414340672, 1031.2277395601602, 
    1032.0131376862532, 1032.7985358123462, 1033.5839339384393, 
    1034.3693320645325, 1035.1547301906255, 1035.9401283167185, 
    1036.7255264428115, 1037.5109245689046, 1038.2963226949976, 
    1039.0817208210906, 1039.8671189471836, 1040.6525170732766, 
    1041.4379151993696, 1042.2233133254629, 1043.0087114515559, 
    1043.7941095776489, 1044.5795077037419, 1045.3649058298349, 
    1046.1503039559279, 1046.935702082021, 1047.721100208114, 
    1048.506498334207, 1049.2918964603, 1050.0772945863932, 
    1050.8626927124863, 1051.6480908385793, 1052.4334889646723, 
    1053.2188870907653, 1054.0042852168583, 1054.7896833429513, 
    1055.5750814690443, 1056.3604795951373, 1057.1458777212304, 
    1057.9312758473236, 1058.7166739734166, 1059.5020720995096, 
    1060.2874702256026, 1061.0728683516957, 1061.8582664777887, 
    1062.6436646038817, 1063.4290627299747, 1064.2144608560677, 
    1064.9998589821607, 1065.785257108254, 1066.570655234347, 
    1067.35605336044, 1068.141451486533, 1068.9268496126263, 
    1069.7122477387193, 1070.4976458648123, 1071.2830439909053, 
    1072.0684421169983, 1072.8538402430913, 1073.6392383691843, 
    1074.4246364952776, 1075.2100346213706, 1075.9954327474636, 
    1076.7808308735566, 1077.5662289996496, 1078.3516271257427, 
    1079.1370252518357, 1079.9224233779287, 1080.7078215040217, 
    1081.4932196301147, 1082.278617756208, 1083.064015882301, 
    1083.849414008394, 1084.634812134487, 1085.42021026058, 
    1086.205608386673, 1086.991006512766, 1087.776404638859, 
    1088.5618027649521, 1089.3472008910451, 1090.1325990171383, 
    1090.9179971432313, 1091.7033952693243, 1092.4887933954174, 
    1093.2741915215104, 1094.0595896476034, 1094.8449877736964, 
    1095.6303858997894, 1096.4157840258824, 1097.2011821519754, 
    1097.9865802780687, 1098.7719784041617, 1099.5573765302547, 
    1100.3427746563477, 1101.1281727824407, 1101.9135709085338, 
    1102.6989690346268, 1103.4843671607198, 1104.2697652868128, 
    1105.0551634129058, 1105.8405615389991, 1106.6259596650921, 
    1107.4113577911851, 1108.1967559172781, 1108.9821540433711, 
    1109.7675521694641, 1110.5529502955571, 1111.3383484216502, 
    1112.1237465477432, 1112.9091446738362, 1113.6945427999294, 
    1114.4799409260224, 1115.2653390521155, 1116.0507371782085, 
    1116.8361353043015, 1117.6215334303945, 1118.4069315564875, 
    1119.1923296825805, 1119.9777278086735, 1120.7631259347668, 
    1121.5485240608598, 1122.3339221869528, 1123.1193203130458, 
    1123.9047184391388, 1124.6901165652318, 1125.4755146913249, 
    1126.2609128174179, 1127.0463109435109, 1127.8317090696039, 
    1128.6171071956971, 1129.4025053217902, 1130.1879034478832, 
    1130.9733015739762, 1131.7586997000692, 1132.5440978261622, 
    1133.3294959522552, 1134.1148940783482, 1134.9002922044413, 
    1135.6856903305343, 1136.4710884566275, 1137.2564865827205, 
    1138.0418847088135, 1138.8272828349066, 1139.6126809609996, 
    1140.3980790870926, 1141.1834772131856, 1141.9688753392786, 
    1142.7542734653716, 1143.5396715914646, 1144.3250697175579, 
    1145.1104678436509, 1145.8958659697439, 1146.6812640958369, 
    1147.4666622219299, 1148.2520603480232, 1149.0374584741162, 
    1149.8228566002092, 1150.6082547263022, 1151.3936528523952, 
    1152.1790509784882, 1152.9644491045813, 1153.7498472306745, 
    1154.5352453567675, 1155.3206434828605, 1156.1060416089535, 
    1156.8914397350466, 1157.6768378611396, 1158.4622359872326, 
    1159.2476341133256, 1160.0330322394186, 1160.8184303655119, 
    1161.6038284916049, 1162.3892266176979, 1163.1746247437909, 
    1163.9600228698839, 1164.7454209959769, 1165.5308191220699, 
    1166.316217248163, 1167.101615374256, 1167.887013500349, 
    1168.6724116264422, 1169.4578097525352, 1170.2432078786283, 
    1171.0286060047213, 1171.8140041308143, 1172.5994022569073, 
    1173.3848003830003, 1174.1701985090933, 1174.9555966351863, 
    1175.7409947612794, 1176.5263928873726, 1177.3117910134656, 
    1178.0971891395586, 1178.8825872656516, 1179.6679853917447, 
    1180.4533835178377, 1181.2387816439307, 1182.0241797700237, 
    1182.8095778961167, 1183.5949760222097, 1184.380374148303, 
    1185.165772274396, 1185.951170400489, 1186.736568526582, 
    1187.521966652675, 1188.307364778768, 1189.092762904861, 
    1189.8781610309541, 1190.6635591570471, 1191.4489572831401, 
    1192.2343554092333, 1193.0197535353263, 1193.8051516614194, 
    1194.5905497875124, 1195.3759479136054, 1196.1613460396984, 
    1196.9467441657914, 1197.7321422918844, 1198.5175404179774, 
    1199.3029385440707, 1200.0883366701637, 1200.8737347962567, 
    1201.6591329223497, 1202.4445310484427, 1203.2299291745358, 
    1204.0153273006288, 1204.8007254267218, 1205.5861235528148, 
    1206.3715216789078, 1207.1569198050011, 1207.9423179310941, 
    1208.7277160571871, 1209.5131141832801, 1210.2985123093731, 
    1211.0839104354661, 1211.8693085615591, 1212.6547066876522, 
    1213.4401048137452, 1214.2255029398382, 1215.0109010659314, 
    1215.7962991920244, 1216.5816973181174, 1217.3670954442105, 
    1218.1524935703035, 1218.9378916963965, 1219.7232898224895, 
    1220.5086879485825, 1221.2940860746755, 1222.0794842007685, 
    1222.8648823268618, 1223.6502804529548, 1224.4356785790478, 
    1225.2210767051408, 1226.0064748312338, 1226.7918729573269, 
    1227.5772710834201, 1228.3626692095131, 1229.1480673356061, 
    1229.9334654616991, 1230.7188635877922, 1231.5042617138852, 
    1232.2896598399784, 1233.0750579660714, 1233.8604560921644, 
    1234.6458542182575, 1235.4312523443505, 1236.2166504704435, 
    1237.0020485965365, 1237.7874467226295, 1238.5728448487225, 
    1239.3582429748155, 1240.1436411009088, 1240.9290392270018, 
    1241.7144373530948, 1242.4998354791878, 1243.2852336052808, 
    1244.0706317313739, 1244.8560298574669, 1245.6414279835599, 
    1246.4268261096529, 1247.2122242357461, 1247.9976223618391, 
    1248.7830204879322, 1249.5684186140252, 1250.3538167401182, 
    1251.1392148662112, 1251.9246129923042, 1252.7100111183972, 
    1253.4954092444902, 1254.2808073705833, 1255.0662054966765, 
    1255.8516036227695, 1256.6370017488625, 1257.4223998749555, 
    1258.2077980010486, 1258.9931961271416, 1259.7785942532346, 
    1260.5639923793276, 1261.3493905054206, 1262.1347886315136, 
    1262.9201867576069, 1263.7055848836999, 1264.4909830097929, 
    1265.2763811358859, 1266.0617792619789, 1266.8471773880719, 
    1267.632575514165, 1268.417973640258, 1269.203371766351, 
    1269.988769892444, 1270.7741680185372, 1271.5595661446303, 
    1272.3449642707233, 1273.1303623968163, 1273.9157605229093, 
    1274.7011586490023, 1275.4865567750953, 1276.2719549011883, 
    1277.0573530272814, 1277.8427511533744, 1278.6281492794676, 
    1279.4135474055606, 1280.1989455316536, 1280.9843436577466, 
    1281.7697417838397, 1282.5551399099327, 1283.3405380360257, 
    1284.1259361621187, 1284.9113342882117, 1285.696732414305, 
    1286.482130540398, 1287.267528666491, 1288.052926792584, 
    1288.838324918677, 1289.62372304477, 1290.409121170863, 
    1291.1945192969561, 1291.9799174230491, 1292.7653155491421, 
    1293.5507136752353, 1294.3361118013283, 1295.1215099274214, 
    1295.9069080535144, 1296.6923061796074, 1297.4777043057004, 
    1298.2631024317934, 1299.0485005578864, 1299.8338986839794, 
    1300.6192968100725, 1301.4046949361657, 1302.1900930622587, 
    1302.9754911883517, 1303.7608893144447, 1304.5462874405378, 
    1305.3316855666308, 1306.117083692724, 1306.902481818817, 
    1307.68787994491, 1308.4732780710031, 1309.2586761970961, 
    1310.0440743231891, 1310.8294724492823, 1311.6148705753753, 
    1312.4002687014683, 1313.1856668275614, 1313.9710649536544, 
    1314.7564630797474, 1315.5418612058404, 1316.3272593319334, 
    1317.1126574580264, 1317.8980555841194, 1318.6834537102127, 
    1319.4688518363057, 1320.2542499623987, 1321.0396480884917, 
    1321.8250462145847, 1322.6104443406778, 1323.3958424667708, 
    1324.1812405928638, 1324.9666387189568, 1325.7520368450498, 
    1326.5374349711431, 1327.3228330972361, 1328.1082312233291, 
    1328.8936293494221, 1329.6790274755151, 1330.4644256016081, 
    1331.2498237277011, 1332.0352218537942, 1332.8206199798872, 
    1333.6060181059804, 1334.3914162320734, 1335.1768143581664, 
    1335.9622124842595, 1336.7476106103525, 1337.5330087364455, 
    1338.3184068625385, 1339.1038049886315, 1339.8892031147245, 
    1340.6746012408175, 1341.4599993669108, 1342.2453974930038, 
    1343.0307956190968, 1343.8161937451898, 1344.6015918712828, 
    1345.3869899973758, 1346.1723881234689, 1346.9577862495619, 
    1347.7431843756549, 1348.5285825017479, 1349.3139806278411, 
    1350.0993787539342, 1350.8847768800272, 1351.6701750061202, 
    1352.4555731322132, 1353.2409712583062, 1354.0263693843992, 
    1354.8117675104922, 1355.5971656365853, 1356.3825637626783, 
    1357.1679618887715, 1357.9533600148645, 1358.7387581409575, 
    1359.5241562670506, 1360.3095543931436, 1361.0949525192366, 
    1361.8803506453296, 1362.6657487714226, 1363.4511468975156, 
    1364.2365450236086, 1365.0219431497019, 1365.8073412757949, 
    1366.5927394018879, 1367.3781375279809, 1368.1635356540739, 
    1368.948933780167, 1369.73433190626, 1370.519730032353, 
    1371.305128158446, 1372.0905262845392, 1372.8759244106323, 
    1373.6613225367253, 1374.4467206628183, 1375.2321187889113, 
    1376.0175169150043, 1376.8029150410973, 1377.5883131671903, 
    1378.3737112932833, 1379.1591094193764, 1379.9445075454696, 
    1380.7299056715626, 1381.5153037976556, 1382.3007019237486, 
    1383.0861000498417, 1383.8714981759347, 1384.6568963020277, 
    1385.4422944281209, 1386.2276925542139, 1387.013090680307, 
    1387.7984888064, 1388.583886932493, 1389.3692850585862, 
    1390.1546831846792, 1390.9400813107723, 1391.7254794368653, 
    1392.5108775629583, 1393.2962756890513, 1394.0816738151443, 
    1394.8670719412373, 1395.6524700673303, 1396.4378681934234, 
    1397.2232663195166, 1398.0086644456096, 1398.7940625717026, 
    1399.5794606977956, 1400.3648588238887, 1401.1502569499817, 
    1401.9356550760747, 1402.7210532021677, 1403.5064513282607, 
    1404.2918494543537, 1405.077247580447, 1405.86264570654, 
    1406.648043832633, 1407.433441958726, 1408.218840084819, 
    1409.004238210912, 1409.789636337005, 1410.5750344630981, 
    1411.3604325891911, 1412.1458307152841, 1412.9312288413773, 
    1413.7166269674703, 1414.5020250935634, 1415.2874232196564, 
    1416.0728213457494, 1416.8582194718424, 1417.6436175979354, 
    1418.4290157240284, 1419.2144138501214, 1419.9998119762147, 
    1420.7852101023077, 1421.5706082284007, 1422.3560063544937, 
    1423.1414044805867, 1423.9268026066798, 1424.7122007327728, 
    1425.4975988588658, 1426.2829969849588, 1427.0683951110518, 
    1427.8537932371451, 1428.6391913632381, 1429.4245894893311, 
    1430.2099876154241, 1430.9953857415171, 1431.7807838676101, 
    1432.5661819937031, 1433.3515801197962, 1434.1369782458892, 
    1434.9223763719822, 1435.7077744980754, 1436.4931726241684, 
    1437.2785707502615, 1438.0639688763545, 1438.8493670024475, 
    1439.6347651285405, 1440.4201632546335, 1441.2055613807265, 
    1441.9909595068195, 1442.7763576329125, 1443.5617557590058, 
    1444.3471538850988, 1445.1325520111918, 1445.9179501372848, 
    1446.7033482633778, 1447.4887463894709, 1448.2741445155639, 
    1449.0595426416569, 1449.8449407677499, 1450.6303388938429, 
    1451.4157370199362, 1452.2011351460292, 1452.9865332721222, 
    1453.7719313982152, 1454.5573295243082, 1455.3427276504012, 
    1456.1281257764942, 1456.9135239025873, 1457.6989220286803, 
    1458.4843201547735, 1459.2697182808665, 1460.0551164069595, 
    1460.8405145330526, 1461.6259126591456, 1462.4113107852386, 
    1463.1967089113316, 1463.9821070374246, 1464.7675051635179, 
    1465.5529032896109, 1466.3383014157039, 1467.1236995417969, 
    1467.9090976678901, 1468.6944957939832, 1469.4798939200762, 
    1470.2652920461692, 1471.0506901722622, 1471.8360882983552, 
    1472.6214864244482, 1473.4068845505412, 1474.1922826766342, 
    1474.9776808027273, 1475.7630789288205, 1476.5484770549135, 
    1477.3338751810065, 1478.1192733070995, 1478.9046714331926, 
    1479.6900695592856, 1480.4754676853786, 1481.2608658114716, 
    1482.0462639375646, 1482.8316620636576, 1483.6170601897509, 
    1484.4024583158439, 1485.1878564419369, 1485.9732545680299, 
    1486.7586526941229, 1487.5440508202159, 1488.329448946309, 
    1489.114847072402, 1489.900245198495, 1490.685643324588, 
    1491.4710414506812, 1492.2564395767743, 1493.0418377028673, 
    1493.8272358289603, 1494.6126339550533, 1495.3980320811463, 
    1496.1834302072393, 1496.9688283333323, 1497.7542264594254, 
    1498.5396245855184, 1499.3250227116116, 1500.1104208377046, 
    1500.8958189637976, 1501.6812170898907, 1502.4666152159837, 
    1503.2520133420767, 1504.0374114681697, 1504.8228095942627, 
    1505.6082077203557, 1506.393605846449, 1507.179003972542, 
    1507.964402098635, 1508.749800224728, 1509.535198350821, 
    1510.320596476914, 1511.105994603007, 1511.8913927291001, 
    1512.6767908551931, 1513.4621889812861, 1514.2475871073793, 
    1515.0329852334723, 1515.8183833595654, 1516.6037814856584, 
    1517.3891796117514, 1518.1745777378444, 1518.9599758639374, 
    1519.7453739900304, 1520.5307721161234, 1521.3161702422165, 
    1522.1015683683097, 1522.8869664944027, 1523.6723646204957, 
    1524.4577627465887, 1525.2431608726818, 1526.0285589987748, 
    1526.8139571248678, 1527.5993552509608, 1528.3847533770538, 
    1529.1701515031468, 1529.9555496292401, 1530.7409477553331, 
    1531.5263458814261, 1532.3117440075191, 1533.0971421336121, 
    1533.8825402597051, 1534.6679383857982, 1535.4533365118912, 
    1536.2387346379842, 1537.0241327640772, 1537.8095308901704, 
    1538.5949290162634, 1539.3803271423565, 1540.1657252684495, 
    1540.9511233945425, 1541.7365215206355, 1542.5219196467285, 
    1543.3073177728215, 1544.0927158989148, 1544.8781140250078, 
    1545.6635121511008, 1546.448910277194, 1547.2343084032871, 
    1548.0197065293801, 1548.8051046554731, 1549.5905027815661, 
    1550.3759009076591, 1551.1612990337521, 1551.9466971598451, 
    1552.7320952859382, 1553.5174934120312, 1554.3028915381244, 
    1555.0882896642174, 1555.8736877903104, 1556.6590859164035, 
    1557.4444840424965, 1558.2298821685895, 1559.0152802946825, 
    1559.8006784207755, 1560.5860765468685, 1561.3714746729615, 
    1562.1568727990548, 1562.9422709251478, 1563.7276690512408, 
    1564.5130671773338, 1565.2984653034268, 1566.0838634295199, 
    1566.8692615556129, 1567.6546596817059, 1568.4400578077989, 
    1569.2254559338919, 1570.0108540599851 ;

 time_resolution = 1, 0.99991675375292488, 0.99966705658901767, 
    0.99925103320562614, 0.99866889131634384, 0.99792092147817368, 
    0.99700749684983814, 0.99592907288151777, 0.99468618693637945, 
    0.99327945784433536, 0.99170958538854992, 0.98997734972529206, 
    0.98808361073780659, 0.98602930732495309, 0.98381545662543546, 
    0.98144315317852182, 0.97891356802222151, 0.97622794772996091, 
    0.97338761338686686, 0.97039395950683527, 0.96724845289162609, 
    0.96395263143329235, 0.96050810286131172, 0.95691654343584853, 
    0.95317969658863388, 0.94929937151300448, 0.94527744170469785, 
    0.94111584345504895, 0.9368165742982858, 0.93238169141466387, 
    0.92781330999122824, 0.92311360154202649, 0.91828479218964265, 
    0.91332916090995009, 0.9082490377420207, 0.90304680196515497, 
    0.89772488024502661, 0.89228574475095934, 0.88673191124637774, 
    0.88106593715448989, 0.87529041960128018, 0.86940799343790043, 
    0.86342132924456017, 0.85733313131802569, 0.85114613564484032, 
    0.84486310786238106, 0.83848684120986927, 0.83202015447144329, 
    0.82546588991340175, 0.81882691121771323, 0.81210610141387485, 
    0.80530636081119467, 0.79843060493354723, 0.79148176245863899, 
    0.78446277316379398, 0.77737658588024849, 0.77022615645791348, 
    0.7630144457425373, 0.75574441756716615, 0.74841903675977051, 
    0.74104126716886298, 0.73361406970890297, 0.72614040042723604, 
    0.7186232085942782, 0.7110654348186104, 0.70347000918860203, 
    0.69583984944213528, 0.68817785916595409, 0.68048692602610872, 
    0.67276992003091896, 0.66502969182782024, 0.65726907103540844, 
    0.64949086461193872, 0.64169785526148138, 0.63389279987887437, 
    0.6260784280345626, 0.61825744050034426, 0.61043250781699399, 
    0.60260626890466762, 0.59478132971693154, 0.58696026193920425, 
    0.57914560173232743, 0.57133984852193231, 0.5635454638341969, 
    0.55576487017853382, 0.54800044997768227, 0.5402545445456215, 
    0.53252945311365796, 0.52482743190497994, 0.51715069325790985, 
    0.50950140479803174, 0.50188168865930449, 0.49429362075421823, 
    0.48673923009299064, 0.4792204981517475, 0.47173935828956981, 
    0.4642976952142418, 0.45689734449647368, 0.44954009213232698, 
    0.44222767415351411, 0.43496177628519561, 0.42774403365084873, 
    0.42057603052373571, 0.41345930012445026, 0.40639532446398102, 
    0.39938553423168055, 0.3924313087274956, 0.38553397583776661, 
    0.37869481205387034, 0.37191504253293983, 0.36519584119986381, 
    0.3585383308897313, 0.35194358352985716, 0.34541262036049158, 
    0.33894641219329241, 0.33254587970660876, 0.32621189377660009, 
    0.31994527584319327, 0.31374679830985747, 0.30761718497615781, 
    0.30155711150202835, 0.2955672059026942, 0.28964804907315034, 
    0.28380017534109975, 0.27802407304723692, 0.27232018515175638, 
    0.26668890986595567, 0.26113060130779969, 0.25564557018030526, 
    0.25023408447160428, 0.24489637017554142, 0.23963261203166256, 
    0.23444295428345352, 0.22932750145368941, 0.22428631913576066, 
    0.21931943479984944, 0.21442683861283396, 0.20960848427081133, 
    0.20486428984313473, 0.20019413862687666, 0.19559788001063907, 
    0.19107533034664609, 0.18662627383006897, 0.18225046338455034, 
    0.17794762155290841, 0.17371744139202355, 0.16955958737092303, 
    0.16547369627110486, 0.16145937808815697, 0.15751621693375248, 
    0.15364377193712017, 0.14984157814511539, 0.14610914742003633, 
    0.14244596933435594, 0.13885151206156271, 0.13532522326232954, 
    0.13186653096525258, 0.12847484444142976, 0.12514955507217193, 
    0.1218900372091677, 0.11869564902644644, 0.11556573336351357, 
    0.11249961855905596, 0.1094966192746424, 0.10655603730787237, 
    0.10367716239445035, 0.10085927299869167, 0.098101637091991795, 
    0.095403512918815894, 0.092764149749795285, 0.090182788621539431, 
    0.087658663062801345, 0.08519099980665816, 0.082779019488394612, 
    0.080421937328802345, 0.078118963802633223, 0.07586930529196742, 
    0.073672164724284325, 0.071526742195044846, 0.069432235574618528, 
    0.067387841099411941, 0.065392753947075805, 0.063446168795691593, 
    0.061547280366858914, 0.0596952839526253, 0.057889375926221856, 
    0.056128754236586344, 0.054412618886674924, 0.052740172395583096, 
    0.051110620244512857, 0.049523171306642133, 0.047977038260968177, 
    0.046471437990212611, 0.045005591962892916, 0.043578726599678215, 
    0.042190073624162723, 0.040838870398203185, 0.039524360241980583, 
    0.038245792738957687, 0.037002424025917018, 0.035793517068273731, 
    0.034618341920869974, 0.033476175974465887, 0.032366304188152492, 
    0.03128801930792053, 0.030240622071626946, 0.02922342140060899, 
    0.028235734578202453, 0.027276887415426679, 0.026346214404106057, 
    0.02544305885770164, 0.024566773040132134, 0.023716718282867637, 
    0.02289226509058297, 0.022092793235661112, 0.021317691841839709, 
    0.020566359457295652, 0.019838204117465379, 0.019132643397898889, 
    0.018449104457447081, 0.017787024072082099, 0.017145848659650856, 
    0.016525034295861073, 0.015924046721799066, 0.01534236134327681, 
    0.014779463222305084, 0.01423484706098713, 0.0137080171781256, 
    0.013198487478832991, 0.012705781417433226, 0.012229431953938852, 
    0.011768981504385601, 0.01132398188530182, 0.010893994252587585, 
    0.010478589035073427, 0.010077345863025101, 0.0096898534918564167, 
    0.009315709721307389, 0.008954521310340597, 0.0086059038880038057, 
    0.0082694818605018039, 0.0079448883147153551, 0.0076317649184002691, 
    0.007329761817293892, 0.0070385375293512235, 0.0067577588363272869, 
    0.0064871006729169444, 0.0062262460136575945, 0.0059748857577948764, 
    0.0057327186123054003, 0.0054994509732652665, 0.0052747968057471843, 
    0.0050584775224232744, 0.0048502218610450435, 0.0046497657609662736, 
    0.0044568522388687814, 0.0042712312638455057, 0.0040926596319895633, 
    0.0039209008406324982, 0.0037557249623692735, 0.003596908519002072, 
    0.0034442343555296192, 0.0032974915143032515, 0.0031564751094657314, 
    0.0030209862017835237, 0.0028908316739780816, 0.0027658241066567286, 
    0.0026457816549385338, 0.0025305279258658951, 0.0024198918566875564, 
    0.0023137075940941961, 0.0022118143744830699, 0.0021140564053236748, 
    0.0020202827476919652, 0.0019303472000364609, 0.0018441081832352528, 
    0.0017614286269989191, 0.0016821758576703553, 0.0016062214874686584, 
    0.0015334413052204604, 0.0014637151686184512, 0.0013969268980432922, 
    0.0013329641719817585, 0.0012717184240705491, 0.0012130847417921053, 
    0.0011569617668456241, 0.0011032515972135167, 0.0010518596909407057, 
    0.0010026947716413773, 0.0009556687357451637, 0.0009106965614922364, 
    0.0008676962196842989, 0.00082658858619618269, 0.00078729735625051418, 
    0.00074974896045579579, 0.00071387248260622684, 0.0006795995792396722, 
    0.00064686440094832286, 0.00061560351543492873, 0.00058575583230575934, 
    0.00055726252958996551, 0.0005300669819735044, 0.00050411469073444789, 
    0.00047935321536517238, 0.00045573210686574231, 0.00043320284269163803, 
    0.00041171876333796406, 0.00039123501054125003, 0.00037170846707908206, 
    0.00035309769814695298, 0.00033536289429094898, 0.00031846581587419804, 
    0.00030236973905436017, 0.00028703940324885494, 0.00027244096006403119, 
    0.00025854192366398004, 0.00024531112255433534, 0.00023271865275600889, 
    0.00022073583234352777, 0.00020933515732239605, 0.00019849025881965395, 
    0.00018817586156170095, 0.00017836774361326783, 0.00016904269735139269, 
    0.00016017849164817207, 0.00015175383523607526, 0.00014374834122963243, 
    0.00013614249277734937, 0.00012891760981782467, 0.0001220558169141256, 
    0.00011554001214066392, 0.00010935383699694832, 0.00010348164732282148, 
    9.790848518997702e-05, 9.2620051744813733e-05, 8.7602680977935573e-05, 
    8.2843314395877014e-05, 7.8329476570942569e-05, 7.404925154533836e-05, 
    6.9991260066120956e-05, 6.61446376278003e-05, 6.2499013299799493e-05, 
    5.9044489316328693e-05, 5.5771621406587196e-05, 5.2671399843603896e-05, 
    4.9735231190389055e-05, 4.6954920722477425e-05, 4.4322655506325462e-05, 
    4.183098811343531e-05, 3.9472820950474326e-05, 3.7241391186069904e-05, 
    3.5130256255369515e-05, 3.3133279923859878e-05, 3.1244618892359799e-05, 
    2.9458709925502941e-05, 2.7770257486446217e-05, 2.6174221860942907e-05, 
    2.4665807754331997e-05, 2.3240453345400792e-05, 2.1893819781478871e-05, 
    2.0621781099527582e-05, 1.942041455838027e-05, 1.8285991367688525e-05, 
    1.7214967799513047e-05, 1.6203976668888393e-05, 1.5249819170066887e-05, 
    1.4349457055523914e-05, 1.3500005145178367e-05, 1.2698724153642407e-05, 
    1.1943013823678244e-05, 1.1230406354388338e-05, 1.0558560113015445e-05, 
    9.9252536195665702e-06, 9.3283797938123319e-06, 8.7659404545376421e-06, 
    8.2360410612435781e-06, 7.736885688813765e-06, 7.2667722259661368e-06, 
    6.8240877886137903e-06, 6.4073043395508461e-06, 6.014974506169662e-06, 
    5.6457275881941253e-06, 5.2982657476897594e-06, 4.9713603738782881e-06, 
    4.6638486155443322e-06, 4.3746300740772478e-06, 4.1026636504370383e-06, 
    3.8469645395753751e-06, 3.606601366075707e-06, 3.3806934550054076e-06, 
    3.1684082321930318e-06, 2.9689587483597384e-06, 2.7816013217421972e-06, 
    2.6056332940467401e-06, 2.4403908947716518e-06, 2.2852472091242498e-06, 
    2.1396102449448874e-06, 2.0029210942282258e-06, 1.8746521850058626e-06, 
    1.7543056195219337e-06, 1.6414115947954368e-06, 1.5355269018202386e-06, 
    1.4362334998051141e-06, 1.3431371620030934e-06, 1.2558661898206589e-06, 
    1.1740701920344971e-06, 1.0974189260750627e-06, 1.0256011984639103e-06, 
    9.583238216144357e-07, 8.9531062432404011e-07, 8.3630151340005453e-07, 
    7.8105158397145208e-07, 7.2933027614459443e-07, 6.8092057576290194e-07, 
    6.3561825712866362e-07, 5.9323116563956299e-07, 5.5357853838312788e-07, 
    5.1649036081982564e-07, 4.818067577691535e-07, 4.4937741699385225e-07, 
    4.1906104375458906e-07, 3.9072484478189732e-07, 3.6424404018334264e-07, 
    3.3950140187237134e-07, 3.1638681717090884e-07, 2.9479687630062572e-07, 
    2.7463448253819391e-07, 2.5580848386752073e-07, 2.3823332501740592e-07, 
    2.218287188259813e-07, 2.0651933592407639e-07, 1.9223451177821351e-07, 
    1.7890797018033705e-07, 1.6647756231588587e-07, 1.5488502058421426e-07, 
    1.4407572638604539e-07, 1.3399849113136725e-07, 1.2460534975830227e-07, 
    1.1585136608882496e-07, 1.076944493810197e-07, 1.0009518146981182e-07, 
    9.3016653918855098e-08, 8.6424314635640398e-08, 8.0285823429839801e-08, 
    7.4570916021608181e-08, 6.9251276031973824e-08, 6.4300414511675431e-08, 
    5.9693556587889473e-08, 5.5407534830241756e-08, 5.1420688958437593e-08, 
    4.7712771533725037e-08, 4.4264859295368824e-08, 4.1059269821305348e-08, 
    3.807948320929376e-08, 3.5310068491153959e-08, 3.2736614508158425e-08, 
    3.0345664990357822e-08, 2.8124657596573327e-08, 2.6061866685066238e-08, 
    2.4146349597477644e-08, 2.2367896250588297e-08, 2.071698184178441e-08, 
    1.9184722484875223e-08, 1.7762833603110601e-08, 1.6443590915915592e-08, 
    1.5219793865032302e-08, 1.4084731334442359e-08, 1.3032149526679467e-08, 
    1.2056221865930904e-08, 1.1151520805715546e-08, 1.031299142590714e-08, 
    9.5359267104892126e-09, 8.8159444036842143e-09, 8.1489653480167704e-09, 
    7.5311932134706844e-09, 6.9590955321894435e-09, 6.4293859581736618e-09, 
    5.9390076761536918e-09, 5.48511788828415e-09, 5.0650733115218025e-09, 
    4.676416622533177e-09, 4.3168637907376198e-09, 3.9842922436392019e-09, 
    3.6767298119508266e-09, 3.3923444051707052e-09, 3.1294343712521135e-09, 
    2.886419496814687e-09, 2.6618326069940426e-09, 2.4543117265218598e-09, 
    2.2625927659788086e-09, 2.0855026993786781e-09, 1.921953201326144e-09, 
    1.7709347139558063e-09, 1.6315109157072795e-09, 1.5028135657314611e-09, 
    1.3840376993591751e-09, 1.2744371516030522e-09, 1.1733203871112639e-09, 
    1.0800466163524301e-09, 9.9402217909099596e-10, 9.1469717741400366e-10, 
    8.4156234170035735e-10, 7.741461139842092e-10, 7.1201193416082635e-10, 
    6.5475571541859729e-10, 6.0200349615893964e-10, 5.5340925648998611e-10, 
    5.0865288815286438e-10, 4.6743830746482554e-10, 4.2949170154324518e-10, 
    3.9455989871240606e-10, 3.6240885459244016e-10, 3.3282224593002208e-10, 
    3.0560016475515347e-10, 2.8055790593992433e-10, 2.5752484169553901e-10, 
    2.3634337697486665e-10, 2.1686798015131896e-10, 1.9896428372239885e-10, 
    1.8250825013962272e-10, 1.6738539819700079e-10, 1.5349008571934665e-10, 
    1.4072484458075282e-10, 1.2899976435368306e-10, 1.182319211417281e-10, 
    1.0834484838494677e-10, 9.9268046647203139e-11, 9.093652960075533e-11, 
    8.3290403615600488e-11, 7.627447854058136e-11, 6.9837907430739869e-11, 
    6.3933853131771061e-11, 5.8519179778235192e-11, 5.3554167398261945e-11, 
    4.9002247944311342e-11, 4.4829761187859082e-11, 4.1005729026124825e-11, 
    3.7501646851707099e-11, 3.4291290731738963e-11, 3.1350539232354169e-11, 
    2.8657208807322638e-11, 2.6190901747045964e-11, 2.3932865756117152e-11, 
    2.1865864294647422e-11, 1.9974056880930497e-11, 1.8242888611027943e-11, 
    1.6658988204811843e-11, 1.5210073938193132e-11, 1.3884866867905667e-11, 
    1.2673010798593804e-11, 1.1564998482243995e-11, 1.0552103577454588e-11, 
    9.6263179308208358e-12, 8.7802937750174517e-12, 8.0072904681643012e-12, 
    7.3011254269046571e-12, 6.6561289314788494e-12, 6.0671025050581166e-12, 
    5.5292805918605613e-12, 5.0382952792099722e-12, 4.5901438278422316e-12, 
    4.1811587925122775e-12, 3.8079805314061108e-12, 3.4675319181114529e-12, 
    3.1569950840279982e-12, 2.8737900321880045e-12, 2.6155549755797617e-12, 
    2.3801282642927073e-12, 2.1655317761964164e-12, 1.9699556554847157e-12, 
    1.7917442923200752e-12, 1.6293834450495486e-12, 1.4814884140841265e-12, 
    1.34679318357974e-12, 1.2241404535751864e-12, 1.1124724912656493e-12, 
    1.0108227356589459e-12, 9.1830809500678064e-13, 8.3412188115682168e-13, 
    7.5752732936297028e-13, 6.8785165614585914e-13, 6.2448061154053494e-13, 
    5.668534855243254e-13, 5.1445853160845614e-13, 4.6682877352064133e-13, 
    4.2353816362173964e-13, 3.8419806420478305e-13, 3.4845402513467473e-13, 
    3.1598283341707533e-13, 2.8648981224825549e-13, 2.5970634890749335e-13, 
    2.3538763252089174e-13, 2.1331058426172731e-13, 1.9327196396734423e-13, 
    1.7508663845548804e-13, 1.5858599802271317e-13, 1.4361650871166007e-13, 
    1.3003838895038489e-13, 1.1772440010195465e-13, 1.0655874132287174e-13, 
    9.6436039920071613e-14, 8.7260429123897223e-14, 7.8944705863404747e-14, 
    7.1409561745261187e-14, 6.4582881002655047e-14, 5.8399099699871829e-14, 
    5.2798620955236834e-14, 4.7727281383245061e-14, 4.3135864359040234e-14, 
    3.8979656077794806e-14, 3.5218040720594113e-14, 3.1814131349620181e-14, 
    2.8734433440937581e-14, 2.5948538225119317e-14, 2.342884324618213e-14, 
    2.1150297769605723e-14, 1.9090170872182027e-14, 1.7227840231580557e-14, 
    1.5544599803192202e-14, 1.4023484727275426e-14, 1.2649111951858372e-14, 
    1.1407535187292198e-14, 1.0286112927810575e-14, 9.2733883848143772e-15, 
    8.3589802767145229e-15, 7.533483511785337e-15, 6.7883788843180718e-15, 
    6.1159509810536627e-15, 5.5092135650271514e-15, 4.9618417681004993e-15, 
    4.4681104821131192e-15, 4.0228383921901122e-15, 3.6213371447477179e-15, 
    3.2593651875066395e-15, 2.933085859726201e-15, 2.6390293482329196e-15, 
    2.3740581589333122e-15, 2.1353357846519834e-15, 1.920298278571578e-15, 
    1.7266284685039609e-15, 1.5522325709030914e-15, 1.3952189851359829e-15, 
    1.2538790682352576e-15, 1.1266697083282015e-15, 1.0121975313249361e-15, 
    9.0920459038580389e-16, 8.165554013036905e-16, 7.3322519934392101e-16, 
    6.582893043877351e-16, 5.9091349152220901e-16, 5.3034527359628216e-16, 
    4.7590601080134818e-16, 4.2698377010768375e-16, 3.8302686446320634e-16, 
    3.4353800809924051e-16, 3.0806903014599323e-16, 2.7621609408916251e-16, 
    2.4761537544541361e-16, 2.2193915444150092e-16, 1.9889228448813054e-16, 
    1.782090008815351e-16, 1.5965003747521782e-16, 1.430000220714523e-16, 
    1.2806512401386807e-16, 1.1467092994362231e-16, 1.0266052593477267e-16, 
    9.1892766270048994e-17, 8.2240710975160813e-17, 7.3590215914958622e-17, 
    6.5838660783990289e-17, 5.8893801711251729e-17, 5.2672736457265944e-17, 
    4.7100971322749198e-17, 4.211157992279737e-17, 3.7644444918448602e-17, 
    3.3645574647586027e-17, 3.0066487367484605e-17, 2.6863656519208622e-17, 
    2.3998011056292495e-17, 2.1434485452672177e-17, 1.9141614523277532e-17, 
    1.7091168660042484e-17, 1.5257825510903418e-17, 1.3618874513811244e-17, 
    1.215395104562311e-17, 1.0844797260410455e-17, 9.6750469763116594e-18, 
    8.6300322274229807e-18, 7.6966093298933196e-18, 6.8630025217105521e-18, 
    6.1186634257547433e-18, 5.454144757442718e-18, 4.8609868534613061e-18, 
    4.331615738237284e-18, 3.8592515713640905e-18, 3.4378264334827609e-18, 
    3.0619105112821089e-18, 2.7266458353928574e-18, 2.4276868089757198e-18, 
    2.1611468406110333e-18, 1.9235504634792436e-18, 1.7117903844956646e-18, 
    1.5230889626728913e-18, 1.3549636661205005e-18, 1.2051961022815616e-18, 
    1.0718042567316825e-18, 9.5301761256147209e-19, 8.4725485541993316e-19, 
    7.5310389907134365e-19, 6.6930399312966087e-19, 5.9472969877571455e-19, 
    5.2837653999294162e-19, 4.6934815741564725e-19, 4.1684480948296305e-19, 
    3.7015308142520877e-19, 3.2863667685181725e-19, 2.9172817951870327e-19, 
    2.5892168437018702e-19, 2.2976620730444645e-19, 2.0385979241810899e-19, 
    1.8084424384887871e-19, 1.604004168496161e-19, 1.4224400947773253e-19, 
    1.2612180234672867e-19, 1.1180829933122799e-19, 9.9102727005058981e-20, 
    8.7826354979870182e-20, 7.7820103249829557e-20, 6.8942406181770551e-20, 
    6.1067305960400539e-20, 5.4082751141937168e-20, 4.7889078519850685e-20, 
    4.2397658793088044e-20, 3.752968857720703e-20, 3.3215113136301841e-20, 
    2.9391665860255336e-20, 2.6004011987208101e-20, 2.3002985392816635e-20, 
    2.034490845159981e-20, 1.7990986035706747e-20, 1.5906765665501446e-20, 
    1.406165667589917e-20, 1.2428502022736129e-20, 1.0983197033810959e-20, 
    9.704350017928784e-21, 8.5729801897345412e-21, 7.5722488550566043e-21, 
    6.6872202368621793e-21, 5.9046487111592617e-21, 5.2127895700849121e-21, 
    4.6012307403235319e-21, 4.0607431627971733e-21, 3.5831477877270584e-21, 
    3.1611973608144914e-21, 2.7884713742215598e-21, 2.4592827327484108e-21, 
    2.1685948433581091e-21, 1.9119479769919164e-21, 1.6853938772540738e-21, 
    1.4854377026328108e-21, 1.3089864889089369e-21, 1.1533034075731364e-21, 
    1.0159671755837359e-21, 8.9483604268277504e-22, 7.8801584567080447e-22, 
    6.938316753503339e-22, 6.1080275201900651e-22, 5.376201500904909e-22, 
    4.7312705223107799e-22, 4.1630124885307884e-22, 3.6623963037166313e-22, 
    3.2214444773179461e-22, 2.8331114172216729e-22, 2.4911756384862458e-22, 
    2.1901443134121554e-22, 1.9251687648300013e-22, 1.6919696611485434e-22, 
    1.4867708110067559e-22, 1.3062405792264917e-22, 1.1474400558502953e-22, 
    1.0077772078901078e-22, 8.8496633035049306e-23, 7.7699219032639877e-23, 
    6.8207832658046016e-23, 5.9865902793169798e-23, 5.2535456788531719e-23, 
    4.609493209595919e-23, 4.0437242879304441e-23, 3.5468072194455872e-23, 
    3.1104363686344561e-23, 2.7272989728213318e-23, 2.3909575569311762e-23, 
    2.0957461399124663e-23, 1.8366786312636027e-23, 1.6093680001772496e-23, 
    1.409954962954029e-23, 1.2350450788965808e-23, 1.0816532729734349e-23, 
    9.4715491699341983e-24, 8.2924270151170881e-24, 7.2588861966086247e-24, 
    6.3531046287195392e-24, 5.5594229817546512e-24, 4.8640845847900348e-24, 
    4.2550063182058294e-24, 3.72157683900541e-24, 3.2544789092250491e-24, 
    2.8455329755947017e-24, 2.4875594827158213e-24, 2.1742576973814012e-24, 
    1.9000990827293165e-24, 1.6602334916250604e-24, 1.4504066525134832e-24, 
    1.266887601053742e-24, 1.1064048698990797e-24, 9.6609038943599696e-25, 
    8.4343017630375889e-25, 7.3622099598390844e-25, 6.4253228236557204e-25, 
    5.6067268244958298e-25, 4.8916066957578107e-25, 4.2669873491072541e-25, 
    3.7215072545429569e-25, 3.2452194842664156e-25, 2.8294170739278329e-25, 
    2.4664797558517706e-25, 2.1497394722814122e-25, 1.8733623881157003e-25, 
    1.6322453969828562e-25, 1.4219253561735094e-25, 1.2384994987959671e-25, 
    1.0785556589270032e-25, 9.3911111051926442e-26, 8.1755896605090242e-26, 
    7.1162120870473363e-26, 6.1930754431627927e-26, 5.3887935825626255e-26, 
    4.6881814942517035e-26, 4.0779789005698361e-26, 3.5466082730823523e-26, 
    3.0839630175337704e-26, 2.6812220989107069e-26, 2.3306878344847174e-26, 
    2.0256439840719298e-26, 1.7602316193326906e-26, 1.5293405636082656e-26, 
    1.3285144657278857e-26, 1.1538678099756384e-26, 1.0020133739905551e-26, 
    8.6999883031889245e-27, 7.5525134874962762e-27, 6.5552919818002366e-27, 
    5.6887947098142026e-27, 4.9360116178311974e-27, 4.2821292812650281e-27, 
    3.7142494419684523e-27, 3.2211433225795691e-27, 2.7930372075729003e-27, 
    2.4214253444923806e-27, 2.0989067127821187e-27, 1.819042640283233e-27, 
    1.5762326263729146e-27, 1.3656060624968485e-27, 1.1829278313020332e-27, 
    1.0245160198116192e-27, 8.8717020457692111e-28, 7.6810896141862612e-28, 
    6.6491542267887484e-28, 5.7548985387125393e-28, 4.9800835188692089e-28, 
    4.3088688082035273e-28, 3.7274996105288747e-28, 3.2240341426586817e-28, 
    2.7881064311221272e-28, 2.4107199072908495e-28, 2.0840678332645423e-28, 
    1.8013770979012081e-28, 1.5567723651567227e-28, 1.345157943487662e-28, 
    1.1621150825474411e-28, 1.0038126979498015e-28, 8.66929781906037e-29, 
    7.4858798179509761e-29, 6.4629302435008968e-29, 5.578838337596356e-29, 
    4.8148834076191769e-29, 4.1548510952368384e-29, 3.584700221679461e-29, 
    3.0922735936164379e-29, 2.6670470124738812e-29, 2.2999114781887134e-29, 
    1.9829842300963213e-29, 1.7094448352276105e-29, 1.4733930285239504e-29, 
    1.2697254397590279e-29, 1.094028716500186e-29, 9.4248687840475911e-30, 
    8.1180102178390718e-30, 6.9911974012675994e-30, 6.0197884091885306e-30, 
    5.1824912575796522e-30, 4.4609116308334646e-30, 3.8391612394522094e-30, 
    3.3035187389607314e-30, 2.8421362068030507e-30, 2.4447851001919149e-30, 
    2.102636422524869e-30, 1.8080705248880467e-30, 1.5545125761299966e-30, 
    1.336290262003699e-30, 1.1485107313934749e-30, 9.8695420475972518e-31, 
    8.4798200456128797e-31, 7.2845706643579926e-31, 6.2567524932375666e-31, 
    5.3730598771990221e-31, 4.613410243542543e-31, 3.9605013078334443e-31, 
    3.3994287003262472e-31, 2.9173558254712697e-31, 2.5032288686573864e-31, 
    2.147530818787132e-31, 1.8420692021001745e-31, 1.5797929387907069e-31, 
    1.3546343541123003e-31, 1.1613729126020863e-31, 9.9551770886383096e-32, 
    8.5320615064618276e-32, 7.3111661808343771e-32, 6.2639318417137216e-32, 
    5.3658074210755892e-32, 4.5956911048160374e-32, 3.9354488217573283e-32, 
    3.369499513230975e-32, 2.8844579831815879e-32, 2.4688273875359926e-32, 
    2.1127345093514623e-32, 1.8077019060662899e-32, 1.5464518270080929e-32, 
    1.3227375004691413e-32, 1.1311979951200042e-32, 9.6723338326718238e-33, 
    8.2689738469078173e-33, 7.068050592390541e-33, 6.0405345240595044e-33, 
    5.1615338804760144e-33, 4.4097085248612866e-33, 3.7667662994257447e-33, 
    3.217030352315182e-33, 2.7470675000093444e-33, 2.3453690702266915e-33, 
    2.0020768616273547e-33, 1.7087478830918229e-33, 1.4581524196975794e-33, 
    1.2441007342786628e-33, 1.0612943695022677e-33, 9.0519858030978818e-34, 
    7.7193291291399946e-34, 6.5817736517849693e-34, 5.6109192349035138e-34, 
    4.7824758125047124e-34, 4.0756721081714212e-34, 3.4727489015258047e-34, 
    2.9585248272247141e-34, 2.5200243884895977e-34, 2.1461593256756507e-34, 
    1.827455734053774e-34, 1.5558204023864122e-34, 1.3243407696475169e-34, 
    1.1271136925659774e-34, 9.5909889982345665e-35, 8.1599359542543573e-35, 
    6.9412517752461005e-35, 5.9035947145188759e-35, 5.0202224692382798e-35, 
    4.2683210796962194e-35, 3.6284311747037723e-35, 3.0839575270831862e-35, 
    2.6207498946757431e-35, 2.2267448472745265e-35, 1.8916597589656929e-35, 
    1.6067314133519511e-35, 1.3644927559748025e-35, 1.1585822596579566e-35, 
    9.8358116655796105e-36, 8.3487455439330367e-36, 7.0853275992447576e-36, 
    6.012101942538044e-36, 5.1005901391267664e-36, 4.3265547930225578e-36, 
    3.6693714669334519e-36, 3.1114930925279995e-36, 2.6379933295183461e-36, 
    2.2361773030396649e-36, 1.8952498345861056e-36, 1.606032723408118e-36, 
    1.3607238679227602e-36, 1.1526920704470245e-36, 9.7630226924384141e-37, 
    8.2676671156559318e-37, 7.0001823903140376e-37, 5.9260241848778244e-37, 
    5.0158573136342194e-37, 4.2447744431792417e-37, 3.5916313387297256e-37, 
    3.0384813640639672e-37, 2.5700944983030287e-37, 2.1735483083576545e-37, 
    1.8378801721465476e-37, 1.5537916312498427e-37, 1.3133971023151673e-37, 
    1.1100103283443821e-37, 9.3796293305251529e-38, 7.9245027867846092e-38, 
    6.6940054118674314e-38, 5.6536352487920816e-38, 4.7741625653840038e-38, 
    4.0308284058502885e-38, 3.4026643265284348e-38, 2.8719150911099332e-38, 
    2.4235488263078357e-38, 2.0448414592453252e-38, 1.7250242327389972e-38, 
    1.4549847752544262e-38, 1.2270136322292306e-38, 1.03458938187073e-38, 
    8.7219649313764827e-39, 7.3517096342961419e-39, 6.1956952156127988e-39, 
    5.2205881750870863e-39, 4.3982156090528036e-39, 3.7047702956577953e-39, 
    3.1201375956212744e-39, 2.6273255988352041e-39, 2.2119827628119086e-39, 
    1.8619896800378051e-39, 1.56711364142023e-39, 1.3187163863913569e-39, 
    1.1095068929501609e-39, 9.3333230219366264e-40, 7.8500112504740603e-40, 
    6.6013377230885801e-40, 5.5503620686369662e-40, 4.6659315951253123e-40, 
    3.9217789466167478e-40, 3.2957597397969574e-40, 2.7692085756811836e-40, 
    2.3263951391259133e-40, 1.9540649093605209e-40, 1.6410513856212732e-40, 
    1.3779487485091846e-40, 1.1568355853407283e-40, 9.7104175359211495e-41, 
    8.1495168047229974e-41, 6.8383843257660938e-41, 5.7372376620013702e-41, 
    4.8126011059029996e-41, 4.0363106385179322e-41, 3.3846751189339936e-41, 
    2.8377692956854361e-41, 2.3788380258825399e-41, 1.993794295316232e-41, 
    1.6707963437459059e-41, 1.3998914904709358e-41, 1.1727161908763685e-41, 
    9.8224348974398615e-42, 8.2257041814419212e-42, 6.8873904694586637e-42, 
    5.7658589464005387e-42, 4.8261521839164921e-42, 4.0389241879682923e-42, 
    3.3795438085684491e-42, 2.8273407319091083e-42, 2.3649714888992337e-42, 
    1.9778864681661533e-42, 1.6538819186530281e-42, 1.3827234538848702e-42, 
    1.1558297001694496e-42, 9.6600652642010762e-43, 8.0722380628138809e-43, 
    6.7442793801589137e-43, 5.6338442148500467e-43, 4.7054569603609779e-43, 
    3.9294020477951097e-43, 3.2807929203857755e-43, 2.7387908061252121e-43, 
    2.2859492987340594e-43, 1.9076645809144246e-43, 1.59171434102382e-43, 
    1.3278711407165291e-43, 1.1075782674129221e-43, 9.2367801969918172e-44, 
    7.7018398323558242e-44, 6.4209020775234603e-44, 5.3521133290621489e-44, 
    4.4604866641557721e-44, 3.716780208312157e-44, 3.0965578981639708e-44, 
    2.5794031134717687e-44, 2.1482604100275487e-44, 1.7888845797383102e-44, 
    1.4893796175259693e-44, 1.2398129892480435e-44, 1.0318929567906844e-44, 
    8.5869869824424568e-45, 7.1445462355759896e-45, 5.9434168046884668e-45, 
    4.9433961485850057e-45, 4.110951301158763e-45, 3.4181171202551926e-45, 
    2.8415757458124182e-45, 2.3618875944547456e-45, 1.9628490548503818e-45, 
    1.6309561003310484e-45, 1.3549564293140803e-45, 1.1254755863549482e-45, 
    9.3470489648230475e-46, 7.7614103772274419e-46, 6.4436874423945573e-46, 
    5.3487952797872035e-46, 4.4392047431810284e-46, 3.6836814398404926e-46, 
    3.0562343049645416e-46, 2.5352390562556022e-46, 2.1027075661173697e-46, 
    1.7436789646735694e-46, 1.4457122784933084e-46, 1.1984637457416485e-46, 
    9.933347357209502e-47, 8.2317852924236991e-47, 6.8205616114347852e-47, 
    5.650331504593058e-47, 4.6801029990232197e-47, 3.8758287845123956e-47, 
    3.209234458242661e-47, 2.6568436622795094e-47, 2.1991671678363119e-47, 
    1.820028449763627e-47, 1.5060028734349154e-47, 1.245951434657354e-47, 
    1.030633177100732e-47, 8.5238306601923996e-48, 7.0484430944279029e-48, 
    5.8274596177700727e-48, 4.817181810371864e-48, 3.981387908009545e-48, 
    3.2900586401738268e-48, 2.7183193361729471e-48, 2.2455617410815779e-48, 
    1.8547151376028148e-48, 1.5316414924947592e-48, 1.2646336093454155e-48, 
    1.0439988167361431e-48, 8.6171367192429863e-49, 7.1113761485982491e-49, 
    5.8677554878297795e-49, 4.840810211038488e-49, 3.9929308945860239e-49, 
    3.2930113084118022e-49, 2.7153282655880508e-49, 2.2386136578827213e-49, 
    1.8452858346751865e-49, 1.5208130724259163e-49, 1.2531865242448894e-49, 
    1.0324838938844401e-49, 8.5050827875273237e-50, 7.0048928297267567e-50, 
    5.7683570613888186e-50, 4.7493094277311843e-50, 3.9096374516910907e-50, 
    3.2178826122512699e-50, 2.6480830293545305e-50, 2.1788166695888897e-50, 
    1.7924104643951085e-50, 1.4742866821533141e-50, 1.2124228263759655e-50, 
    9.9690541810650115e-51, 8.1956140570864558e-51, 6.7365374924881947e-51, 
    5.5363004895893718e-51, 4.5491501025442113e-51, 3.7373912984825217e-51, 
    3.0699730536915209e-51, 2.5213216159541482e-51, 2.0703778895602632e-51, 
    1.6998033666085699e-51, 1.3953252049869981e-51, 1.1451961619608793e-51, 
    9.3974931661309715e-52, 7.7103100692373948e-52, 6.3249829430524061e-52, 
    5.1876965449628657e-52, 4.2541956544141797e-52, 3.4880929181925519e-52, 
    2.8594751155975044e-52, 2.343755411033157e-52, 1.9207283392842378e-52, 
    1.5737918461384048e-52, 1.2893069620612621e-52, 1.0560708491868979e-52, 
    8.6488322203797886e-53, 7.0818965726536997e-53, 5.7978820717521797e-53, 
    4.7458812322693942e-53, 3.8841146772291656e-53, 3.1783001783402534e-53, 
    2.6003120643171338e-53, 2.1270794890026535e-53, 1.7396811544837406e-53, 
    1.4226015849097187e-53, 1.1631202254937646e-53, 9.5080973023535239e-54, 
    7.7712399271509193e-54, 6.3505992482748282e-54, 5.1887982881667799e-54, 
    4.2388354590711796e-54, 3.462214887605054e-54, 2.8274124798076278e-54, 
    2.3086176512263243e-54, 1.8847013574867472e-54, 1.5383698689929307e-54, 
    1.255470975659207e-54, 1.0244252612545966e-54, 8.3575998047297339e-55, 
    6.8172709331004053e-55, 5.5599031556810009e-55, 4.5336875877465362e-55, 
    3.6962696237258765e-55, 3.0130295202311345e-55, 2.4556746125382989e-55, 
    2.0010868788338894e-55, 1.6303796968649619e-55, 1.3281259511834971e-55, 
    1.0817264706035098e-55, 8.8089337163345565e-56, 7.1722747380877371e-56, 
    5.8387271721592731e-56, 4.7523359910706088e-56, 3.8674417694344488e-56, 
    3.1467925933393839e-56, 2.5600010614607921e-56, 2.0822835187330454e-56, 
    1.6934300739629393e-56, 1.376963299211346e-56, 1.1194511632000473e-56, 
    9.0994601863543311e-57, 7.3952659455396219e-57, 6.0092414491443944e-57, 
    4.8821734204900067e-57, 3.9658331626758968e-57, 3.2209454402184407e-57, 
    2.6155316929980993e-57, 2.1235588231086627e-57, 1.723837382768294e-57, 
    1.3991232825029608e-57, 1.1353855509010785e-57, 9.2120955223496337e-58, 
    7.4731068605206176e-58, 6.0613818256321132e-58, 4.9155235678920657e-58, 
    3.98561746402706e-58, 3.2310905852861749e-58, 2.6189689211709904e-58, 
    2.122458688438552e-58, 1.7197916548024222e-58, 1.3932855044282811e-58, 
    1.1285793265972796e-58, 9.1401169477552055e-59, 7.4011482717060573e-59, 
    5.9920323201319228e-59, 4.8503924573306861e-59, 3.9256113690520934e-59, 
    3.1766210967746697e-59, 2.5701070868192321e-59, 2.0790489404863747e-59, 
    1.6815349424505487e-59, 1.3597991657369935e-59, 1.0994394964426995e-59, 
    8.8878269269477611e-60, 7.183689185891788e-60, 5.8053334286396805e-60, 
    4.690665821768942e-60, 3.7893917806722359e-60, 3.0607807004690761e-60, 
    2.4718528298816248e-60, 1.9959088135481357e-60, 1.6113373431056489e-60, 
    1.3006484821395668e-60, 1.0496900850413422e-60, 8.4701273846389474e-61, 
    6.8335516121133119e-61, 5.5122728463921999e-61, 4.4457252931342606e-61, 
    3.5849428054791914e-61, 2.8903439663136276e-61, 2.3299388195941388e-61, 
    1.8778772285567951e-61, 1.5132739784311159e-61, 1.2192580256830955e-61, 
    9.8220326165688278e-62, 7.9110624199084582e-62, 6.3708288875265885e-62, 
    5.1296148777345196e-62, 4.1295361297895411e-62, 3.3238810249654024e-62, 
    2.6749604211268122e-62, 2.1523700541166567e-62, 1.7315865820392664e-62, 
    1.3928334007275439e-62, 1.120164548988523e-62, 9.0072489308067309e-63, 
    7.2415277123489504e-63, 5.8209774765320109e-63, 4.6783136056349965e-63, 
    3.7593298505129824e-63, 3.020363585835492e-63, 2.4262508938455034e-63, 
    1.9486770990142267e-63, 1.5648465058396743e-63, 1.2564097496978676e-63, 
    1.0085990190635037e-63, 8.0953098334411917e-64, 6.496449985486622e-64, 
    5.2125041472495477e-64, 4.1816185916604099e-64, 3.3540544806568284e-64, 
    2.6898217288590781e-64, 2.1567736684782349e-64, 1.7290730351363685e-64, 
    1.385957119054446e-64, 1.1107439064263619e-64, 8.9003231543179712e-65, 
    7.1305873040438386e-65, 5.7117937646547339e-65, 4.5745399496768176e-65, 
    3.6631105160920972e-65, 2.9327855553456341e-65, 2.3476766794367485e-65, 
    1.8789877704003879e-65, 1.5036172907137696e-65, 1.2030352677994206e-65, 
    9.6238112648208998e-66, 7.6973906104216836e-66, 6.1555610702667926e-66, 
    4.9217489034898139e-66, 3.9345851841574583e-66, 3.1448949384558522e-66, 
    2.513280843653642e-66, 2.0081844078046899e-66, 1.6043305395732543e-66, 
    1.2814799063910286e-66, 1.0234283453003566e-66, 8.1720454205551564e-67, 
    6.5242680026356031e-67, 5.2078744235183005e-67, 4.1563958724616058e-67, 
    3.3166603303957468e-67, 2.6461397576773454e-67, 2.1108251007256272e-67, 
    1.6835243878348546e-67, 1.3424999072749706e-67, 1.0703770946967516e-67, 
    8.5327110634928752e-68, 6.8008776638560207e-68, 5.4196417029475043e-68, 
    4.3182111986039864e-68, 3.4400509350938643e-68, 2.7400188897544266e-68, 
    2.1820762929345069e-68, 1.7374567205143881e-68, 1.3832024508775375e-68, 
    1.1009946142455318e-68, 8.7621832063394324e-69, 6.9721569457990968e-69, 
    5.5468914889283548e-69, 4.412247601479976e-69, 3.5091163774323105e-69, 
    2.790380045766112e-69, 2.2184857009909025e-69, 1.7635086749186075e-69, 
    1.4016069976043406e-69, 1.1137881783149951e-69, 8.8492535990368598e-70, 
    7.0297255275514542e-70, 5.5833877078783098e-70, 4.4338897894381419e-70, 
    3.5204622516897745e-70, 2.7947449507054525e-70, 2.2182595435321641e-70, 
    1.7603954091800015e-70, 1.3968050169175229e-70, 1.1081257205512336e-70, 
    8.7896174695726113e-71, 6.9707355033042544e-71, 5.5273240160458581e-71, 
    4.3820661982748882e-71, 3.4735266415697544e-71, 2.7528973938427985e-71, 
    2.181409023558515e-71, 1.7282711333883886e-71, 1.3690343255230597e-71, 
    1.084287593456348e-71, 8.5862262890685821e-72, 6.7981049003744446e-72, 
    5.3814719853268794e-72, 4.2593369315682399e-72, 3.3706262474495137e-72, 
    2.6669009800836776e-72, 2.1097494085988574e-72, 1.6687164487863288e-72, 
    1.3196595657152311e-72, 1.0434435615542477e-72, 8.249045656920339e-73, 
    6.5202784275501509e-73, 5.152953998347018e-73, 4.0716841349221121e-73, 
    3.2167668487574228e-73, 2.5409304583192104e-73, 2.0067518139107415e-73, 
    1.5846094422957825e-73, 1.2510610550383937e-73, 9.8755765689448062e-74, 
    7.7942459591932487e-74, 6.1505427663251188e-74, 4.8526667629750936e-74, 
    3.828028702920567e-74, 3.0192396921596216e-74, 2.380935822468511e-74, 
    1.8772645387658294e-74, 1.4798951739028052e-74, 1.1664446124662203e-74, 
    9.1923167183855245e-75, 7.2429173178621402e-75, 5.7059737030755853e-75, 
    4.4944204126540684e-75, 3.5395276808275502e-75, 2.7870491141135918e-75, 
    2.194176812392547e-75, 1.7271351012747015e-75, 1.359279259308208e-75, 
    1.0695935124105838e-75, 8.4150464993194647e-76, 6.6194509802717756e-76, 
    5.2061312274318187e-76, 4.0938878535663336e-76, 3.2187293675808471e-76, 
    2.5302339207560184e-76, 1.9886784840315547e-76, 1.5627739618431315e-76, 
    1.2278786510635856e-76, 9.64589256406926e-77, 7.57629859596654e-77, 
    5.9497598291341066e-77, 4.671641177638466e-77, 3.6674754107382935e-77, 
    2.8786749845691617e-77, 2.2591535351542878e-77, 1.7726645133418533e-77, 
    1.3907050910048169e-77, 1.0908655543189045e-77, 8.5552972339613695e-78, 
    6.7085192006794267e-78, 5.2595177094098477e-78, 4.1228056888406935e-78, 
    3.2312272425094416e-78, 2.5320357138348894e-78, 1.9838089375910788e-78, 
    1.5540233795984078e-78, 1.2171467512995806e-78, 9.5313853976452143e-79, 
    7.4627141498094359e-79, 5.8420500512357463e-79, 4.5725812404093841e-79, 
    3.5783702730234603e-79, 2.7998632138854603e-79, 2.1903627347509823e-79, 
    1.7132587549459952e-79, 1.3398542794577066e-79, 1.0476588014125854e-79, 
    8.1904894307119776e-80, 6.4021748766945323e-80, 5.0034884501431698e-80, 
    3.9097227432721705e-80, 3.0545462819686697e-80, 2.3860258767221242e-80, 
    1.8635080750876197e-80, 1.4551745777949347e-80, 1.1361262886269998e-80, 
    8.8688193614428146e-81, 6.9220176112274681e-81, 5.4016604481218363e-81, 
    4.2145339018519503e-81, 3.2877554993596568e-81, 2.5643491965696945e-81, 
    1.9997813137273067e-81, 1.5592492284002956e-81, 1.2155596065403152e-81, 
    9.4746826456318351e-82, 7.3838144512319434e-82, 5.7533999793876188e-82, 
    4.4822497370390194e-82, 3.4913647562284043e-82, 2.7190806356124769e-82, 
    2.1172719337010813e-82, 1.6483858751060378e-82, 1.2831245620498961e-82, 
    9.9863421746331763e-83, 7.7709078188559304e-83, 6.0459529333341607e-83, 
    4.703113469643361e-83, 3.6579169589975743e-83, 2.8445260632290997e-83, 
    2.2116361649753087e-83, 1.7192741711377552e-83, 1.3363009734846383e-83, 
    1.0384632238346552e-83, 8.0687386273177457e-84, 6.2682724409849513e-84, 
    4.8687533187960769e-84, 3.7810756635535203e-84, 2.935895920613143e-84, 
    2.2792587622472243e-84, 1.7691892866132345e-84, 1.373038322269799e-84, 
    1.065414754881653e-84, 8.2657534193778322e-85, 6.4117100441024746e-85, 
    4.9727084003572623e-85, 3.8560246546378828e-85, 2.9896083740904729e-85, 
    2.3174826467881742e-85, 1.7961655835539469e-85, 1.3918868779829789e-85, 
    1.0784231466086291e-85, 8.3541477357746206e-86, 6.4705737526116761e-86, 
    5.0108467722047526e-86, 3.8797803900124867e-86, 3.0035222592803188e-86, 
    2.3247821177292368e-86, 1.7991250400612921e-86, 1.3920926163982199e-86, 
    1.0769675111360847e-86, 8.3303790753500318e-87, 6.4425028164707708e-87, 
    4.9816379352311433e-87, 3.8513890640835204e-87, 2.9770787043282211e-87, 
    2.3008638969369081e-87, 1.7779487301331795e-87, 1.373647269354751e-87, 
    1.0611063445670146e-87, 8.1954024568603298e-88, 6.3286248201091274e-88, 
    4.8862547421227575e-88, 3.7719901494884079e-88, 2.9113383761251171e-88, 
    2.2466866802210648e-88, 1.7334847531850589e-88, 1.3372888760818595e-88, 
    1.0314736266107704e-88, 7.9546067504751131e-89, 6.1334805292648873e-89, 
    4.728495256293838e-89, 3.6447405167057515e-89, 2.8089108897778639e-89, 
    2.1643973782820827e-89, 1.6674918763782246e-89, 1.2844527847414472e-89, 
    9.8923677443819727e-90, 7.6174576949524638e-90, 5.8647234715173605e-90, 
    4.5145318171270074e-90, 3.4746061745188028e-90, 2.6737829293014802e-90, 
    2.0571899575191685e-90, 1.5825241095522678e-90, 1.2171776381752442e-90, 
    9.3602033738763613e-91, 7.1968805608458362e-91, 5.5326219531577463e-91, 
    4.2525104189793736e-91, 3.2680407802114226e-91, 2.5110608577387625e-91, 
    1.9290998162971534e-91, 1.4817667704256404e-91, 1.1379749260419459e-91, 
    8.7380238341974867e-92, 6.7084385690435428e-92, 5.1494086665273824e-92, 
    3.9520366390225137e-92, 3.0325799207426173e-92, 2.3266509711945589e-92, 
    1.7847521404616581e-92, 1.3688386995521834e-92, 1.0496737309853687e-92, 
    8.0479278208524771e-93, 6.169379795917748e-93, 4.7285352534455159e-93, 
    3.6235932823490343e-93, 2.7763866705994325e-93, 2.1269052621687385e-93, 
    1.6290860732989861e-93, 1.2475777091754459e-93, 9.5525401601409433e-94, 
    7.3130379664503506e-94, 5.5976336835095184e-94, 4.2838949315704593e-94, 
    3.2779387719445343e-94, 2.5077864645103251e-94, 1.9182621648881673e-94, 
    1.467077505771194e-94, 1.1218268898370324e-94, 8.5768205460603633e-95, 
    6.5562346882051747e-95, 5.0108378512786606e-95, 3.8290752182578174e-95, 
    2.92553390895595e-95, 2.234827799555867e-95, 1.706910240784803e-95, 
    1.3034818646413524e-95, 9.9523809809561671e-96, 7.5976045006951285e-96, 
    5.799012730147529e-96, 4.4254672605611827e-96, 3.3766954489688333e-96, 
    2.5760384618064807e-96, 1.9649001407073033e-96, 1.498498507416315e-96, 
    1.1426147758106757e-96, 8.711060846092533e-97, 6.6400285832274162e-97, 
    5.0605362561231528e-97, 3.8561225068928139e-97, 2.9378714919748424e-97, 
    2.2379091785148031e-97, 1.7044325137142935e-97, 1.2979108205606862e-97, 
    9.8818347313459347e-98, 7.52242748008082e-98, 5.7254038168749719e-98, 
    4.3569434886335708e-98, 3.3150144133016394e-98, 2.5218346360993947e-98, 
    1.9181187015082667e-98, 1.4586867711973423e-98, 1.109114285934271e-98, 
    8.4317601551823064e-99, 6.4089647022706625e-99, 4.8706307381986187e-99, 
    3.7009244621286895e-99, 2.8116608061731443e-99, 2.135715124369163e-99, 
    1.6220020904808274e-99, 1.2316496456731406e-99, 9.3508405846398291e-100, 
    7.0980950422985236e-100, 5.3871697136894149e-100, 
    4.0879652461880655e-100, 3.1015688246759428e-100, 
    2.3527909482917729e-100, 1.7844851936340952e-100, 1.353225731371052e-100, 
    1.0260186046380703e-100, 7.7779995676207863e-101, 
    5.8953322168954418e-101, 4.4676211986568231e-101, 
    3.3851045960915942e-101, 2.5644576543278136e-101, 
    1.9424357479526288e-101, 1.4710433877101613e-101, 
    1.1138635505781361e-101, 8.4326911249590761e-102, 
    6.3830476127025884e-102, 4.8307845089566458e-102, 
    3.6554002415200878e-102, 2.7655397025052875e-102, 
    2.0919560169479612e-102, 1.5821690737037402e-102, 
    1.1964124489351252e-102, 9.0455847220081968e-103, 
    6.8378576931075302e-103, 5.1681030048643042e-103, 
    3.9054398550604506e-103, 2.950777322482862e-103, 2.2291054338833839e-103, 
    1.6836525567542704e-103, 1.271458027286272e-103, 9.6001777040351351e-104, 
    7.2474329544398255e-104, 5.4703716271222679e-104, 
    4.1283560471836119e-104, 3.1150509227702265e-104, 
    2.3500702557774342e-104, 1.7726550456120406e-104, 
    1.3368888672316551e-104, 1.0080778506738616e-104, 
    7.6001213848420227e-105, 5.7289452905213976e-105, 
    4.3177402423432963e-105, 3.2536140745945873e-105, 
    2.4513383240756465e-105, 1.8465801473877701e-105, 
    1.3907874384655357e-105, 1.0473239790959584e-105, 
    7.8854961651230399e-106, 5.9361476261320276e-106, 
    4.4679473946038055e-106, 3.3623204308516049e-106, 2.529867863035451e-106, 
    1.9031992904561955e-106, 1.4315231848675426e-106, 
    1.0765648490458967e-106, 8.0948665801207292e-107, 
    6.0856487865948243e-107, 4.574375003496359e-107, 3.4378295086308076e-107, 
    2.5832390399014656e-107, 1.9407631884353123e-107, 
    1.4578343766322851e-107, 1.0948925936636419e-107, 
    8.2217172929719733e-108, 6.1727864242329141e-108, 
    4.6336972232857117e-108, 3.4777771082916901e-108, 
    2.6097777650080179e-108, 1.9580915761705223e-108, 
    1.4688930015427332e-108, 1.1017295918204135e-108, 
    8.2620450277377476e-109, 6.1948071479038318e-109, 4.644037460648669e-109, 
    3.4808982447605131e-109, 2.608642898617258e-109, 1.9546347973614102e-109, 
    1.4643480404320337e-109, 1.09685870162962e-109, 8.2145683915964379e-110, 
    6.1510110152113762e-110, 4.6050669658065199e-110, 
    3.4470936740986112e-110, 2.5798705271895493e-110, 
    1.9305027605652953e-110, 1.4443439715550826e-110, 
    1.0804347138610203e-110, 8.0807954945722355e-111, 
    6.0427884817154281e-111, 4.5180221910304438e-111, 
    3.3774351344146075e-111, 2.5243720576794096e-111, 
    1.8864591355206691e-111, 1.4095131430070195e-111, 
    1.0529761824635325e-111, 7.864944388735913e-112, 5.8735470860659788e-112, 
    4.3856396378564312e-112, 3.2741089150169911e-112, 
    2.4438862702549005e-112, 1.8238812173239963e-112, 
    1.3609425749679653e-112, 1.0153382337001205e-112, 
    7.5737221823393515e-113, 5.6485332639586651e-113, 4.21201298246786e-113, 
    3.1403018989688814e-113, 2.3408888483914508e-113, 
    1.7446884012289694e-113, 1.3001176231850884e-113, 
    9.6866834295777363e-114, 7.2159789657245103e-114, 
    5.3745622895870939e-114, 4.0023828857008233e-114, 
    2.9800383653719818e-114, 2.2184659529545705e-114, 
    1.6512444496396292e-114, 1.2288465765836701e-114, 
    9.1434826943346362e-115, 6.8022614568739587e-115, 
    5.0596757341261278e-115, 3.7628745400788105e-115, 
    2.7979792069200089e-115, 2.0801608439259505e-115, 
    1.5462404907642034e-115, 1.1491715261539196e-115, 
    8.5392624522076194e-116, 6.3442977490308938e-116, 
    4.7127504384212019e-116, 3.5002012714597026e-116, 2.599197521289129e-116, 
    1.9298041692507068e-116, 1.432566815304602e-116, 1.0632716227862377e-116, 
    7.8904405160533988e-117, 5.8544481927331274e-117, 
    4.3430854527843043e-117, 3.2213541419237172e-117, 
    2.3889455962558906e-117, 1.7713392154959319e-117, 1.313181953188507e-117, 
    9.7336508534975549e-118, 7.2136374709022422e-118, 
    5.3451580509415483e-118, 3.9599935668010458e-118, 
    2.9332974157428908e-118, 2.1724280869090359e-118, 
    1.6086531315247535e-118, 1.1909872127213948e-118, 
    8.8161603115955422e-119, 6.5249854718874397e-119, 
    4.8284452310794766e-119, 3.5724220421549508e-119, 
    2.6426880527088416e-119, 1.9545947706139814e-119, 
    1.4454239747170696e-119, 1.0687139186337378e-119, 
    7.9005143713015757e-120, 5.8395174354781672e-120, 
    4.3154515168495113e-120, 3.1886232927764818e-120, 
    2.3556343413402417e-120, 1.7399638684459511e-120, 1.284991553915891e-120, 
    9.4882912344489291e-121, 7.0049240376624938e-121, 
    5.1706666972528312e-121, 3.8160789219972913e-121, 
    2.8158910160568918e-121, 2.0775047560591279e-121, 
    1.5324838322277392e-121, 1.1302576789432814e-121, 
    8.3346376096637697e-122, 6.1450251797898723e-122, 
    4.5298967407295303e-122, 3.3387248389613224e-122, 
    2.4603712534091778e-122, 1.8127935629235712e-122, 
    1.3354380518590242e-122, 9.8361882860474211e-123, 
    7.2436525442486789e-123, 5.3335463977499967e-123, 
    3.9264695587554284e-123, 2.8901213772554836e-123, 
    2.1269516621522279e-123, 1.5650450672394745e-123, 1.151393481091911e-123, 
    8.4693167307292143e-124, 6.2287467460827782e-124, 
    4.5801601324035187e-124, 3.3673506375343046e-124, 
    2.4752764532631206e-124, 1.8192264850066086e-124, 
    1.3368341145330774e-124, 9.8219102124828697e-125, 
    7.2150955997012239e-125, 5.2992683243039493e-125, 
    3.8915034591874101e-125, 2.8572393436800107e-125, 
    2.0975074531099774e-125, 1.5395297793642198e-125, 
    1.1297968652995364e-125, 8.2897288831580208e-126, 6.081461742757003e-126, 
    4.4607031325451913e-126, 3.2713450432986975e-126, 
    2.3987063016935818e-126, 1.7585531096069601e-126, 
    1.2890257465088275e-126, 9.4470319706310541e-127, 
    6.9224028345729445e-127, 5.0716122504135174e-127, 
    3.7150349692377648e-127, 2.7208679199690626e-127, 
    1.9924145495870212e-127, 1.4587458685193321e-127, 1.067842652601356e-127, 
    7.8156045808883543e-128, 5.7193356405022932e-128, 
    4.1846224376135726e-128, 3.0612208666095271e-128, 2.239034270222284e-128, 
    1.6373989476145567e-128, 1.1972255132329606e-128, 8.752358731624153e-129, 
    6.3973770268323548e-129, 4.6752675956176937e-129, 
    3.4161638334503856e-129, 2.4957357376050822e-129, 
    1.8229980139903327e-129, 1.331378328181114e-129, 9.721750282357321e-130, 
    7.09765898973421e-130, 5.1809987572021495e-130, 3.7812860875510338e-130, 
    2.7592641331390977e-130, 2.0131433686615302e-130, 
    1.4685333855425845e-130, 1.0710768526798897e-130, 
    7.8106132449085467e-131, 5.694784883456347e-131, 4.1514250711904553e-131, 
    3.025831740298645e-131, 2.2050580893978823e-131, 1.6066563164261136e-131, 
    1.1704520506388214e-131, 8.5253449079917708e-132, 
    6.2086614602496741e-132, 4.5207624964687626e-132, 
    3.2911910507534578e-132, 2.3956434737770197e-132, 
    1.7434880219308124e-132, 1.2686547231714842e-132, 
    9.2298704114814742e-133, 6.7139090934099727e-133, 
    4.8829581246812021e-133, 3.5507347737044e-133, 2.581553662425753e-133, 
    1.8766002551699141e-133, 1.363923697826467e-133, 9.9114243286260582e-134, 
    7.201280940231802e-134, 5.2313181010278843e-134, 3.7996202540307333e-134, 
    2.7592874730600872e-134, 2.0034633158945741e-134, 
    1.4544323658536124e-134, 1.0556825827111768e-134, 
    7.6612718414878611e-135, 5.5589923813947958e-135, 
    4.0329141339439943e-135, 2.925294281563936e-135, 2.1215234629112229e-135, 
    1.5383452200098051e-135, 1.1152891156768555e-135, 
    8.0844189522807791e-136, 5.8591936155646636e-136, 
    4.2457515565331031e-136, 3.0760897020887564e-136, 
    2.2282868859217403e-136, 1.6138787494006427e-136, 
    1.1686874814686881e-136, 8.4616210406090188e-137, 
    6.1254280177540686e-137, 4.4335029349222878e-137, 
    3.2083759347695954e-137, 2.3214064682939151e-137, 
    1.6793639280013337e-137, 1.2146919154722651e-137, 
    8.7844616606733493e-138, 6.3517274242456568e-138, 4.591940412858012e-138, 
    3.3191610480666038e-138, 2.3987671723678023e-138, 
    1.7333072701212581e-138, 1.2522490492913e-138, 9.0455203059266631e-139, 
    6.5328710421484085e-139, 4.7173957132350838e-139, 
    3.4058712060187147e-139, 2.4585657323134423e-139, 
    1.7744473484098879e-139, 1.280477940410714e-139, 9.238655537801538e-140, 
    6.6645854216756485e-140, 4.8069011688916805e-140, 
    3.4664499770913958e-140, 2.4993804709427404e-140, 
    1.8018037937024837e-140, 1.2987044004974187e-140, 
    9.3592450282263393e-141, 6.7437119704837456e-141, 
    4.8583063731426301e-141, 3.4994393794387471e-141, 
    2.5202274692237883e-141, 1.8147161208565929e-141, 1.306487755627114e-141, 
    9.4043694221496163e-142, 6.7683328453552089e-142, 
    4.8703640500427311e-142, 3.5040382040895024e-142, 
    2.5205999905930654e-142, 1.81287023404383e-142, 1.3036385555782992e-142, 
    9.3729298097542258e-143, 6.7378482159824362e-143, 
    4.8427803570103776e-143, 3.480134358672084e-143, 2.5004889545350647e-143, 
    1.7963111264192504e-143, 1.2902262385409998e-143, 9.265692208479196e-144, 
    6.6530005548115124e-144, 4.776226787293932e-144, 3.4283094086750803e-144, 
    2.4603833044926732e-144, 1.7654410572389274e-144, 
    1.2665763182767688e-144, 9.085256540900285e-145, 6.5158445796391073e-145, 
    4.6723129991336871e-145, 3.3498150593568266e-145 ;

 frequency_resolution = 1, 0.99261774516933099, 0.97079636050239726, 
    0.93548820017660983, 0.88820365913169719, 0.83090404247139049, 
    0.76586682126361416, 0.69553615292009763, 0.622372266754739, 
    0.54871246348221436, 0.47665426958208207, 0.40796811316024911, 
    0.34404323452402669, 0.28586691435094636, 0.2340339353901679, 
    0.18878081076006786, 0.15003788311580848, 0.11749194111254087, 
    0.090652398571217541, 0.068915131623251372, 0.051619518608300566, 
    0.038095824730339192, 0.02770160163770502, 0.019847072173656798, 
    0.014010450115364264, 0.009744774573919401, 0.0066781408662551422, 
    0.0045092407602355875, 0.0029999591579678501, 0.0019664881335663019, 
    0.0012700809080201608, 0.00080823102076036778, 0.00050676161583864949, 
    0.00031306605390129697, 0.00019056025082514889, 0.00011428591828011938, 
    6.753317969967008e-05, 3.9319296985640725e-05, 2.2555806479683745e-05, 
    1.2748968416909115e-05, 7.0999583390887694e-06, 3.8958356308625014e-06, 
    2.1062480683728268e-06, 1.1219732027087135e-06, 5.8887012031205955e-07, 
    3.0452336657006711e-07, 1.5516215259126554e-07, 7.7895978909022787e-08, 
    3.8530828955133e-08, 1.8778709147316588e-08, 9.017521534215219e-09, 
    4.2665094362927225e-09, 1.9889428422427242e-09, 9.135576623570703e-10, 
    4.1344114640211354e-10, 1.8435524482647913e-10, 8.0995589150602872e-11, 
    3.5061566001196529e-11, 1.4954273537233289e-11, 6.2843939335640229e-12, 
    2.6021093958042384e-12, 1.0615776604428162e-12, 4.2671907844331635e-13, 
    1.6900378059331838e-13, 6.5950007457414576e-14, 2.5356969478790034e-14, 
    9.6060295118521347e-15, 3.5855398608161929e-15, 1.3186491620066904e-15, 
    4.7782408961678024e-16, 1.7059680319517759e-16, 6.0011959305108679e-17, 
    2.0800261419799363e-17, 7.1033604053906331e-18, 2.3901380010066185e-18, 
    7.9240311339391141e-19, 2.5884122076058104e-19, 8.3307629196209175e-20, 
    2.641801491111585e-20, 8.2542887342006454e-21, 2.5411084569313597e-21, 
    7.7078067316551929e-22, 2.3035757665043587e-22, 6.7832567481344019e-23, 
    1.9680588450170413e-23, 5.6260290928610951e-24, 1.5846375296304793e-24, 
    4.3976632540830865e-25, 1.2024805872123126e-25, 3.2396511461358676e-26, 
    8.5996839268655335e-27, 2.249214123320825e-27, 5.7961976176996076e-28, 
    1.4717011728022023e-28, 3.6817996969304753e-29, 9.075378545527232e-30, 
    2.2041107373001261e-30, 5.2743159397270448e-31, 1.2435491123068966e-31, 
    2.8888421510327814e-32, 6.6122421915388192e-33, 1.4912064117168108e-33, 
    3.3135295045426587e-34, 7.2545084589830411e-35, 1.5649094409568821e-35, 
    3.3260938523799135e-36, 6.9653646616543403e-37, 1.4372002584955368e-37, 
    2.9218289297508565e-38, 5.8527012034687326e-39, 1.1551064008190923e-39, 
    2.2462169383074462e-40, 4.3037345341003211e-41, 8.1246249464356996e-42, 
    1.5112114611276017e-42, 2.7695628499163051e-43, 5.0010509748114035e-44, 
    8.8976518222953907e-45, 1.5597450027341015e-45, 2.6939893114371518e-46, 
    4.5846079534028693e-47, 7.6872783786545756e-48, 1.2700098319022286e-48, 
    2.067310105318453e-49, 3.3156466525963878e-50, 5.2395612990899403e-51, 
    8.1580371625676894e-52, 1.2515278052088468e-52, 1.8917310663439212e-53, 
    2.817360094513939e-54, 4.1341800945745467e-55, 5.9772372462253003e-56, 
    8.5148238160788401e-57, 1.1951293395894031e-57, 1.6527920676535225e-58, 
    2.252089269347806e-59, 3.0235492871624356e-60, 3.9995632887330613e-61, 
    5.2128132209785886e-62, 6.6941559329651766e-63, 8.4700028164416734e-64, 
    1.0559305492500143e-64, 1.2970335929363968e-65, 1.5697524292675667e-66, 
    1.8718677975248016e-67, 2.199293810372404e-68, 2.5459824207693195e-69, 
    2.9039666139657635e-70, 3.2635622976979149e-71, 3.613734694177164e-72, 
    3.9426179327858826e-73, 4.2381584593050646e-74, 4.4888361951812808e-75, 
    4.6844045543159969e-76, 4.8165835848175498e-77, 4.8796410672238694e-78, 
    4.8708047836429318e-79, 4.7904646509845745e-80, 4.6421441852538504e-81, 
    4.4322442063079156e-82, 4.1695847554126759e-83, 3.8647908933476904e-84, 
    3.5295819177440887e-85, 3.1760300313711097e-86, 2.8158531656030214e-87, 
    2.4597981948505653e-88, 2.1171567922801799e-89, 1.7954389216793835e-90, 
    1.5002109078106513e-91, 1.235088482359726e-92, 1.0018619771452083e-93, 
    8.0072204784350036e-95, 6.3055031815650929e-96, 4.8923980130095541e-97, 
    3.7401402059662941e-98, 2.8172024297406402e-99, 2.0907990567393596e-100, 
    1.5288701675150353e-101, 1.1015215224165497e-102, 
    7.8195081679025091e-104, 5.4692774834770614e-105, 
    3.7691597765791946e-106, 2.5593118499102693e-107, 
    1.7122451194432216e-108, 1.1286849552883625e-109, 
    7.3306689123104159e-111, 4.6911416188130479e-112, 
    2.9578595777676105e-113, 1.8375562003669485e-114, 
    1.1247805000429278e-115, 6.7835807052818862e-117, 4.031013788468421e-118, 
    2.3601175857254664e-119, 1.3614981886510525e-120, 
    7.7386385882020221e-122, 4.3338725059226871e-123, 
    2.3913974801949678e-124, 1.3001440513607172e-125, 
    6.9645850936371457e-127, 3.6758949742489017e-128, 
    1.9115911432053671e-129, 9.7946967532132999e-131, 
    4.9448264013864242e-132, 2.4596605399142604e-133, 
    1.2054893226606119e-134, 5.821241704344082e-136, 2.7696951196676384e-137, 
    1.2984115474494407e-138, 5.9973147564389372e-140, 
    2.7293886764820397e-141, 1.2238776337607487e-142, 
    5.4072279790613825e-144, 2.353831838221619e-145, 1.0095788756516719e-146, 
    4.266474424441769e-148, 1.7764873039571162e-149, 7.2881808255309154e-151, 
    2.9460508608709526e-152, 1.1733441462336998e-153, 
    4.6044170293504101e-155, 1.7802785602960485e-156, 
    6.7821180004211994e-158, 2.5456974728070847e-159, 
    9.4148262794002735e-161, 3.4306933455879086e-162, 
    1.2317301131624612e-163, 4.3572581195031965e-165, 
    1.5187108174459813e-166, 5.2155601041134374e-168, 
    1.7647812972350999e-169, 5.883623857247137e-171, 1.9326934632452811e-172, 
    6.255256531111281e-174, 1.9947631742181154e-175, 6.2676051501405565e-177, 
    1.9403317279309654e-178, 5.9185376065443674e-180, 
    1.7787581684165074e-181, 5.2672444379295681e-183, 
    1.5367885237609006e-184, 4.4178281070912298e-186, 
    1.2513177034128535e-187, 3.4921302496194261e-189, 
    9.6023459419342241e-191, 2.6015269689410139e-192, 
    6.9445384432090263e-194, 1.8265119172032965e-195, 
    4.7333182271780889e-197, 1.2085732203195848e-198, 
    3.0404950441791857e-200, 7.5366735213561459e-202, 
    1.8406837366103459e-203, 4.4293777257780722e-205, 1.050195926376258e-206, 
    2.4533641290500819e-208, 5.6469996732503559e-210, 1.280671025213314e-211, 
    2.8616826790569151e-213, 6.3004190447103977e-215, 
    1.3667260307718786e-216, 2.921174940467678e-218, 6.1517366627393808e-220, 
    1.2764446168217088e-221, 2.6095780192898865e-223, 
    5.2565725746841254e-225, 1.0432757527580585e-226, 
    2.0401384107686173e-228, 3.9308296307644725e-230, 
    7.4623030031569328e-232, 1.3958077565403403e-233, 2.572423125504091e-235, 
    4.6711441818543642e-237, 8.3573426759520755e-239, 
    1.4732526023576454e-240, 2.5588822022313727e-242, 
    4.3791259889473833e-244, 7.3839484562568223e-246, 
    1.2267439997560149e-247, 2.0080905769189012e-249, 
    3.2387447627115265e-251, 5.1467635784049818e-253, 
    8.0585292012334813e-255, 1.2432011945059032e-256, 
    1.8896924297306722e-258, 2.8301203067149123e-260, 
    4.1762139672168086e-262, 6.0719006273879886e-264, 
    8.6982250257053972e-266, 1.2277238484593332e-267, 
    1.7073981836665045e-269, 2.3395536450640561e-271, 
    3.1586046497952372e-273, 4.2016667376437636e-275, 
    5.5069610482308847e-277, 7.1115861655226747e-279, 
    9.0486755819602377e-281, 1.1344036865505223e-282, 
    1.4012457559161842e-284, 1.7053952969945372e-286, 
    2.0450309330144292e-288, 2.4162327791986835e-290, 
    2.8128186426399482e-292, 3.2263298152102294e-294, 
    3.6461947473000952e-296, 4.0600841072516216e-298, 
    4.4544518556700546e-300, 4.8152360102394827e-302, 
    5.1286723740060519e-304, 5.3821575300345176e-306, 
    5.5650865495734418e-308, 5.6695881332244625e-310, 
    5.6910862600134632e-312, 5.6286325200651865e-314, 
    5.4849754973548085e-316, 5.2663593541203904e-318, 
    4.9821579726631302e-320, 4.6442170709077175e-322, 
    4.9406564584124654e-324, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Sqw-Na =
  // Sqw-Na(0, 0-1999)
    0.16264072692879217, 0.16163257848253348, 0.15864830524097015, 
    0.15380570101777902, 0.14729227422649277, 0.1393529049829865, 
    0.13027421238165435, 0.12036703785866419, 0.10994854774441158, 
    0.099325389898964125, 0.088779125206158091, 0.078554831919026888, 
    0.068853397569099167, 0.05982762052057522, 0.051581887789100937, 
    0.044174913331709552, 0.037624833261251663, 0.031915867747493928, 
    0.027005766431617083, 0.022833337302982808, 0.019325494364034173, 
    0.016403421526530165, 0.013987615589680959, 0.012001721148744262, 
    0.010375192330736877, 0.0090449041687208076, 0.0079558896245315331, 
    0.0070614004092815832, 0.0063224871289086935, 0.0057072743011411008, 
    0.0051900757016506514, 0.0047504615294206264, 0.0043723557698662763, 
    0.0040432129985164961, 0.0037533003457054397, 0.0034950928787026393, 
    0.0032627788560909443, 0.0030518642765093923, 0.0028588627781215735, 
    0.0026810561490415719, 0.0025163115241599011, 0.002362943016592504, 
    0.0022196075258861031, 0.0020852264394558718, 0.0019589267136818551, 
    0.0018399963127058981, 0.0017278501915436709, 0.0016220039669631238, 
    0.001522053168610509, 0.001427656546725377, 0.0013385223662748873, 
    0.0012543969661180524, 0.0011750551238691907, 0.0011002919554563425, 
    0.0010299162034266575, 0.00096374483964920985, 0.00090159893628688167, 
    0.00084330075437357571, 0.00078867197286897398, 0.00073753294321786725, 
    0.00068970281480533067, 0.00064500034338050584, 0.00060324517361416143, 
    0.00056425938223462048, 0.00052786908090270536, 0.00049390590692964759, 
    0.00046220827168717198, 0.00043262228602611557, 0.00040500233317873797, 
    0.00037921130639832328, 0.00035512056572562363, 0.00033260969209477205, 
    0.00031156612589054326, 0.00029188477166745223, 0.00027346763365601004, 
    0.00025622352201122166, 0.00024006784231879317, 0.00022492245540425986, 
    0.00021071557490092102, 0.0001973816588974677, 0.0001848612502577813, 
    0.00017310072727418354, 0.00016205194025493142, 0.00015167172769201142, 
    0.00014192132468821879, 0.00013276569339274922, 0.00012417281789467864, 
    0.00011611301277335089, 0.00010855829464474789, 0.00010148185983642885, 
    9.4857699815077202e-05, 8.8660370826504318e-05, 8.2864917386790365e-05, 
    7.7446932903463197e-05, 7.2382726781161552e-05, 6.7649557508543077e-05, 
    6.3225886517836007e-05, 5.909160849437447e-05, 5.5228220013136196e-05, 
    5.1618898958375329e-05, 4.8248480650193816e-05, 4.5103331137022437e-05, 
    4.2171131789946984e-05, 3.9440600417947242e-05, 3.6901181281536682e-05, 
    3.4542738894707059e-05, 3.2355288316079234e-05, 3.0328788354086857e-05, 
    2.8453014883469911e-05, 2.6717520769670902e-05, 2.5111678285035699e-05, 
    2.362479079428225e-05, 2.2246253950661644e-05, 2.0965743272646359e-05, 
    1.9773404834604647e-05, 1.8660028509518935e-05, 1.7617187992257118e-05, 
    1.6637337762149264e-05, 1.5713863239073085e-05, 1.4841085809203355e-05, 
    1.401422854167139e-05, 1.3229350986358418e-05, 1.2483262427337687e-05, 
    1.1773422606697655e-05, 1.1097837626670552e-05, 1.0454956945832788e-05, 
    9.8435755348879621e-06, 9.2627436786713707e-06, 8.7116857852452672e-06, 
    8.1897289313576323e-06, 7.696241644910662e-06, 7.2305834370203447e-06, 
    6.7920656518965519e-06, 6.3799241390100485e-06, 5.9933039602043999e-06, 
    5.6312558074513229e-06, 5.2927430816839639e-06, 4.9766577956078203e-06, 
    4.6818427633988492e-06, 4.4071170767439933e-06, 4.1513017433762254e-06, 
    3.9132426258744412e-06, 3.6918284331876573e-06, 3.4860023923829978e-06, 
    3.294767220538698e-06, 3.117183972082918e-06, 2.9523661081286031e-06, 
    2.7994706216760577e-06, 2.6576882040465809e-06, 2.5262342714338308e-06, 
    2.4043422475198572e-06, 2.2912599248189876e-06, 2.1862491136169302e-06, 
    2.088588242108871e-06, 1.9975771677728278e-06, 1.9125432418757164e-06, 
    1.8328476346935284e-06, 1.7578910512970481e-06, 1.6871181937481541e-06, 
    1.6200206020138964e-06, 1.5561377777890878e-06, 1.4950567285461269e-06, 
    1.4364102379812757e-06, 1.3798742701413283e-06, 1.3251649492124918e-06, 
    1.2720355374277117e-06, 1.2202737694552978e-06, 1.1696998061152002e-06, 
    1.1201649497671718e-06, 1.0715511314250923e-06, 1.0237710431244339e-06, 
    9.7676866510927133e-07, 9.3051983809929946e-07, 8.850324751639291e-07, 
    8.4034600351368094e-07, 7.9652968325010407e-07, 7.5367956080246276e-07, 
    7.1191396903692076e-07, 6.7136766094700533e-07, 6.3218483548480164e-07, 
    5.9451145569821162e-07, 5.5848735207609659e-07, 5.2423863469905011e-07, 
    4.918709071649597e-07, 4.6146369040841038e-07, 4.3306634508658776e-07, 
    4.0669564520913009e-07, 3.8233502648814279e-07, 3.5993542363930336e-07, 
    3.3941753350694615e-07, 3.2067529389463536e-07, 3.0358034884818413e-07, 
    2.8798726768087818e-07, 2.7373928836375806e-07, 2.606743559371359e-07, 
    2.4863121920095422e-07, 2.3745533438564102e-07, 2.2700430863288038e-07, 
    2.1715260700556404e-07, 2.0779525497315452e-07, 1.9885030152162628e-07, 
    1.9025987025577935e-07, 1.8198971617593746e-07, 1.7402731719862969e-07, 
    1.663786499940158e-07, 1.5906391502040607e-07, 1.5211256976803961e-07, 
    1.4555809009313585e-07, 1.3943289664613182e-07, 1.3376385525077894e-07, 
    1.2856868838591681e-07, 1.2385353017036809e-07, 1.1961173144454013e-07, 
    1.1582389213896391e-07, 1.1245897973736687e-07, 1.0947630020045536e-07, 
    1.0682802998552604e-07, 1.044620001183413e-07, 1.0232444348244411e-07, 
    1.0036246919149325e-07, 9.8526101368389122e-08, 9.6769802613752922e-08, 
    9.5053480043969816e-08, 9.3343035092002745e-08, 9.1610557171163964e-08, 
    8.9834275185361633e-08, 8.799836954240932e-08, 8.6092718464331006e-08, 
    8.4112613548511848e-08, 8.2058442083201209e-08, 7.9935304825886133e-08, 
    7.7752525642509542e-08, 7.5523013909483722e-08, 7.3262461804575728e-08, 
    7.0988389215571508e-08, 6.8719083130187381e-08, 6.6472506257634571e-08, 
    6.4265266308839474e-08, 6.2111737419170023e-08, 6.0023409826978803e-08, 
    5.8008514440414183e-08, 5.6071933086154225e-08, 5.4215367693802213e-08, 
    5.2437711582700315e-08, 5.073554647900259e-08, 4.9103684389543702e-08, 
    4.7535682409813539e-08, 4.6024279452306953e-08, 4.4561730559602182e-08, 
    4.3140042852471218e-08, 4.1751140225903892e-08, 4.0386999192450213e-08, 
    3.9039801638474811e-08, 3.7702143785648653e-08, 3.6367323912904944e-08, 
    3.5029710339940477e-08, 3.3685167643429987e-08, 3.2331499717195678e-08, 
    3.0968854272107942e-08, 2.9600029164161917e-08, 2.823062519888494e-08, 
    2.6869003679875119e-08, 2.552602628219724e-08, 2.4214578551765745e-08, 
    2.2948901378353813e-08, 2.1743776149704485e-08, 2.0613624734609852e-08, 
    1.957159491126936e-08, 1.862870319739614e-08, 1.7793102529785414e-08, 
    1.7069530022813104e-08, 1.6458974843504615e-08, 1.5958586689454311e-08, 
    1.5561826058305581e-08, 1.5258838111544944e-08, 1.5037015679045862e-08, 
    1.4881703798298116e-08, 1.4776990379476189e-08, 1.4706523936708856e-08, 
    1.4654301684896106e-08, 1.4605377339510312e-08, 1.4546448200555613e-08, 
    1.4466293559620362e-08, 1.4356050271012631e-08, 1.4209324475017011e-08, 
    1.4022150965296082e-08, 1.3792820727745597e-08, 1.3521604476946394e-08, 
    1.3210402961988037e-08, 1.2862355979912288e-08, 1.2481439592272277e-08, 
    1.207207816976796e-08, 1.1638792571804243e-08, 1.118590185196657e-08, 
    1.0717290340998574e-08, 1.0236248764019173e-08, 9.7453935144050893e-09, 
    9.246665460979893e-09, 8.7414054023445546e-09, 8.2304998698198029e-09, 
    7.7145858297471687e-09, 7.1942983393083553e-09, 6.6705398200214513e-09, 
    6.1447457298902035e-09, 5.6191185683155749e-09, 5.0968023597402675e-09, 
    4.5819723838062789e-09, 4.0798215563053788e-09, 3.5964337173727778e-09, 
    3.1385456363987849e-09, 2.7132112393665572e-09, 2.3273930008524025e-09, 
    1.9875140921950616e-09, 1.6990103593175831e-09, 1.4659221366590354e-09, 
    1.2905627171755098e-09, 1.1732930469622912e-09, 1.1124222589287892e-09, 
    1.1042421290333812e-09, 1.1431918380084855e-09, 1.2221387115077132e-09, 
    1.3327523661027547e-09, 1.4659435674621129e-09, 1.6123362014649737e-09, 
    1.7627404204343814e-09, 1.9085971916758906e-09, 2.0423684343276672e-09, 
    2.1578521306229122e-09, 2.250407901611656e-09, 2.317085188608316e-09, 
    2.3566519728950854e-09, 2.369528407206113e-09, 2.3576341112513817e-09, 
    2.3241627361227064e-09, 2.2732999581115088e-09, 2.2099034101762752e-09, 
    2.1391638643167716e-09, 2.0662671269451393e-09, 1.9960750226325177e-09, 
    1.9328424390146308e-09, 1.8799846863737183e-09, 1.8399067844642959e-09, 
    1.8139024013127369e-09, 1.8021262993301131e-09, 1.8036396251775722e-09, 
    1.8165230987753943e-09, 1.8380484140887598e-09, 1.8648948276320069e-09, 
    1.8933943307026476e-09, 1.9197874350394556e-09, 1.9404707383098777e-09, 
    1.9522188780215301e-09, 1.9523657259952027e-09, 1.938933826607267e-09, 
    1.9107056539654908e-09, 1.8672357458254624e-09, 1.8088076492931094e-09, 
    1.7363446209727257e-09, 1.6512859872353882e-09, 1.5554437293501611e-09, 
    1.4508539237807577e-09, 1.3396369289390521e-09, 1.223877675327437e-09, 
    1.1055341527720968e-09, 9.8637806903523996e-10, 8.6796782447882832e-10, 
    7.5165008494438767e-10, 6.3858355418262768e-10, 5.2977652019831336e-10, 
    4.2612929864458675e-10, 3.2847296748666408e-10, 2.3759750926955134e-10, 
    1.5426449868264165e-10, 7.9202340595521989e-11, 1.3084520895671373e-11, 
    -4.3505793847508545e-11, -9.0120062403379232e-11, 
    -1.2649108253969106e-10, -1.5257562076746813e-10, 
    -1.6858668085857119e-10, -1.750103863435112e-10, -1.7260414005314914e-10, 
    -1.6237491156455852e-10, -1.4553854455846273e-10, 
    -1.2346333015638636e-10, -9.7602368182166071e-11, 
    -6.9420900884182669e-11, -4.0324635731177646e-11, 
    -1.1595266206309359e-11, 1.5662004736058736e-11, 4.0555257989856584e-11, 
    6.242571480021104e-11, 8.0850812200399406e-11, 9.5632739772862435e-11, 
    1.0677580246958537e-10, 1.1445679067358515e-10, 1.1899230232142253e-10, 
    1.2080671546317031e-10, 1.2040315616265553e-10, 1.1833865059957782e-10, 
    1.1520330901949069e-10, 1.1160258007197254e-10, 1.0814070254741679e-10, 
    1.0540382293040344e-10, 1.0394121990794773e-10, 1.0424427381005786e-10, 
    1.0672336801817418e-10, 1.1168421817048503e-10, 1.1930549788958144e-10, 
    1.2962039392826371e-10, 1.425043275503109e-10, 1.5767111716485829e-10, 
    1.7467876560703889e-10, 1.9294546996793794e-10, 2.1177527283415584e-10, 
    2.3039205068245363e-10, 2.4797970402627275e-10, 2.6372594204458005e-10, 
    2.7686672058862324e-10, 2.8672854843208799e-10, 2.9276584532744587e-10, 
    2.9459109874506703e-10, 2.9199598748695845e-10, 2.8496232888652536e-10, 
    2.7366230182763667e-10, 2.5844833531674772e-10, 2.3983345671714751e-10, 
    2.1846380678029976e-10, 1.9508534744717175e-10, 1.705072301452547e-10, 
    1.455642594226014e-10, 1.2108090735167219e-10, 9.7838947347400517e-11, 
    7.655015382886518e-11, 5.7835032364032758e-11, 4.2207946622051549e-11, 
    3.0068240239366635e-11, 2.1696850112631614e-11, 1.7257402031483812e-11, 
    1.6800922318670858e-11, 2.0273250815662766e-11, 2.7524611724149585e-11, 
    3.8320692172235045e-11, 5.2355217091120651e-11, 6.9263515986014304e-11, 
    8.8637076876273661e-11, 1.1003848978773684e-10, 1.3301639894575338e-10, 
    1.571196435627112e-10, 1.819098541207434e-10, 2.0697161129480933e-10, 
    2.3191962406683601e-10, 2.5640248984455549e-10, 2.8010304908856658e-10, 
    3.027357847260682e-10, 3.2404198488499656e-10, 3.4378378454478259e-10, 
    3.6173839367298849e-10, 3.7769367133307655e-10, 3.9144623894841162e-10, 
    4.0280286284828748e-10, 4.1158549394510361e-10, 4.1763979916761529e-10, 
    4.2084658494864562e-10, 4.2113493463581449e-10, 4.1849571344356997e-10, 
    4.1299367274585851e-10, 4.047766123920876e-10, 3.9408001846046146e-10, 
    3.8122615556938814e-10, 3.6661690362730053e-10, 3.5072044465643448e-10, 
    3.3405233885803e-10, 3.1715221859741394e-10, 3.0055774515231743e-10, 
    2.8477774685374702e-10, 2.7026649967986369e-10, 2.5740115194387208e-10, 
    2.4646372116670142e-10, 2.3762901024063317e-10, 2.3095896146724846e-10, 
    2.2640378105587224e-10, 2.2380936003924863e-10, 2.2293043858183999e-10, 
    2.2344832632149079e-10, 2.2499201350284313e-10, 2.271612075888363e-10, 
    2.2954983695509464e-10, 2.3176864461056854e-10, 2.3346553249600852e-10, 
    2.3434244577841725e-10, 2.3416813774708382e-10, 2.3278601548485387e-10, 
    2.3011708569515852e-10, 2.2615797095827716e-10, 2.2097467648738324e-10, 
    2.1469273455155969e-10, 2.0748483839796045e-10, 1.9955696673440476e-10, 
    1.9113414631208666e-10, 1.8244675039979665e-10, 1.7371825552414284e-10, 
    1.651548620433722e-10, 1.5693755773065247e-10, 1.4921653754719938e-10, 
    1.4210810765593552e-10, 1.3569378590591674e-10, 1.300213654716798e-10, 
    1.2510758180804318e-10, 1.2094201177886112e-10, 1.1749181823232293e-10, 
    1.1470696841023303e-10, 1.1252550848991137e-10, 1.1087862048846546e-10, 
    1.0969507570815651e-10, 1.0890493010607932e-10, 1.0844221804173686e-10, 
    1.08246633518944e-10, 1.0826417998347794e-10, 1.0844695185082823e-10, 
    1.0875219618770828e-10, 1.0914094772026353e-10, 1.0957648428551006e-10, 
    1.100229247551502e-10, 1.1044413004071618e-10, 1.108031467527919e-10, 
    1.1106226449222286e-10, 1.1118368355056469e-10, 1.1113066577857106e-10, 
    1.1086910326074116e-10, 1.103691932453622e-10, 1.096070711211595e-10, 
    1.0856607615084749e-10, 1.0723755999531218e-10, 1.0562104094657534e-10, 
    1.037236755677225e-10, 1.0155906469602793e-10, 9.9145561891246686e-11, 
    9.6504189694480303e-11, 9.3656492303744411e-11, 9.0622474514597188e-11, 
    8.7418971170051765e-11, 8.405859571779226e-11, 8.0549413854640695e-11, 
    7.6895446990517256e-11, 7.3097962643840086e-11, 6.9157368799529997e-11, 
    6.5075640497028971e-11, 6.0858914221494415e-11, 5.6519992848081668e-11, 
    5.2080427544345173e-11, 4.7571937171514398e-11, 4.3036894850032709e-11, 
    3.8527796307448289e-11, 3.4105620080496348e-11, 2.9837205256753701e-11, 
    2.5791793716363555e-11, 2.203704405185166e-11, 1.8634785276934984e-11, 
    1.5636998812857476e-11, 1.308225556535617e-11, 1.0993065293162959e-11, 
    9.374293226730507e-12, 8.2128918468824181e-12, 7.4788698196434699e-12, 
    7.1275600744228097e-12, 7.1028929154709556e-12, 7.3414358454668135e-12, 
    7.7768495678256987e-12, 8.3443975795042134e-12, 8.9850982084030325e-12, 
    9.6492643898913284e-12, 1.0299130821103168e-11, 1.0910394948356826e-11, 
    1.147267071416399e-11, 1.1988848520657034e-11, 1.2473470966344571e-11, 
    1.2950377841738236e-11, 1.3449727990857821e-11, 1.4004820752579701e-11, 
    1.4648759629124697e-11, 1.5411370563473783e-11, 1.6316433101513066e-11, 
    1.7379497453291902e-11, 1.8606300631727764e-11, 1.9992010225457815e-11, 
    2.1521209767504773e-11, 2.3168749574084733e-11, 2.4901306696192104e-11, 
    2.6679668390030006e-11, 2.8461451101450163e-11, 3.0204181514152566e-11, 
    3.1868343072141551e-11, 3.3420257688544934e-11, 3.483437674722822e-11, 
    3.6094890512784074e-11, 3.7196398255423498e-11, 3.814363630263793e-11, 
    3.8950213804061631e-11, 3.963660828834884e-11, 4.0227564077625229e-11, 
    4.0749253343276972e-11, 4.1226481027268436e-11, 4.1680313898436094e-11, 
    4.2126297238988986e-11, 4.2573553466167008e-11, 4.3024697939717599e-11, 
    4.3476660948314724e-11, 4.3922166193259763e-11, 4.4351730354111443e-11, 
    4.4755801147496509e-11, 4.5126895956280863e-11, 4.5461316053688928e-11, 
    4.5760372722217242e-11, 4.6030872003272702e-11, 4.6284919771275614e-11, 
    4.6538970738980814e-11, 4.6812352265541842e-11, 4.7125338214794281e-11, 
    4.749707032729074e-11, 4.7943445785338983e-11, 4.8475261204458285e-11, 
    4.9096695314532645e-11, 4.9804343205777428e-11, 5.0586770239077266e-11, 
    5.142470755973527e-11, 5.2291784058206112e-11, 5.3155830344505891e-11, 
    5.3980531256579458e-11, 5.4727479043151285e-11, 5.5358376193885012e-11, 
    5.5837343866216244e-11, 5.6133105972501764e-11, 5.6220993020681382e-11, 
    5.6084604804587709e-11, 5.5717004306674626e-11, 5.5121331462591127e-11, 
    5.4310877066633954e-11, 5.3308462258480421e-11, 5.2145296681148578e-11, 
    5.0859303044210882e-11, 4.9493052420405395e-11, 4.80914808434743e-11, 
    4.6699528137148714e-11, 4.5359839403807503e-11, 4.4110740123402207e-11, 
    4.2984547341145335e-11, 4.2006348136674481e-11, 4.1193253445084451e-11, 
    4.0554159495597304e-11, 4.0090019045574768e-11, 3.979450695634121e-11, 
    3.965502158991759e-11, 3.9653958726023878e-11, 3.9770120141831303e-11, 
    3.9980171285641721e-11, 4.0260025097019329e-11, 4.058608828415792e-11, 
    4.0936301525485406e-11, 4.1290893443829695e-11, 4.1632839177019792e-11, 
    4.1948027783099369e-11, 4.2225149045349231e-11, 4.2455394059169701e-11, 
    4.2631947272184141e-11, 4.274946689235216e-11, 4.2803577718162215e-11, 
    4.2790472246920686e-11, 4.2706655511485266e-11, 4.2548889772097695e-11, 
    4.2314382986155482e-11, 4.2001120193443396e-11, 4.1608297785735095e-11, 
    4.1136837817974489e-11, 4.0589803459590461e-11, 3.9972731007002929e-11, 
    3.9293704949946539e-11, 3.8563234520249016e-11, 3.7793831571619467e-11, 
    3.6999408930236068e-11, 3.6194437552532069e-11, 3.5393089264093476e-11, 
    3.4608303462165583e-11, 3.3850999793050035e-11, 3.3129447186387286e-11, 
    3.2448867069339475e-11, 3.1811288503553751e-11, 3.1215704735820212e-11, 
    3.065840816109144e-11, 3.0133558422990182e-11, 2.9633838824079013e-11, 
    2.9151178501811069e-11, 2.8677404426112311e-11, 2.8204872459452009e-11, 
    2.772691023021855e-11, 2.7238169337188849e-11, 2.6734767993278382e-11, 
    2.6214345477510249e-11, 2.5675964047098202e-11, 2.5119973108906419e-11, 
    2.454777261038781e-11, 2.3961621354780187e-11, 2.3364409373081178e-11, 
    2.2759521571759623e-11, 2.2150667275586892e-11, 2.1541820679776531e-11, 
    2.0937139033293868e-11, 2.0340927380563168e-11, 1.975759638838682e-11, 
    1.9191652728255463e-11, 1.8647590049873494e-11, 1.8129855410721831e-11, 
    1.7642728240288075e-11, 1.7190242410951899e-11, 1.6776020369304519e-11, 
    1.6403188385390405e-11, 1.6074255684718562e-11, 1.5791019242675474e-11, 
    1.5554478727458016e-11, 1.5364792927639646e-11, 1.5221236537177296e-11, 
    1.5122208639274433e-11, 1.5065236925272726e-11, 1.5047025074214451e-11, 
    1.5063505435623194e-11, 1.5109929019568358e-11, 1.5180943454831697e-11, 
    1.5270732453156703e-11, 1.5373150233279877e-11, 1.5481888356999839e-11, 
    1.5590701080038657e-11, 1.5693622786566367e-11, 1.5785269480446582e-11, 
    1.5861122266469196e-11, 1.5917816905739533e-11, 1.5953450543614434e-11, 
    1.5967789123147122e-11, 1.596242759635355e-11, 1.5940822078339234e-11, 
    1.5908157038497124e-11, 1.5871093202353636e-11, 1.5837325244931673e-11, 
    1.5815031074901073e-11, 1.5812228333813333e-11, 1.5836073546525477e-11, 
    1.589223176138545e-11, 1.5984315700119424e-11, 1.6113490710139268e-11, 
    1.6278306340224865e-11, 1.6474780916807182e-11, 1.6696641196621753e-11, 
    1.6935845935215503e-11, 1.7183251309676697e-11, 1.7429359720171798e-11, 
    1.7665082598930708e-11, 1.7882460764116533e-11, 1.8075225405345083e-11, 
    1.8239215307734022e-11, 1.8372555890078759e-11, 1.8475633550330425e-11, 
    1.855084513358636e-11, 1.8602195277838581e-11, 1.8634759609048017e-11, 
    1.8654089174579383e-11, 1.8665593164037338e-11, 1.8674032027033732e-11, 
    1.8683022726757506e-11, 1.8694744096681572e-11, 1.8709791944726801e-11, 
    1.8727202942784334e-11, 1.8744570842340484e-11, 1.8758390126051824e-11, 
    1.8764421178621987e-11, 1.875814662486949e-11, 1.8735250385741131e-11, 
    1.8692080409321894e-11, 1.862599933154184e-11, 1.8535732466439415e-11, 
    1.8421504268517902e-11, 1.8285131021181145e-11, 1.8129939368243121e-11, 
    1.7960608048857592e-11, 1.7782883154327958e-11, 1.7603233953859344e-11, 
    1.7428478427170194e-11, 1.7265372663206312e-11, 1.7120204002595447e-11, 
    1.6998442040001574e-11, 1.6904395463465738e-11, 1.684097500453896e-11, 
    1.6809457782701077e-11, 1.6809377518912858e-11, 1.6838480554375518e-11, 
    1.6892749761684041e-11, 1.6966530221664339e-11, 1.7052750856900846e-11, 
    1.7143218774525676e-11, 1.7229048832092222e-11, 1.7301097004865348e-11, 
    1.7350524510591679e-11, 1.7369316483665606e-11, 1.7350829787957318e-11, 
    1.7290222961170212e-11, 1.7184855234221425e-11, 1.7034464738275647e-11, 
    1.6841222704764184e-11, 1.6609578275401423e-11, 1.6345958767781668e-11, 
    1.6058268011765267e-11, 1.5755327713072103e-11, 1.5446251502952792e-11, 
    1.5139808846481507e-11, 1.4843886652913127e-11, 1.4565052474645025e-11, 
    1.430825176455145e-11, 1.4076705683236858e-11, 1.3871925358013447e-11, 
    1.3693907757997095e-11, 1.3541386908916996e-11, 1.3412157387085549e-11, 
    1.3303410729614715e-11, 1.3212029152412274e-11, 1.313480130470627e-11, 
    1.306860044515804e-11, 1.3010431298008221e-11, 1.2957461240018447e-11, 
    1.2906986017652201e-11, 1.285637291231432e-11, 1.2803048151065244e-11, 
    1.2744470232607283e-11, 1.2678194116831173e-11, 1.2601956192600687e-11, 
    1.2513808605062129e-11, 1.2412267070492276e-11, 1.2296499192976061e-11, 
    1.2166445132666915e-11, 1.20229621088225e-11, 1.1867865211468011e-11, 
    1.1703948723128366e-11, 1.1534900457585095e-11, 1.1365203814892231e-11, 
    1.1199914217219612e-11, 1.1044446567767931e-11, 1.0904286750659304e-11, 
    1.0784697291228809e-11, 1.0690402723584993e-11, 1.0625302285542441e-11, 
    1.0592218401267003e-11, 1.0592655743557556e-11, 1.0626668215356941e-11, 
    1.0692794138608283e-11, 1.0788066925840631e-11, 1.09081400733499e-11, 
    1.104748972121088e-11, 1.1199678723037328e-11, 1.1357707113223118e-11, 
    1.151434876652367e-11, 1.1662506338735526e-11, 1.1795531295238234e-11, 
    1.1907454976545937e-11, 1.1993191915226202e-11, 1.2048630011018802e-11, 
    1.2070633147494133e-11, 1.2057010128913096e-11, 1.2006438633359283e-11, 
    1.1918378456663068e-11, 1.1792977259966118e-11, 1.1631044226431e-11, 
    1.1434028950488677e-11, 1.120407905838919e-11, 1.0944087469962116e-11, 
    1.0657797545459145e-11, 1.0349825868729031e-11, 1.0025732712401871e-11, 
    9.6919378618208633e-12, 9.3556318104718715e-12, 9.0245631241352423e-12, 
    8.7067897131209309e-12, 8.4103197365353918e-12, 8.1427757464342588e-12, 
    7.9110074824868368e-12, 7.7207730873476269e-12, 7.5764188354212118e-12, 
    7.4806790130586137e-12, 7.4345264642756117e-12, 7.4371478464583669e-12, 
    7.4859576969409011e-12, 7.5767379427734871e-12, 7.7037977878598756e-12, 
    7.8602471223373934e-12, 8.0382250854895849e-12, 8.2292043642628425e-12, 
    8.4243093293184665e-12, 8.6146290955236975e-12, 8.7915253767226121e-12, 
    8.9469656097728999e-12, 9.0738078920762561e-12, 9.1661288041269725e-12, 
    9.2194573275822439e-12, 9.2310122373647301e-12, 9.1998731481183409e-12, 
    9.1270693549303566e-12, 9.0155709265985086e-12, 8.8701991321786096e-12, 
    8.6974099538062318e-12, 8.5049890261354281e-12, 8.3016539879684041e-12, 
    8.0966031474855424e-12, 7.899010527617566e-12, 7.7175524559863652e-12, 
    7.5599404763006152e-12, 7.4325428835156909e-12, 7.3400977737539184e-12, 
    7.285553789218727e-12, 7.2700014086085683e-12, 7.292757880091159e-12, 
    7.3515263606005827e-12, 7.4426519084399256e-12, 7.5614083528782828e-12, 
    7.7023228463642535e-12, 7.8594769056274222e-12, 8.026784715036005e-12, 
    8.1982271886199051e-12, 8.3680337500572402e-12, 8.5308040404228486e-12, 
    8.6815922804213741e-12, 8.8159664259786714e-12, 8.9300548026316843e-12, 
    9.020556762826949e-12, 9.0847939067105309e-12, 9.1207525931437145e-12, 
    9.1271199904523017e-12, 9.103352104605324e-12, 9.0497314348221216e-12, 
    8.9673743261391792e-12, 8.8582714733846572e-12, 8.7252426273633451e-12, 
    8.5719171141605284e-12, 8.4026056754558014e-12, 8.2222042597187448e-12, 
    8.0360133003336217e-12, 7.8496038400696755e-12, 7.6685647811420121e-12, 
    7.4983442404720674e-12, 7.344018369430321e-12, 7.2101210034552729e-12, 
    7.100427856626778e-12, 7.0178325486879401e-12, 6.9641670675959121e-12, 
    6.9401452173729809e-12, 6.9452606074744405e-12, 6.9778356366548448e-12, 
    7.0350092709261003e-12, 7.1128890963561756e-12, 7.2066822697054659e-12, 
    7.3109430504200204e-12, 7.4198004105891055e-12, 7.5272608266683442e-12, 
    7.6275006568865277e-12, 7.7151509701914554e-12, 7.7855566173322694e-12, 
    7.834994137795061e-12, 7.8608215703030481e-12, 7.8615796017945989e-12, 
    7.8370128588047544e-12, 7.7880436647976292e-12, 7.7166654623654707e-12, 
    7.6258236971910191e-12, 7.519236306762063e-12, 7.4012094052144708e-12, 
    7.2764187350081046e-12, 7.1497146788280587e-12, 7.0258966311206812e-12, 
    6.909487965120891e-12, 6.8045556660090619e-12, 6.7145240160178681e-12, 
    6.6419725963640595e-12, 6.588512745787599e-12, 6.5546735207651051e-12, 
    6.5398481222930114e-12, 6.5422512415067201e-12, 6.5590047341118025e-12, 
    6.5862145102830544e-12, 6.6191500504083107e-12, 6.6524636325795607e-12, 
    6.6804739514384957e-12, 6.6974437013692669e-12, 6.6979251881944997e-12, 
    6.6770659902507694e-12, 6.630916530003743e-12, 6.55669696557621e-12, 
    6.4530319981618657e-12, 6.320074179071806e-12, 6.1595903107524697e-12, 
    5.9749442220488514e-12, 5.7710053950994559e-12, 5.5539343045585116e-12, 
    5.3309370983911489e-12, 5.1099199579766566e-12, 4.8990945705267015e-12, 
    4.7065800047342381e-12, 4.5399587800621524e-12, 4.4058697483521701e-12, 
    4.3096587269871125e-12, 4.2550601742578905e-12, 4.2439823671558782e-12, 
    4.2763686219968799e-12, 4.3501760024075121e-12, 4.4614587988934872e-12, 
    4.6045718990378629e-12, 4.7724521871593607e-12, 4.9570207488631225e-12, 
    5.1496282521759026e-12, 5.3415550062388341e-12, 5.524541539950003e-12, 
    5.6912601549759339e-12, 5.835782748229022e-12, 5.9539205907228012e-12, 
    6.0434555120655775e-12, 6.1042129632371258e-12, 6.1380076386368441e-12, 
    6.1483949993461528e-12, 6.1403123602277e-12, 6.119572578861865e-12, 
    6.0923311224057992e-12, 6.0645030503103507e-12, 6.0412333671896278e-12, 
    6.0264513193064391e-12, 6.0225779762520405e-12, 6.0303703566620033e-12, 
    6.0489696472406394e-12, 6.0760858131013339e-12, 6.1083534198408219e-12, 
    6.1417577666127992e-12, 6.1721137489482522e-12, 6.1955340272269139e-12, 
    6.2088261198867157e-12, 6.2097761599012877e-12, 6.1973113928806657e-12, 
    6.1714971681551149e-12, 6.1334208395481016e-12, 6.0849490697876342e-12, 
    6.0284180214193415e-12, 5.9662999241340894e-12, 5.9008792151591483e-12, 
    5.8339994500967317e-12, 5.7668884342834312e-12, 5.7001073407123726e-12, 
    5.6336052854095053e-12, 5.5668507799924949e-12, 5.4990870312404283e-12, 
    5.4296026468484888e-12, 5.3579543347586858e-12, 5.2842266403326041e-12, 
    5.2091618444502125e-12, 5.1342161145613774e-12, 5.0614958710818504e-12, 
    4.9936023811926131e-12, 4.9333759634788723e-12, 4.8836086586230098e-12, 
    4.8467218382171676e-12, 4.8244851948239547e-12, 4.8177827840448901e-12, 
    4.826472021395975e-12, 4.8493471793198249e-12, 4.8842268576784275e-12, 
    4.9280952140321708e-12, 4.9773696941458244e-12, 5.0281714568954572e-12, 
    5.0766311008824593e-12, 5.1191707345982229e-12, 5.1527269667779809e-12, 
    5.1749391854184195e-12, 5.1842310331564158e-12, 5.1798513540241634e-12, 
    5.1618312776784346e-12, 5.130892964635903e-12, 5.0883269560329294e-12, 
    5.0358621491191532e-12, 4.9755022259543758e-12, 4.9094068069697349e-12, 
    4.8397396124893928e-12, 4.7685618359465264e-12, 4.6977256039123853e-12, 
    4.6287791503611216e-12, 4.5628802615495644e-12, 4.5007416528583022e-12, 
    4.4425856950676903e-12, 4.3881014087753239e-12, 4.3364737603822934e-12, 
    4.2864243668935665e-12, 4.2362984309025899e-12, 4.1842063707153485e-12, 
    4.1281683307576856e-12, 4.0663349035770021e-12, 3.9971636462542725e-12, 
    3.9196270264329925e-12, 3.8333753277652499e-12, 3.7388422435829133e-12, 
    3.6373090290170466e-12, 3.5308936119605076e-12, 3.4224530141899691e-12, 
    3.3154594414346273e-12, 3.2137934274949215e-12, 3.1215252740152694e-12, 
    3.0426739364935904e-12, 2.9809786839532355e-12, 2.9396851785250888e-12, 
    2.9213741284285195e-12, 2.9278531748939974e-12, 2.9600284671399378e-12, 
    3.0179047980614278e-12, 3.1005685876099358e-12, 3.2062319001358184e-12, 
    3.3323004706052683e-12, 3.4754992479354253e-12, 3.6319777947055311e-12, 
    3.7974855646648945e-12, 3.9675553238335835e-12, 4.1377187004287796e-12, 
    4.3036930993643941e-12, 4.4616110590489999e-12, 4.6081883432455277e-12, 
    4.7408985649540204e-12, 4.8580351203413824e-12, 4.9587360397349451e-12, 
    5.0429449340474002e-12, 5.1112627046527465e-12, 5.1647544327019719e-12, 
    5.2047056379134924e-12, 5.2323550133438911e-12, 5.2486528553095099e-12, 
    5.2540522629208967e-12, 5.2483753025997087e-12, 5.2307841966847874e-12, 
    5.1998339822544967e-12, 5.1536254332594084e-12, 5.0900701387651203e-12, 
    5.0071600408112717e-12, 4.9032859284717343e-12, 4.7775649512408518e-12, 
    4.6300717379014274e-12, 4.4620261759668569e-12, 4.2758638331352661e-12, 
    4.0751988239034642e-12, 3.8646340153217863e-12, 3.6495447609528307e-12, 
    3.4357180169503887e-12, 3.2289578689489165e-12, 3.0346738932434751e-12, 
    2.8575156828587054e-12, 2.701033881196925e-12, 2.5674655091564079e-12, 
    2.4576096967049441e-12, 2.3708499388026193e-12, 2.3052775654369353e-12, 
    2.2579631308506897e-12, 2.2252746880478356e-12, 2.2032668837477867e-12, 
    2.1880514289247662e-12, 2.1761871717456399e-12, 2.1649493690659663e-12, 
    2.152529333393108e-12, 2.1381054331019298e-12, 2.1218264768348131e-12, 
    2.1046610230863615e-12, 2.0881723155379328e-12, 2.0742258094898661e-12, 
    2.0647016950858634e-12, 2.0611621089619099e-12, 2.0646232768204614e-12, 
    2.0753371144343876e-12, 2.0927116609915085e-12, 2.1152720215640703e-12, 
    2.1407853643134016e-12, 2.166396743857742e-12, 2.1889345621928977e-12, 
    2.2051818596652084e-12, 2.2122327225147974e-12, 2.2078173734802114e-12, 
    2.1906038106313172e-12, 2.1604059285558594e-12, 2.1183560237238497e-12, 
    2.0669008307738569e-12, 2.009738900737146e-12, 1.951583022897179e-12, 
    1.8978987275735308e-12, 1.8544753911416745e-12, 1.8270432564670613e-12, 
    1.8207857826903114e-12, 1.8399908418691698e-12, 1.8876584322473275e-12, 
    1.9653015559630786e-12, 2.0727986382192511e-12, 2.2083986887300755e-12, 
    2.3688419768250595e-12, 2.5495934126118477e-12, 2.7451542886166679e-12, 
    2.9494313615892583e-12, 3.1561160530721926e-12, 3.3590720509267793e-12, 
    3.5526448369863948e-12, 3.7319588691325481e-12, 3.893079586041931e-12, 
    4.0331332021628669e-12, 4.1502963125098907e-12, 4.2437599505424742e-12, 
    4.313563073929786e-12, 4.360437520019059e-12, 4.3855650080318052e-12, 
    4.3903662296622713e-12, 4.37624950214294e-12, 4.3444379955419659e-12, 
    4.2957992703635847e-12, 4.2307377756392439e-12, 4.1491715265337115e-12, 
    4.0505767705693242e-12, 3.9340919988985143e-12, 3.7987261684493569e-12, 
    3.643585636319239e-12, 3.4681556798038873e-12, 3.2725837573307475e-12, 
    3.0579177151800784e-12, 2.8263152127301049e-12, 2.5811409153490707e-12, 
    2.3269698136050119e-12, 2.0694655335500057e-12, 1.8151493975635771e-12, 
    1.571058826362618e-12, 1.344348344060464e-12, 1.1418259821009989e-12, 
    9.6953339323593325e-13, 8.3232885055917429e-13, 7.3357363362935459e-13, 
    6.7491441828666115e-13, 6.5623303362405415e-13, 6.7564000837968427e-13, 
    7.2969143308006623e-13, 8.1360264910826911e-13, 9.216474909747129e-13, 
    1.047479618986123e-12, 1.1845810796362678e-12, 1.3265792123780104e-12, 
    1.4676359854514544e-12, 1.602647970706989e-12, 1.7275114323845297e-12, 
    1.8391667830731914e-12, 1.9357082560407298e-12, 2.0163075424537748e-12, 
    2.0811744727446362e-12, 2.1313953818594398e-12, 2.1688206545233382e-12, 
    2.195836839550751e-12, 2.2152358225351421e-12, 2.229970588546919e-12, 
    2.2430354420750155e-12, 2.2572499832486555e-12, 2.2751468246673303e-12, 
    2.2988253723339205e-12, 2.3298792417309029e-12, 2.3692681064316239e-12, 
    2.4173139402494665e-12, 2.4736511687068632e-12, 2.5372460637383205e-12, 
    2.6064381667525506e-12, 2.6790264108045816e-12, 2.7523733615092842e-12, 
    2.8235907546843841e-12, 2.8896962294731172e-12, 2.9478498184181603e-12, 
    2.9955524751493827e-12, 3.0308734190417429e-12, 3.0526195444096195e-12, 
    3.0604913395759002e-12, 3.0551360572590733e-12, 3.0381570831242077e-12, 
    3.0120239022515733e-12, 2.9799201990615157e-12, 2.9454844526218061e-12, 
    2.912564569363032e-12, 2.8848722002736062e-12, 2.8656963019549999e-12, 
    2.8576051689734832e-12, 2.862242058129183e-12, 2.8801460725781381e-12, 
    2.9107095178634944e-12, 2.9521909033056685e-12, 3.0018637360333862e-12, 
    3.0561891784347565e-12, 3.1111021748965943e-12, 3.1623189555928933e-12, 
    3.2056600493481424e-12, 3.2373629396553301e-12, 3.2543810070316817e-12, 
    3.2545925753924153e-12, 3.2369678070477085e-12, 3.2016342970763536e-12, 
    3.1498657236016574e-12, 3.0839641442094248e-12, 3.007094690226196e-12, 
    2.9230212913706117e-12, 2.8358266213377561e-12, 2.7496055730094794e-12, 
    2.6681617748058174e-12, 2.5947298533599528e-12, 2.5317608993723979e-12, 
    2.4807586004337226e-12, 2.4422227708681412e-12, 2.4156347394193153e-12, 
    2.3995653708506607e-12, 2.391817850875549e-12, 2.3896675855544955e-12, 
    2.3900845871964781e-12, 2.3900084004776497e-12, 2.3865963018134055e-12, 
    2.3774550209766713e-12, 2.3607829834028081e-12, 2.335500124353467e-12, 
    2.3012757808506219e-12, 2.2585119545025942e-12, 2.2082491788796737e-12, 
    2.1520458653864786e-12, 2.0918248415591956e-12, 2.0297084786343898e-12, 
    1.9678588105580794e-12, 1.9083689475265475e-12, 1.8531307091285623e-12, 
    1.8037839830568723e-12, 1.7616778960614898e-12, 1.7278695113977321e-12, 
    1.7031157307015024e-12, 1.687913997425064e-12, 1.6825055086305902e-12, 
    1.6869071190701882e-12, 1.7009380145592363e-12, 1.7241777267816759e-12, 
    1.7560398605602768e-12, 1.7957700920699677e-12, 1.842450009280847e-12, 
    1.8950469448438742e-12, 1.9524234258011125e-12, 2.0133887262027988e-12, 
    2.0766985433601019e-12, 2.1411091689182889e-12, 2.2053350005965304e-12, 
    2.2680662543418536e-12, 2.3279211736134598e-12, 2.38343102446005e-12, 
    2.432983180545867e-12, 2.4748239230394838e-12, 2.5070520231373285e-12, 
    2.5276729825664751e-12, 2.5346775079839808e-12, 2.5261706339563016e-12, 
    2.500520291843971e-12, 2.456554690543113e-12, 2.3937037228367792e-12, 
    2.3121822083439514e-12, 2.2130596961788356e-12, 2.0983289616350169e-12, 
    1.9708248201439803e-12, 1.8341331019703242e-12, 1.6923562608095489e-12, 
    1.5498556389080978e-12, 1.4109420608098071e-12, 1.2795714891199813e-12, 
    1.1590439857204115e-12, 1.0517740954850491e-12, 9.591409579772618e-13, 
    8.8142391771340793e-13, 8.178552039344173e-13, 7.667477403257196e-13, 
    7.2572283297579823e-13, 6.9198481360513359e-13, 6.6261895760273965e-13, 
    6.3490038236264897e-13, 6.0657344055890792e-13, 5.7605789855036948e-13, 
    5.4263144552474297e-13, 5.0649291003203602e-13, 4.6876707668956836e-13, 
    4.3142989646226177e-13, 3.9718049834955073e-13, 3.6923598042357927e-13, 
    3.5112136496410011e-13, 3.4641734598995061e-13, 3.5850751852951753e-13, 
    3.9035134457663178e-13, 4.4425918363017435e-13, 5.2174177980093898e-13, 
    6.233634857808742e-13, 7.486969678471883e-13, 8.9631247346024798e-13, 
    1.0638314713440137e-12, 1.2480364670565821e-12, 1.4450516610791373e-12, 
    1.6504882576726583e-12, 1.8596835012007246e-12, 2.067886401956894e-12, 
    2.2704520079975253e-12, 2.4629930424036583e-12, 2.6415037458917725e-12, 
    2.802435523520815e-12, 2.9427598570907253e-12, 3.0599634301089463e-12, 
    3.1520714633258489e-12, 3.2176268057381528e-12, 3.2557027472366589e-12, 
    3.2659065042244883e-12, 3.2484329515366239e-12, 3.2040779236339736e-12, 
    3.1343221928480821e-12, 3.0413423619558026e-12, 2.9280684914408423e-12, 
    2.798156607716513e-12, 2.6559592515994962e-12, 2.5064005259606639e-12, 
    2.3548313370617566e-12, 2.2068082330690125e-12, 2.067865562867246e-12, 
    1.9432012750922201e-12, 1.8374478026737676e-12, 1.7543607381137394e-12, 
    1.6966178416144003e-12, 1.6656666106159515e-12, 1.661659792960605e-12, 
    1.6834254755072255e-12, 1.728578341652946e-12, 1.7937014124003002e-12, 
    1.8745837931539213e-12, 1.9664815195407836e-12, 2.0644413188142804e-12, 
    2.1635871260601624e-12, 2.2593773963503302e-12, 2.3478422987784812e-12, 
    2.4257304336104124e-12, 2.4906099076304624e-12, 2.5408901813243017e-12, 
    2.5758066132036546e-12, 2.5953504980667603e-12, 2.6001623075417629e-12, 
    2.5914067676914759e-12, 2.5706594114389195e-12, 2.5397674694204119e-12, 
    2.5007417314966716e-12, 2.4556414485623571e-12, 2.4064785419407523e-12, 
    2.3551344316679211e-12, 2.3032834356721144e-12, 2.2523184737583766e-12, 
    2.2033064649920898e-12, 2.1569364513294669e-12, 2.1135059852345272e-12, 
    2.072933297377564e-12, 2.0347565283642374e-12, 1.998217848185248e-12, 
    1.9623095699500443e-12, 1.9259065035175426e-12, 1.8878510265069361e-12, 
    1.8470798090686974e-12, 1.8027223034952098e-12, 1.7542047964983511e-12, 
    1.7012866923896866e-12, 1.6441094324274234e-12, 1.5831762425610436e-12, 
    1.5193401669722222e-12, 1.4537096112502951e-12, 1.3875915484874619e-12, 
    1.3223928160775052e-12, 1.2595525884093077e-12, 1.2004573614773554e-12, 
    1.1464089705753036e-12, 1.0985719180128316e-12, 1.0580037245153389e-12, 
    1.0256141406220891e-12, 1.0021946642181243e-12, 9.8841443611964333e-13, 
    9.8480356360666107e-13, 9.9170651646178965e-13, 1.0092385204392484e-12, 
    1.037175317416857e-12, 1.0748784985191313e-12, 1.1211999778310348e-12, 
    1.1744189710506273e-12, 1.2322007263102997e-12, 1.291631953791459e-12, 
    1.3493053735160067e-12, 1.4014756881349663e-12, 1.444265612458982e-12, 
    1.4739373262462877e-12, 1.4871576774548258e-12, 1.4812877630556931e-12, 
    1.4546145236761584e-12, 1.4065674955739921e-12, 1.337791410922579e-12, 
    1.2501649903735898e-12, 1.1467473950912466e-12, 1.0315933434661964e-12, 
    9.0949136287476126e-13, 7.8566991640795126e-13, 6.6545801105746965e-13, 
    5.539466903479381e-13, 4.5565299175331605e-13, 3.7426843691954508e-13, 
    3.124265060446082e-13, 2.7158030505527171e-13, 2.5194121371249701e-13, 
    2.5251430573767073e-13, 2.7119237548263473e-13, 3.0495695558138841e-13, 
    3.5007045918721955e-13, 4.0236952811410823e-13, 4.5752756965534371e-13, 
    5.1136677463620434e-13, 5.6009723855921227e-13, 6.005909348972859e-13, 
    6.3053127513672236e-13, 6.485866725258455e-13, 6.5444221002806752e-13, 
    6.48823606172552e-13, 6.3338821964996329e-13, 6.1060331908655451e-13, 
    5.8351527891442043e-13, 5.5554083195610059e-13, 5.3015170072981825e-13, 
    5.1063089283898276e-13, 4.9979899405679452e-13, 4.9982500852718647e-13, 
    5.120451316327915e-13, 5.3689252290741207e-13, 5.7390421651270931e-13, 
    6.2177320707130474e-13, 6.7853076565704999e-13, 7.4170266665182314e-13, 
    8.0858813078427785e-13, 8.7647664515606285e-13, 9.4291530290297612e-13, 
    1.0058676196280073e-12, 1.0639223648037393e-12, 1.1163387924228788e-12, 
    1.1630926815389544e-12, 1.2047973752863682e-12, 1.2426224571703794e-12, 
    1.2780773201134572e-12, 1.312852603237771e-12, 1.3485398364256559e-12, 
    1.3864656606421008e-12, 1.4274509122222423e-12, 1.4716926340613059e-12, 
    1.5186469165368795e-12, 1.567045061008361e-12, 1.6149058064086586e-12, 
    1.6597290206968417e-12, 1.698645191821898e-12, 1.7287019017486105e-12, 
    1.7471062387305847e-12, 1.7515307789103489e-12, 1.7403249486785214e-12, 
    1.7127527497061535e-12, 1.6690690645971675e-12, 1.6105969073592793e-12, 
    1.5396510045239402e-12, 1.4594071041947123e-12, 1.3736726990900317e-12, 
    1.2866481857325042e-12, 1.2026019402972961e-12, 1.1256037963049787e-12, 
    1.0592311571318529e-12, 1.0063711732905504e-12, 9.69050508968595e-13, 
    9.4837196380571596e-13, 9.4450294668021174e-13, 9.567650759310711e-13, 
    9.837287717512235e-13, 1.023421348262696e-12, 1.0735188353402421e-12, 
    1.1315229638789003e-12, 1.194941118657419e-12, 1.2614624921161505e-12, 
    1.3290307497080558e-12, 1.395931764317694e-12, 1.4607839882880178e-12, 
    1.5225295839604418e-12, 1.5803610055661469e-12, 1.6336592506589129e-12, 
    1.6819071069547795e-12, 1.72463895185268e-12, 1.7613909655652403e-12, 
    1.79169879126914e-12, 1.815125281190018e-12, 1.8313321989300977e-12, 
    1.8401699525956477e-12, 1.8417633694809689e-12, 1.8366197865862035e-12, 
    1.8256975028010847e-12, 1.8104187090553791e-12, 1.7926814536701804e-12, 
    1.7747668017715071e-12, 1.7591963491997451e-12, 1.7485634415291876e-12, 
    1.7453195533483904e-12, 1.7515450720239975e-12, 1.7687424030941579e-12, 
    1.7976728950857551e-12, 1.8382367821316433e-12, 1.8894364109958848e-12, 
    1.9493984283950284e-12, 2.0154902302344014e-12, 2.0845037618846063e-12, 
    2.1528538606859346e-12, 2.216856986373923e-12, 2.2729698512922392e-12, 
    2.3180219009734475e-12, 2.3494172924188707e-12, 2.365268163929496e-12, 
    2.3644666522299109e-12, 2.3467198335056711e-12, 2.3124916589264074e-12, 
    2.2629166802688944e-12, 2.199657386511253e-12, 2.1247818094791138e-12, 
    2.040569453583908e-12, 1.9493989379985419e-12, 1.8535947205389139e-12, 
    1.7553190342114375e-12, 1.6564890938735565e-12, 1.5587335891569827e-12, 
    1.4633526607233258e-12, 1.3713359286592501e-12, 1.2833718748344327e-12, 
    1.1998942980425271e-12, 1.1211307356124034e-12, 1.0471529762412042e-12, 
    9.7795503687206527e-13, 9.1349572453910455e-13, 8.5374644123001924e-13, 
    7.9874981914210805e-13, 7.4862956082899284e-13, 7.0360768429534796e-13, 
    6.6398884954250917e-13, 6.3014534112135141e-13, 6.0246885684121533e-13, 
    5.8131907120367625e-13, 5.6696980936398972e-13, 5.59541168847199e-13, 
    5.5895431571948521e-13, 5.649009446173654e-13, 5.7683110884590037e-13, 
    5.9396619465200054e-13, 6.1532648779262126e-13, 6.3982278551523928e-13, 
    6.6633609992350441e-13, 6.9380544520845931e-13, 7.2135152512063571e-13, 
    7.4834556824043009e-13, 7.7448285919610743e-13, 7.9980929825908733e-13, 
    8.2470667664024657e-13, 8.4982908638593312e-13, 8.7599893744239896e-13, 
    9.0406487019523748e-13, 9.3475649136845911e-13, 9.6850451598321933e-13, 
    1.0053139388641827e-12, 1.0446593844240457e-12, 1.0854275985142406e-12, 
    1.1259340544772745e-12, 1.1639948809269092e-12, 1.1970435679249063e-12, 
    1.2223428460049316e-12, 1.2371495498303653e-12, 1.2389456450245862e-12, 
    1.2256310895164154e-12, 1.195676271277857e-12, 1.1482435543530481e-12, 
    1.0832459136610955e-12, 1.0013427624703197e-12, 9.0390332605576248e-13, 
    7.9291721756586705e-13, 6.7088468647262193e-13, 5.406929707220018e-13, 
    4.0548705099735115e-13, 2.6856003530958428e-13, 1.332314469145158e-13, 
    2.7570099446772153e-15, -1.1973486502970301e-13, -2.3136186407481648e-13, 
    -3.2951951805722323e-13, -4.1198027505081182e-13, 
    -4.7694574890103166e-13, -5.2311300781561541e-13, 
    -5.4974496087074669e-13, -5.5669226199770378e-13, 
    -5.4442002637314802e-13, -5.1400839330806445e-13, 
    -4.6711945240375426e-13, -4.0591126644449689e-13, 
    -3.3294639355577724e-13, -2.5107226228014424e-13, 
    -1.6327185830777632e-13, -7.252149340520573e-14, 1.8363732288275432e-14, 
    1.0686172772519543e-13, 1.908643907152167e-13, 2.6875264509165656e-13, 
    3.3947214494405363e-13, 4.0254022162578195e-13, 4.5802417068300667e-13, 
    5.065282876173006e-13, 5.491189933399639e-13, 5.8722023396010403e-13, 
    6.2251362658470288e-13, 6.5682932024262929e-13, 6.9201366088243194e-13, 
    7.2981520282579606e-13, 7.7175783465133022e-13, 8.1903836278452759e-13, 
    8.7245128375441483e-13, 9.3232901822566399e-13, 9.9849609722121376e-13, 
    1.0702930483187358e-12, 1.1466014007900906e-12, 1.2259175965983125e-12, 
    1.3064398376357036e-12, 1.3862043132950173e-12, 1.4632040435820631e-12, 
    1.5355348111454277e-12, 1.6015144124960889e-12, 1.6597987204754561e-12, 
    1.7094597925730219e-12, 1.7500286493064268e-12, 1.781489263373084e-12, 
    1.8042496748827109e-12, 1.819043201071157e-12, 1.8268212356586624e-12, 
    1.8286020382199004e-12, 1.8253147379824385e-12, 1.817649552397808e-12, 
    1.8059358383384531e-12, 1.7900602027586652e-12, 1.769418702418536e-12, 
    1.7429513741728003e-12, 1.7092303696429237e-12, 1.66660708602252e-12, 
    1.6134089279635721e-12, 1.5481646211758091e-12, 1.4698266192414954e-12, 
    1.3779883203091146e-12, 1.273048651560851e-12, 1.1563122757835945e-12, 
    1.0300152403194301e-12, 8.9726737862110609e-13, 7.6189834335267792e-13, 
    6.2825387273751056e-13, 5.0090950496283846e-13, 3.8438336808997944e-13, 
    2.8282393531464173e-13, 1.997179851172699e-13, 1.3767669603094608e-13, 
    9.8274815981680654e-14, 8.1929470912001693e-14, 8.7920561579284417e-14, 
    1.1446759411181484e-13, 1.5887511977151008e-13, 2.1774608387103745e-13, 
    2.872134098720325e-13, 3.6320730967368928e-13, 4.4169795274019462e-13, 
    5.1891712610915735e-13, 5.9154036122512144e-13, 6.5681276658926882e-13, 
    7.1260703311908157e-13, 7.574558428008041e-13, 7.9048862993798726e-13, 
    8.1138016505650701e-13, 8.2023771133467169e-13, 8.1750570942644399e-13, 
    8.0386439737826143e-13, 7.8016357805638291e-13, 7.473459669925588e-13, 
    7.0645083548244203e-13, 6.5862866248070396e-13, 6.0513734081756856e-13, 
    5.4737688706034175e-13, 4.8693826489092896e-13, 4.2559622141508603e-13, 
    3.652887975637396e-13, 3.0806389206790074e-13, 2.5600719127547217e-13, 
    2.1113134276910187e-13, 1.7524805341773999e-13, 1.4985364136708089e-13, 
    1.3601100199633575e-13, 1.3426783173552705e-13, 1.4461070852366054e-13, 
    1.6645338725113428e-13, 1.9868223472825989e-13, 2.3974453440087973e-13, 
    2.8774840418495107e-13, 3.4061311319114654e-13, 3.9622048537907249e-13, 
    4.5258140106328401e-13, 5.0794740584705186e-13, 5.6096783005882664e-13, 
    6.1074861627845371e-13, 6.5692883340194665e-13, 6.9968061691763849e-13, 
    7.3968937620853298e-13, 7.7806929133449552e-13, 8.1626971009788139e-13, 
    8.5591787230374707e-13, 8.9865169788291401e-13, 9.4593663166616412e-13, 
    9.9891533457877479e-13, 1.0581928063778921e-12, 1.1237341705288164e-12, 
    1.1947740936573359e-12, 1.269776742742326e-12, 1.3464622342672073e-12, 
    1.4218870328003671e-12, 1.4925885754220414e-12, 1.5547806388291328e-12, 
    1.6045692561010417e-12, 1.6381961728932926e-12, 1.6522888251684538e-12, 
    1.6440751636092216e-12, 1.6116035712063536e-12, 1.5538931490272521e-12, 
    1.4710558842902452e-12, 1.3643443459538827e-12, 1.2361814262402559e-12, 
    1.090074363913798e-12, 9.3054814549898682e-13, 7.6296508805191478e-13, 
    5.9332865529453752e-13, 4.2800972099291003e-13, 2.7351473673980584e-13, 
    1.361441184562915e-13, 2.1709067644894642e-14, -6.4788478890081987e-14, 
    -1.1940440560940836e-13, -1.3949411962161516e-13, 
    -1.2385190540381007e-13, -7.2815804685763257e-14, 1.175236688022789e-14, 
    1.265482600358375e-13, 2.6701461375295182e-13, 4.2758386974139908e-13, 
    6.0198401829082855e-13, 7.8357271235798748e-13, 9.656940179635968e-13, 
    1.1420079098436259e-12, 1.3067864712803145e-12, 1.4551430553947562e-12, 
    1.5832259452674586e-12, 1.6882967110088627e-12, 1.7687700929212438e-12, 
    1.8241664558824152e-12, 1.8550329157872736e-12, 1.8627890017716737e-12, 
    1.8496028559067042e-12, 1.8182109022075343e-12, 1.7717674573712615e-12, 
    1.713697371339216e-12, 1.6475828057887157e-12, 1.577035514721594e-12, 
    1.5056182121105399e-12, 1.4367458150619178e-12, 1.3736023073384025e-12, 
    1.3190361138338267e-12, 1.2754774669653783e-12, 1.2448136081271621e-12, 
    1.2282952286942514e-12, 1.2264091687463824e-12, 1.2388304113596579e-12, 
    1.2643472520769925e-12, 1.3008891511745321e-12, 1.3455457546348857e-12, 
    1.3947254181099763e-12, 1.4443227245595071e-12, 1.4899572247301001e-12, 
    1.5272265382356713e-12, 1.5520424453528621e-12, 1.5608650786947118e-12, 
    1.5509876644909174e-12, 1.5207075652506909e-12, 1.4694468406789138e-12, 
    1.3977745943109987e-12, 1.3073431700263514e-12, 1.200712657925943e-12, 
    1.0811850272477992e-12, 9.5250951538363711e-13, 8.1862335758107125e-13, 
    6.8337417249513831e-13, 5.5031842691098282e-13, 4.2250419522629037e-13, 
    3.0239439775464468e-13, 1.9178478707177339e-13, 9.1830622634930818e-14, 
    3.0826872748652638e-15, -7.4403054958768818e-14, -1.4098413428390207e-13, 
    -1.9728748098524156e-13, -2.4412620370185146e-13, 
    -2.8238064453840346e-13, -3.1293127089687764e-13, 
    -3.3656992140475641e-13, -3.5395157769834159e-13, -3.655423774590527e-13, 
    -3.7159719431339673e-13, -3.7212510992782646e-13, 
    -3.6689151933954217e-13, -3.5543648909994572e-13, 
    -3.3711899631033817e-13, -3.1117999008103872e-13, 
    -2.7684168020681152e-13, -2.3341580246280116e-13, 
    -1.8044332613450607e-13, -1.1779405821254034e-13, 
    -4.5822816876976509e-14, 3.4597531456366505e-14, 1.2203916554670113e-13, 
    2.1448087785746833e-13, 3.0941872821732755e-13, 4.0397359676689546e-13, 
    4.9505492760236687e-13, 5.7956885784436364e-13, 6.5462403913574542e-13, 
    7.1775136486192844e-13, 7.6708685581647508e-13, 8.0153903751612354e-13, 
    8.2086639825773898e-13, 8.2574049352249479e-13, 8.1769956993842791e-13, 
    7.9904950780833702e-13, 7.727077632200827e-13, 7.4199219355981884e-13, 
    7.1037027283498489e-13, 6.8121678403872418e-13, 6.5756111391541772e-13, 
    6.4187673471572159e-13, 6.35911216162548e-13, 6.4061151752244913e-13, 
    6.5608553998625181e-13, 6.8167940497345427e-13, 7.1609417202433974e-13, 
    7.575702671797596e-13, 8.0409830012491932e-13, 8.5363697556496098e-13, 
    9.0430470391574083e-13, 9.5454479357125813e-13, 1.0032134124414631e-12, 
    1.0496254052055526e-12, 1.0935016400352295e-12, 1.1348962144629357e-12, 
    1.1740726101777853e-12, 1.2113307439675411e-12, 1.2468746431827288e-12, 
    1.2806824558024262e-12, 1.3124273514157321e-12, 1.3414321648653679e-12, 
    1.3666919935684747e-12, 1.3869489623824774e-12, 1.4008022912606007e-12, 
    1.4068405221539462e-12, 1.403811987197288e-12, 1.3907426787329455e-12, 
    1.3670872491677202e-12, 1.3327916303122409e-12, 1.2883455035980231e-12, 
    1.2347676706141396e-12, 1.1735687933115679e-12, 1.1066332116786041e-12, 
    1.0361059675228711e-12, 9.6423324647729978e-13, 8.9322757904281034e-13, 
    8.2507924303088179e-13, 7.6144280344606234e-13, 7.0351455424274507e-13, 
    6.5196204644809024e-13, 6.0686530025520706e-13, 5.6774954800508959e-13, 
    5.3360837445592423e-13, 5.0302186830130731e-13, 4.7426956725540844e-13, 
    4.4551151876673405e-13, 4.1496157857454922e-13, 3.8107533018835181e-13, 
    3.4273523165000522e-13, 2.993849047656424e-13, 2.5113458421354472e-13, 
    1.9880151436519213e-13, 1.4388477928106755e-13, 8.8463244855751633e-14, 
    3.5047467819237819e-14, -1.3646844066863611e-14, -5.492153368078892e-14, 
    -8.6365932240388135e-14, -1.0605800186574626e-13, -1.1277200243503933e-13,
  // Sqw-Na(1, 0-1999)
    0.11872328912208698, 0.11819983744539017, 0.11664686818370407, 
    0.11411550385130845, 0.11068758830953912, 0.10647094766968056, 
    0.10159332370119023, 0.096195471925616893, 0.090423960419904886, 
    0.084424195065253116, 0.078334137276820925, 0.072279081477697599, 
    0.066367735871672148, 0.06068971712669298, 0.055314442453006901, 
    0.050291293763977771, 0.04565084684837141, 0.04140690808548185, 
    0.03755908227121272, 0.034095604107041051, 0.030996196846769016, 
    0.02823476721087434, 0.025781798518910035, 0.023606357379002071, 
    0.021677677927550806, 0.01996632795072923, 0.018444991380297426, 
    0.017088921294231028, 0.015876127499016124, 0.014787364637505492, 
    0.013805982562000614, 0.01291769251293869, 0.012110292348481468, 
    0.011373383246421911, 0.010698100108976726, 0.010076869094415276, 
    0.0095031986600669534, 0.0089715053151828168, 0.0084769718217362986, 
    0.0080154335867995731, 0.0075832881407558476, 0.0071774225645549654, 
    0.0067951542214380609, 0.0064341809218618007, 0.006092537522766628, 
    0.0057685568095720589, 0.0054608332561317981, 0.0051681888670935738, 
    0.0048896407682209146, 0.0046243705301103289, 0.0043716954062430957, 
    0.0041310417593102009, 0.0039019209637076104, 0.0036839080299766623, 
    0.0034766231196735483, 0.0032797160245671866, 0.0030928535862731351, 
    0.0029157099415010801, 0.0027479594002076117, 0.0025892717020757736, 
    0.0024393093515427669, 0.002297726702485466, 0.0021641704496526901, 
    0.0020382811841617283, 0.0019196956842028412, 0.0018080496388161429, 
    0.00170298054094489, 0.0016041305336693093, 0.0015111490471137517, 
    0.0014236951185297993, 0.0013414393395273776, 0.0012640654177449215, 
    0.0011912713719533707, 0.0011227703980511456, 0.0010582914491062744, 
    0.00099757956800351506, 0.00094039600023208695, 0.00088651810139012946, 
    0.00083573904325481081, 0.00078786731687924467, 0.00074272603265190503, 
    0.00070015202542600408, 0.00065999478602590713, 0.0006221152560018623, 
    0.0005863845373467486, 0.00055268258013456536, 0.00052089691647830532, 
    0.0004909215076125701, 0.0004626557621301581, 0.00043600376830961517, 
    0.00041087376373461127, 0.0003871778432580825, 0.00036483188428096462, 
    0.00034375564874824979, 0.00032387300634819288, 0.0003051122147433105, 
    0.00028740619114542011, 0.00027069271523473749, 0.00025491451552077415, 
    0.00024001920819333194, 0.00022595907716776761, 0.00021269070393534103, 
    0.0002001744735424403, 0.0001883739964561056, 0.00017725549377110768, 
    0.00016678719456434806, 0.00015693878947826791, 0.00014768097492365829, 
    0.00013898510934817995, 0.00013082298887506766, 0.00012316673631740461, 
    0.00011598878685345751, 0.00010926194667779901, 0.0001029594982093091, 
    9.7055326716269136e-05, 9.1524047699719852e-05, 8.6341120837864094e-05, 
    8.1482943367513653e-05, 7.6926922176000521e-05, 7.2651528613523281e-05, 
    6.8636342543224754e-05, 6.4862092336067181e-05, 6.1310695717914913e-05, 
    5.7965303244208876e-05, 5.4810342528058535e-05, 5.1831558012126068e-05, 
    4.9016038741473252e-05, 4.6352225724201909e-05, 4.382989121996369e-05, 
    4.1440084551752281e-05, 3.9175042415579631e-05, 3.7028065626290655e-05, 
    3.4993368162401568e-05, 3.3065907670245052e-05, 3.1241208775076553e-05, 
    2.9515191331842935e-05, 2.7884015050064526e-05, 2.634394989237801e-05, 
    2.4891278603729818e-05, 2.3522234142059385e-05, 2.2232971160282096e-05, 
    2.1019567515627099e-05, 1.9878049428210587e-05, 1.8804432598517055e-05, 
    1.7794771363146506e-05, 1.6845208701436631e-05, 1.5952021351090911e-05, 
    1.5111656134158924e-05, 1.4320755507322215e-05, 1.3576172056971376e-05, 
    1.2874972965100344e-05, 1.2214436288680302e-05, 1.1592041227925267e-05, 
    1.1005454492977797e-05, 1.0452514538716131e-05, 9.931214965972586e-06, 
    9.4396879059004207e-06, 8.976187806309077e-06, 8.5390757739711743e-06, 
    8.1268045111733188e-06, 7.7379038991174698e-06, 7.3709673926466069e-06, 
    7.0246395507412455e-06, 6.6976051923493276e-06, 6.3885807891478723e-06, 
    6.0963087543456603e-06, 5.8195552299335653e-06, 5.557111805823715e-06, 
    5.3078013234842183e-06, 5.0704875490558623e-06, 4.8440880835880094e-06, 
    4.6275894672575137e-06, 4.4200630899618462e-06, 4.2206803052460132e-06, 
    4.0287251025025386e-06, 3.843602851081993e-06, 3.6648439799609864e-06, 
    3.4921019623633218e-06, 3.3251455678185751e-06, 3.1638459428153756e-06, 
    3.0081595971963106e-06, 2.8581087345179457e-06, 2.7137605217684202e-06, 
    2.5752068363415505e-06, 2.4425457791193004e-06, 2.3158658601387842e-06, 
    2.1952333216169752e-06, 2.0806826450240226e-06, 1.9722099614200487e-06, 
    1.8697688950257604e-06, 1.7732683299535611e-06, 1.6825716829564022e-06, 
    1.597497443598392e-06, 1.5178209493779374e-06, 1.4432775336878265e-06, 
    1.3735672711668028e-06, 1.3083615180523871e-06, 1.2473113060612011e-06, 
    1.190057419930924e-06, 1.1362417181957607e-06, 1.0855189981924386e-06, 
    1.0375685146938474e-06, 9.9210417794709338e-07, 9.4888250533855567e-07, 
    9.0770757834843184e-07, 8.6843254170036666e-07, 8.3095753169292564e-07, 
    7.952242873298785e-07, 7.6120802786560437e-07, 7.289074327622731e-07, 
    6.9833370389900881e-07, 6.694997155534989e-07, 6.4241017044719277e-07, 
    6.1705350313748169e-07, 5.9339603549711635e-07, 5.7137863053138181e-07, 
    5.5091584310991033e-07, 5.3189735747198781e-07, 5.1419134826148928e-07, 
    4.9764931114249694e-07, 4.8211187599761136e-07, 4.6741512988949868e-07, 
    4.5339702165423953e-07, 4.399034807817457e-07, 4.2679394588920655e-07, 
    4.1394605607576758e-07, 4.012593086002047e-07, 3.8865753220176969e-07, 
    3.7609007173123081e-07, 3.6353163414024888e-07, 3.5098081048477073e-07, 
    3.3845736566501033e-07, 3.2599847076703152e-07, 3.1365413492983224e-07, 
    3.0148216206482314e-07, 2.8954300229465462e-07, 2.7789487821991884e-07, 
    2.665895389133673e-07, 2.5566892951770695e-07, 2.4516297021994347e-07, 
    2.3508852512250123e-07, 2.2544952549814746e-07, 2.1623810608488852e-07, 
    2.0743653191209016e-07, 1.9901964321755956e-07, 1.9095753265966532e-07, 
    1.832181884232452e-07, 1.7576988434669741e-07, 1.6858316249052017e-07, 
    1.6163232561752446e-07, 1.5489642474320493e-07, 1.4835978319517827e-07, 
    1.4201213648589521e-07, 1.3584848570562016e-07, 1.2986876051920588e-07, 
    1.24077371421177e-07, 1.1848270308111351e-07, 1.1309657025328309e-07, 
    1.0793362839329336e-07, 1.030107111064186e-07, 9.8346057085593044e-08, 
    9.3958394048540613e-08, 8.9865864243157671e-08, 8.6084804036420468e-08, 
    8.2628422781489908e-08, 7.9505459991247235e-08, 7.6718926690959447e-08, 
    7.4265053176509243e-08, 7.2132565858310091e-08, 7.030239972989845e-08, 
    6.8747919625941213e-08, 6.7435677448751268e-08, 6.6326677743049927e-08, 
    6.5378069148578199e-08, 6.4545129959954593e-08, 6.3783381162116695e-08, 
    6.3050643387863628e-08, 6.2308859875921559e-08, 6.1525533725043505e-08, 
    6.0674673102116437e-08, 5.9737194586687355e-08, 5.8700796841211295e-08, 
    5.7559373948340128e-08, 5.6312084061559729e-08, 5.4962216871883533e-08, 
    5.3516011473819465e-08, 5.1981562513519919e-08, 5.0367922358879634e-08, 
    4.8684463704939478e-08, 4.6940520346359682e-08, 4.5145278447032359e-08, 
    4.3307856232190293e-08, 4.1437488130095141e-08, 3.9543725437881294e-08, 
    3.7636575479893738e-08, 3.5726525363584628e-08, 3.382442631866013e-08, 
    3.194124766803644e-08, 3.0087737027831885e-08, 2.8274043543663904e-08, 
    2.6509368124981949e-08, 2.480170114312814e-08, 2.3157691985327933e-08, 
    2.1582672686436262e-08, 2.0080830533151331e-08, 1.865549972494234e-08, 
    1.7309521230024165e-08, 1.6045608420310958e-08, 1.4866653493661446e-08, 
    1.377591809170794e-08, 1.2777067236410301e-08, 1.1874028534607143e-08, 
    1.1070682647999695e-08, 1.037041517791184e-08, 9.7755791731952478e-09, 
    9.2869309502636169e-09, 8.9031066519098612e-09, 8.6202046575838139e-09, 
    8.4315283877247928e-09, 8.3275286373755245e-09, 8.2959644903904201e-09, 
    8.3222815030489948e-09, 8.390184883454795e-09, 8.4823682468626315e-09, 
    8.5813445799186106e-09, 8.670317934943027e-09, 8.7340312218927368e-09, 
    8.7595284199121785e-09, 8.7367769237719755e-09, 8.6591081478539483e-09, 
    8.5234487699634097e-09, 8.3303321100317511e-09, 8.0836950337329434e-09, 
    7.7904817699805703e-09, 7.4600881761690393e-09, 7.1036900372864878e-09, 
    6.7335039415989973e-09, 6.3620313354361794e-09, 6.001333511812699e-09, 
    5.6623803101767379e-09, 5.354506731383951e-09, 5.0850026599228261e-09, 
    4.8588499499777273e-09, 4.6786112986140641e-09, 4.5444652022649482e-09, 
    4.454373339507752e-09, 4.4043592597560647e-09, 4.3888726628423938e-09, 
    4.4012099586961439e-09, 4.4339609769465816e-09, 4.4794520823572245e-09, 
    4.5301589698992144e-09, 4.5790661499757773e-09, 4.6199559847887451e-09, 
    4.6476160762125766e-09, 4.6579607571748002e-09, 4.6480686917529936e-09, 
    4.6161447707539132e-09, 4.5614190387295308e-09, 4.4839992707439829e-09, 
    4.3846954324475192e-09, 4.2648349483959487e-09, 4.1260861254942509e-09, 
    3.970304895668849e-09, 3.7994158769040023e-09, 3.6153345087977747e-09, 
    3.4199318252017299e-09, 3.2150386574867254e-09, 3.0024813452046696e-09, 
    2.7841378394885126e-09, 2.5620004151894929e-09, 2.3382309861799597e-09, 
    2.1151956620386491e-09, 1.8954681443864828e-09, 1.6817952781175588e-09, 
    1.4770232716269514e-09, 1.2839879518208867e-09, 1.1053776662731112e-09, 
    9.4358114621136113e-10, 8.0053539569874993e-10, 6.7758938768319377e-10, 
    5.7539849176608426e-10, 4.9386178407128605e-10, 4.3211046125009867e-10, 
    3.8855054774159643e-10, 3.6095800551290246e-10, 3.4661911691213911e-10, 
    3.4250502497537856e-10, 3.4546613546582179e-10, 3.5243054663423912e-10, 
    3.6059058979695961e-10, 3.6756327319674356e-10, 3.7151295867220823e-10, 
    3.7122854931730765e-10, 3.6615164880137634e-10, 3.563566162956463e-10, 
    3.4248728415237487e-10, 3.2565852347761982e-10, 3.0733289446316623e-10, 
    2.8918369525182278e-10, 2.7295551296234172e-10, 2.6033228022479604e-10, 
    2.528207247166549e-10, 2.5165486386846683e-10, 2.5772451802403094e-10, 
    2.7152871539900629e-10, 2.9315286151719228e-10, 3.2226760729580106e-10, 
    3.581464014781902e-10, 3.9969899006880749e-10, 4.4551804373910265e-10, 
    4.939367700590657e-10, 5.4309546635002295e-10, 5.9101528536531768e-10, 
    6.3567717888362285e-10, 6.7510380297415348e-10, 7.0744150042376044e-10, 
    7.310390337516204e-10, 7.4451926868998722e-10, 7.4684019871679465e-10, 
    7.3734168161201257e-10, 7.1577524002755636e-10, 6.8231523679244171e-10, 
    6.3755101852833291e-10, 5.824609339420027e-10, 5.183705102432388e-10, 
    4.4689777666101619e-10, 3.6988962734479599e-10, 2.8935301137404559e-10, 
    2.0738483513328241e-10, 1.2610363916614995e-10, 4.7585709838576737e-11, 
    -2.6192683206053831e-11, -9.3405796083101957e-11, 
    -1.5242127549548909e-10, -2.0183504585133093e-10, -2.404984782240578e-10, 
    -2.6753775108931719e-10, -2.8236565578116575e-10, 
    -2.8468577557617966e-10, -2.7448934578648868e-10, 
    -2.5204496693752602e-10, -2.1788187512315469e-10, 
    -1.7276746555785011e-10, -1.1768035369558666e-10, 
    -5.3780146725166742e-11, 1.762458574105226e-11, 9.5108989972451067e-11, 
    1.771642031196574e-10, 2.6222862140553903e-10, 3.4871787079362105e-10, 
    4.3505365270024724e-10, 5.1969166079457423e-10, 6.0114908502144693e-10, 
    6.7803181655140919e-10, 7.4906147112926576e-10, 8.1310177964892085e-10, 
    8.6918374554305713e-10, 9.1652840474880868e-10, 9.5456611829716643e-10, 
    9.8295099949292206e-10, 1.0015694021198458e-09, 1.0105415354291546e-09, 
    1.0102156613185678e-09, 1.0011547822936779e-09, 9.8411608923082363e-10, 
    9.6002391095822774e-10, 9.2993724272145845e-10, 8.9501312325161766e-10, 
    8.5646743225087711e-10, 8.1553464803883067e-10, 7.734282055801499e-10, 
    7.3130292999698117e-10, 6.9022099060814234e-10, 6.5112250707070647e-10, 
    6.1480179792107007e-10, 5.8188993796478878e-10, 5.5284404229390649e-10, 
    5.2794337693882169e-10, 5.0729223636542263e-10, 4.9082907356634479e-10, 
    4.7834143719067598e-10, 4.6948575074195236e-10, 4.6381111162233838e-10, 
    4.6078588053483468e-10, 4.5982599476453921e-10, 4.6032368739720519e-10, 
    4.6167544377881871e-10, 4.6330799421177663e-10, 4.6470139286714262e-10, 
    4.6540813641971042e-10, 4.650678345171403e-10, 4.6341681328464404e-10, 
    4.6029253437984159e-10, 4.5563272902395073e-10, 4.4946955725282752e-10, 
    4.419191201152985e-10, 4.3316704383108562e-10, 4.2345085282908816e-10, 
    4.1304020194634069e-10, 4.0221605766879949e-10, 3.9125012071406174e-10, 
    3.8038580658232382e-10, 3.6982213258743331e-10, 3.5970161228593368e-10, 
    3.5010320343329549e-10, 3.4104077477249931e-10, 3.3246732277876949e-10, 
    3.2428444543434684e-10, 3.1635630019004758e-10, 3.085266068244645e-10, 
    3.0063713882591399e-10, 2.925458611767854e-10, 2.8414300578838332e-10, 
    2.7536358631026724e-10, 2.6619529848955783e-10, 2.5668118933006261e-10, 
    2.4691718148282569e-10, 2.3704489330525988e-10, 2.2724080368824846e-10, 
    2.1770291528055151e-10, 2.0863636828831387e-10, 2.002392610573543e-10, 
    1.926898625757223e-10, 1.8613604957640722e-10, 1.8068752064871305e-10, 
    1.7641099990966818e-10, 1.7332840162686175e-10, 1.7141752809988455e-10, 
    1.7061507994893665e-10, 1.7082125948307893e-10, 1.7190562041678734e-10, 
    1.7371351728295574e-10, 1.7607287276319695e-10, 1.7880077306410884e-10, 
    1.8170973944599048e-10, 1.8461337331675532e-10, 1.8733136005987236e-10, 
    1.8969370757064672e-10, 1.9154435064878904e-10, 1.9274406324696242e-10, 
    1.9317292598237463e-10, 1.9273233939055752e-10, 1.9134676710705296e-10, 
    1.8896514890876193e-10, 1.8556210174859044e-10, 1.8113865257897205e-10, 
    1.7572256301491169e-10, 1.6936794611412264e-10, 1.6215412119214245e-10, 
    1.541835079355749e-10, 1.4557863816646434e-10, 1.3647819184540022e-10, 
    1.2703234550987855e-10, 1.1739754348206237e-10, 1.0773108007058727e-10, 
    9.8185738854593502e-11, 8.8904880371555997e-11, 8.0018190429344996e-11, 
    7.1638391339191142e-11, 6.3858940612612348e-11, 5.6752875426501675e-11, 
    5.0372652346398149e-11, 4.475094903691729e-11, 3.9902134601081316e-11, 
    3.5824309471415742e-11, 3.2501605330569006e-11, 2.9906624336029057e-11, 
    2.8002751272909136e-11, 2.6746373012725203e-11, 2.6088823757413631e-11, 
    2.5978193686619347e-11, 2.636094803656395e-11, 2.718346047363771e-11, 
    2.8393487560932804e-11, 2.9941592420486876e-11, 3.1782422791526021e-11, 
    3.3875820993382835e-11, 3.6187503945410099e-11, 3.8689342183901895e-11, 
    4.1358916477646883e-11, 4.4178518519295808e-11, 4.7133466616641724e-11, 
    5.0210021185676592e-11, 5.3393031341836396e-11, 5.6663719970336667e-11, 
    5.9997847915312846e-11, 6.3364637752496746e-11, 6.6726551453558088e-11, 
    7.0040135080184709e-11, 7.3257751327065678e-11, 7.6330110993454987e-11, 
    7.9209198634167121e-11, 8.1851308594795386e-11, 8.4219689245188395e-11, 
    8.6286587268331104e-11, 8.8034315832707454e-11, 8.9455337679739556e-11, 
    9.0551269341867778e-11, 9.1331108936399566e-11, 9.1808820948361714e-11, 
    9.200077742172844e-11, 9.19232907683795e-11, 9.159074011906e-11, 
    9.1014441657463342e-11, 9.0202583469565923e-11, 8.9161111538438854e-11, 
    8.7895638636137761e-11, 8.6414029008811252e-11, 8.4729415594302108e-11, 
    8.2863167802901541e-11, 8.0847491934303852e-11, 7.8727146292250151e-11, 
    7.6560070104749558e-11, 7.4416603315698699e-11, 7.2377347906040781e-11, 
    7.0529613502441709e-11, 6.8962835431239215e-11, 6.776317573999549e-11, 
    6.7007889602211835e-11, 6.6759797449802764e-11, 6.7062489919235056e-11, 
    6.7936533564296677e-11, 6.9377142287911937e-11, 7.1353368126523618e-11, 
    7.3808997706034517e-11, 7.6664971796137071e-11, 7.9823234073372195e-11, 
    8.3171599511168416e-11, 8.6589423046236208e-11, 8.9953586627784292e-11, 
    9.3144525786364945e-11, 9.6051839064008776e-11, 9.8579293670877982e-11, 
    1.0064891236856277e-10, 1.0220398899861195e-10, 1.0321089240185178e-10, 
    1.0365968024111036e-10, 1.0356343265678429e-10, 1.0295650266627109e-10, 
    1.0189173150516899e-10, 1.004368695908597e-10, 9.8670414412580009e-11, 
    9.6677138169666775e-11, 9.454354915381146e-11, 9.2353604787407568e-11, 
    9.0184856329545089e-11, 8.8105298100636144e-11, 8.6170978239707022e-11, 
    8.4424551675779717e-11, 8.2894714215046556e-11, 8.1596545181555763e-11, 
    8.0532540235988798e-11, 7.9694359130204976e-11, 7.9064938017901846e-11, 
    7.8620892157509503e-11, 7.8334922204523767e-11, 7.8178103336484205e-11, 
    7.812183271125193e-11, 7.8139374581157351e-11, 7.8206821891488439e-11, 
    7.8303595440803635e-11, 7.8412343586016834e-11, 7.8518489665309707e-11, 
    7.8609424262715216e-11, 7.8673566874604481e-11, 7.8699458367364036e-11, 
    7.8675024975822413e-11, 7.8587139214489658e-11, 7.8421567401648098e-11, 
    7.8163353839022784e-11, 7.779758139509832e-11, 7.7310426243568103e-11, 
    7.6690414507250315e-11, 7.5929679140623811e-11, 7.5025127083223879e-11, 
    7.3979254493403951e-11, 7.2800649113585756e-11, 7.1503934669353965e-11, 
    7.0109286652352028e-11, 6.8641400750682396e-11, 6.7128162290614829e-11, 
    6.5598943603720629e-11, 6.4082852935244255e-11, 6.2606966035357484e-11, 
    6.1194776760103543e-11, 5.9864905435464808e-11, 5.8630263318657966e-11, 
    5.7497607086428538e-11, 5.6467583480836982e-11, 5.553515503771164e-11, 
    5.4690379973068609e-11, 5.3919398024344993e-11, 5.3205581888663466e-11, 
    5.2530680150357483e-11, 5.1875954696859377e-11, 5.1223150191281395e-11, 
    5.0555367996127689e-11, 4.9857729838143784e-11, 4.9117943941827221e-11, 
    4.832668231666284e-11, 4.7477879529157659e-11, 4.6568908256253979e-11, 
    4.5600674549385301e-11, 4.4577579958255447e-11, 4.3507404141457534e-11, 
    4.2401020345323405e-11, 4.1271987038816775e-11, 4.0135976949626614e-11, 
    3.9010099140849997e-11, 3.7912062481638025e-11, 3.6859333838443664e-11, 
    3.5868250110715882e-11, 3.4953228517937727e-11, 3.4126056289024054e-11, 
    3.3395385926064711e-11, 3.2766444957922075e-11, 3.2240960030603177e-11, 
    3.1817300753627407e-11, 3.1490845991941293e-11, 3.1254457924399095e-11, 
    3.1099105370443119e-11, 3.1014470252331284e-11, 3.0989574819808657e-11, 
    3.1013323940110189e-11, 3.1074967558674548e-11, 3.1164428175371701e-11, 
    3.1272547010190118e-11, 3.1391218719440066e-11, 3.1513468282139095e-11, 
    3.1633481649890434e-11, 3.1746625577571803e-11, 3.1849482385662676e-11, 
    3.1939891263274467e-11, 3.2016989638780945e-11, 3.2081287714508332e-11, 
    3.2134679095984109e-11, 3.2180425202102324e-11, 3.2223048224266721e-11, 
    3.2268132346622445e-11, 3.2322006612523107e-11, 3.2391343107495879e-11, 
    3.2482655208124938e-11, 3.2601764549891809e-11, 3.2753249572889606e-11, 
    3.2939970842345729e-11, 3.3162669848355979e-11, 3.3419749538306676e-11, 
    3.3707229988914781e-11, 3.4018942756150024e-11, 3.4346879236389689e-11, 
    3.4681775191500306e-11, 3.5013837994548204e-11, 3.5333557160027124e-11, 
    3.5632506269064227e-11, 3.5904115927518833e-11, 3.614425557818912e-11, 
    3.6351629124666839e-11, 3.6527887400085572e-11, 3.6677447585960596e-11, 
    3.680700107121101e-11, 3.6924784657889727e-11, 3.7039635499533052e-11, 
    3.7159948741779093e-11, 3.7292616214369212e-11, 3.7442116271259428e-11, 
    3.7609736176972677e-11, 3.7793167556732682e-11, 3.7986401296463864e-11, 
    3.818004108164773e-11, 3.8361894581541644e-11, 3.8517938340909525e-11, 
    3.8633429175083235e-11, 3.8694136869482442e-11, 3.8687564695278451e-11, 
    3.860402917713678e-11, 3.843749007520733e-11, 3.8186139001462934e-11, 
    3.7852571340453609e-11, 3.7443678645418645e-11, 3.6970185220750064e-11, 
    3.6445945489206175e-11, 3.5887001653390139e-11, 3.5310573719637368e-11, 
    3.4733963535894478e-11, 3.4173556829291656e-11, 3.3643863771352881e-11, 
    3.3156784760737029e-11, 3.2721005098484547e-11, 3.2341666643388997e-11, 
    3.2020181472622908e-11, 3.1754321013845627e-11, 3.1538468770363634e-11, 
    3.1364071770236381e-11, 3.1220197011730171e-11, 3.109427316340163e-11, 
    3.0972850357104153e-11, 3.0842467052448986e-11, 3.0690463931968216e-11, 
    3.0505813263407808e-11, 3.0279805901514799e-11, 3.0006646627803665e-11, 
    2.9683824939057603e-11, 2.9312322589814709e-11, 2.8896523914067458e-11, 
    2.8443932624895247e-11, 2.7964625803219931e-11, 2.7470554251056547e-11, 
    2.6974640842414877e-11, 2.6489876934232938e-11, 2.6028393758197112e-11, 
    2.5600620760392228e-11, 2.5214611227978527e-11, 2.4875589900835872e-11, 
    2.4585716745748111e-11, 2.4344135631674823e-11, 2.414724876038465e-11, 
    2.3989208757511404e-11, 2.3862534746247408e-11, 2.3758823561953446e-11, 
    2.3669472856498294e-11, 2.3586341763496727e-11, 2.350229026283378e-11, 
    2.341158515173701e-11, 2.3310109864267132e-11, 2.3195402406616534e-11, 
    2.3066546809510164e-11, 2.2923901184619736e-11, 2.276877946315741e-11, 
    2.2603069152096674e-11, 2.2428880928222986e-11, 2.2248261067758085e-11, 
    2.2062984795447961e-11, 2.1874490580419551e-11, 2.1683917793923437e-11, 
    2.1492265065195811e-11, 2.130062859521334e-11, 2.1110474109951362e-11, 
    2.0923919940949377e-11, 2.0743960393432473e-11, 2.0574604298169655e-11, 
    2.04208841460095e-11, 2.0288730407718451e-11, 2.0184706562329417e-11, 
    2.011558364527557e-11, 2.0087848325248874e-11, 2.010711985035062e-11, 
    2.0177574117962916e-11, 2.0301374174214327e-11, 2.0478225016820582e-11, 
    2.0705043410976862e-11, 2.0975807494341992e-11, 2.128160138926603e-11, 
    2.1610867479753146e-11, 2.1949843654897156e-11, 2.2283181352742878e-11, 
    2.2594684668351578e-11, 2.2868132562638693e-11, 2.3088116526907464e-11, 
    2.3240844219452795e-11, 2.3314853115939753e-11, 2.3301592100567237e-11, 
    2.3195821377894444e-11, 2.299583655286781e-11, 2.2703497680216062e-11, 
    2.2324100338354464e-11, 2.1866049517700898e-11, 2.1340470122080621e-11, 
    2.076066620572433e-11, 2.0141575186316451e-11, 1.9499150465652574e-11, 
    1.8849788438192834e-11, 1.8209732930356138e-11, 1.7594562881712744e-11, 
    1.7018686896569528e-11, 1.6494926062162503e-11, 1.6034166662395946e-11, 
    1.5645089855377449e-11, 1.5333966692521908e-11, 1.5104577469448553e-11, 
    1.4958168378447126e-11, 1.4893549104296004e-11, 1.4907198351869683e-11, 
    1.4993481731482237e-11, 1.5144877804757665e-11, 1.5352279249702609e-11, 
    1.5605242753559953e-11, 1.5892323327588855e-11, 1.6201345938072217e-11, 
    1.6519744179754576e-11, 1.6834825984982855e-11, 1.7134121928129422e-11, 
    1.7405687129826979e-11, 1.7638467872452647e-11, 1.7822617540030865e-11, 
    1.79498727478548e-11, 1.8013849041358055e-11, 1.8010371511059097e-11, 
    1.7937676594499854e-11, 1.7796590213348493e-11, 1.7590579244453264e-11, 
    1.7325702124964537e-11, 1.7010427324078096e-11, 1.6655343325742569e-11, 
    1.6272735900704175e-11, 1.5876088609679275e-11, 1.5479496541802549e-11, 
    1.5097051971486479e-11, 1.4742209009158593e-11, 1.4427189267637387e-11, 
    1.4162462541217351e-11, 1.3956311579623089e-11, 1.3814533355263158e-11, 
    1.3740283752138003e-11, 1.3734044716697895e-11, 1.3793765339686188e-11, 
    1.3915082861874341e-11, 1.4091676163922504e-11, 1.4315650532588352e-11, 
    1.4577980783805345e-11, 1.4868937154446159e-11, 1.5178491831216702e-11, 
    1.549668402609043e-11, 1.5813926142502598e-11, 1.6121234022552488e-11, 
    1.6410405464046122e-11, 1.6674143860944625e-11, 1.6906126688835491e-11, 
    1.710103641201448e-11, 1.725457608290302e-11, 1.7363452884784602e-11, 
    1.7425375714183816e-11, 1.7439043476706061e-11, 1.7404159363542874e-11, 
    1.7321415177343773e-11, 1.7192520972816598e-11, 1.702021015361424e-11, 
    1.6808246156379474e-11, 1.6561391225273516e-11, 1.6285356782231596e-11, 
    1.5986699247196524e-11, 1.5672692873954341e-11, 1.535109117627394e-11, 
    1.5029906750224106e-11, 1.4717108944393381e-11, 1.4420330431137636e-11, 
    1.4146533382729711e-11, 1.390175361561801e-11, 1.3690803386539077e-11, 
    1.3517118500694649e-11, 1.3382596887810119e-11, 1.3287593971728693e-11, 
    1.3230902156304058e-11, 1.320990511518149e-11, 1.3220700500826006e-11, 
    1.3258369644012977e-11, 1.3317195021892361e-11, 1.3390972319108033e-11, 
    1.3473275420728356e-11, 1.355777434996365e-11, 1.3638472629297149e-11, 
    1.3709998660575378e-11, 1.3767786825998033e-11, 1.380831448307957e-11, 
    1.3829216055273865e-11, 1.3829443148041578e-11, 1.3809292627760219e-11, 
    1.3770467669698626e-11, 1.3716014158503175e-11, 1.3650253485068027e-11, 
    1.3578578529189798e-11, 1.3507248138129008e-11, 1.3443029516035362e-11, 
    1.339280687919719e-11, 1.3363128992290584e-11, 1.3359715219316844e-11, 
    1.3386914160192207e-11, 1.3447232315063994e-11, 1.3540899028732126e-11, 
    1.36655625123202e-11, 1.3816094077154536e-11, 1.3984625586252587e-11, 
    1.4160717288797273e-11, 1.4331769775091226e-11, 1.4483607526933193e-11, 
    1.4601208581404656e-11, 1.4669542237853714e-11, 1.4674487541184439e-11, 
    1.4603699385142172e-11, 1.4447456641561119e-11, 1.4199355203387722e-11, 
    1.3856874451896415e-11, 1.3421673772465241e-11, 1.2899731671013918e-11, 
    1.230122299528527e-11, 1.1640175522416776e-11, 1.0933921603565716e-11, 
    1.0202393535365386e-11, 9.4672509604883854e-12, 8.7509638769903552e-12, 
    8.0757983626974105e-12, 7.4628525171030704e-12, 6.9310972944504831e-12, 
    6.4965650728314875e-12, 6.1716138385688438e-12, 5.9644134028009494e-12, 
    5.878578184364254e-12, 5.9130509087830262e-12, 6.0621902534316506e-12, 
    6.3160826682546517e-12, 6.661080104899046e-12, 7.0805159157566511e-12, 
    7.5555796870166638e-12, 8.0663087666672704e-12, 8.5926333200832532e-12, 
    9.1154206440041631e-12, 9.6174590975408954e-12, 1.0084303928807523e-11, 
    1.0504917486220222e-11, 1.0872082123472127e-11, 1.1182535405397407e-11, 
    1.1436795774717342e-11, 1.1638729472756561e-11, 1.1794851762950302e-11, 
    1.1913454539707285e-11, 1.200363404204068e-11, 1.2074280511532222e-11, 
    1.2133176384974881e-11, 1.2186250788493381e-11, 1.2237083417589909e-11, 
    1.2286691716460245e-11, 1.2333628763066455e-11, 1.2374354820439329e-11, 
    1.2403860392499896e-11, 1.2416419349986912e-11, 1.2406436409971362e-11, 
    1.2369208651515649e-11, 1.2301601670929259e-11, 1.220247933286239e-11, 
    1.2072910595823219e-11, 1.1916079713628598e-11, 1.1736979215054169e-11, 
    1.1541872661625075e-11, 1.1337671185059673e-11, 1.1131227921060958e-11, 
    1.0928720675068952e-11, 1.0735131646734452e-11, 1.0553926498298808e-11, 
    1.0386932248118284e-11, 1.0234421202606531e-11, 1.009539933147327e-11, 
    9.968027197729104e-12, 9.850062875098404e-12, 9.7393619511780362e-12, 
    9.6342762936521012e-12, 9.5339452160136926e-12, 9.4384296223042838e-12, 
    9.3486997505129871e-12, 9.2664641578020031e-12, 9.1939039770151946e-12, 
    9.1333239600582541e-12, 9.0868132373287013e-12, 9.0559099138222331e-12, 
    9.0413618940470797e-12, 9.0429740453877795e-12, 9.0595677589382551e-12, 
    9.0890309595702041e-12, 9.1284732907977345e-12, 9.1744200709497332e-12, 
    9.2230554174882229e-12, 9.2704633723287551e-12, 9.3128541590657487e-12, 
    9.3467822368758772e-12, 9.369290910669394e-12, 9.3780451284992155e-12, 
    9.3714225449956441e-12, 9.3485392749220314e-12, 9.3092719046351674e-12, 
    9.2542226868420542e-12, 9.1846456168370731e-12, 9.1023502789508586e-12, 
    9.0095455182119539e-12, 8.9086666750128649e-12, 8.8021755664709207e-12, 
    8.6923518093784914e-12, 8.5810819107572984e-12, 8.4697147935794413e-12, 
    8.3589321876262115e-12, 8.2486995963851718e-12, 8.1383041338381645e-12, 
    8.0264562318447733e-12, 7.9114798943987348e-12, 7.7915453610980012e-12, 
    7.6649176853129747e-12, 7.5302313895015528e-12, 7.3867151070071797e-12, 
    7.2343682241585434e-12, 7.0740754181505906e-12, 6.9076203980409704e-12, 
    6.7376448122669785e-12, 6.5675268384805909e-12, 6.4012130819956943e-12, 
    6.2430300309171052e-12, 6.0974775705233298e-12, 5.9690412667299804e-12, 
    5.862036248630658e-12, 5.7804581005004405e-12, 5.7278894102847847e-12, 
    5.70741478880355e-12, 5.7215750613853377e-12, 5.7722789545166335e-12, 
    5.8607717664586817e-12, 5.9875547627039592e-12, 6.1523213478710747e-12, 
    6.3538816543828408e-12, 6.5901260541004563e-12, 6.8579662979888097e-12, 
    7.1533505997349391e-12, 7.4713158930008482e-12, 7.8060949874582984e-12, 
    8.1512613667557406e-12, 8.4999313580739812e-12, 8.8449985189755397e-12, 
    9.1793856672755799e-12, 9.4962691201703543e-12, 9.7892890724685657e-12, 
    1.0052736509500439e-11, 1.0281647299378388e-11, 1.0471866393234067e-11, 
    1.0620045428739974e-11, 1.0723592312938304e-11, 1.0780613836812555e-11, 
    1.0789829112201091e-11, 1.0750513262960128e-11, 1.0662469219618859e-11, 
    1.0526037479073676e-11, 1.0342151014471755e-11, 1.0112452627518186e-11, 
    9.8393874310389204e-12, 9.5263346216158116e-12, 9.1777126974966175e-12, 
    8.7990088662204539e-12, 8.3967576547091898e-12, 7.9784216546572688e-12, 
    7.5521637503021319e-12, 7.1265294097918995e-12, 6.7100878935120268e-12, 
    6.310996399277156e-12, 5.9365780266952637e-12, 5.592922284128294e-12, 
    5.2845860049754683e-12, 5.0143810138517311e-12, 4.7833112155236053e-12, 
    4.5906434237231695e-12, 4.4341070745885321e-12, 4.3102011058339479e-12, 
    4.2145858145491272e-12, 4.1424767501589024e-12, 4.0890381105346906e-12, 
    4.0497062606068764e-12, 4.0204228021328839e-12, 3.9977764497024597e-12, 
    3.9790028060616748e-12, 3.9619334047432481e-12, 3.9448512902721618e-12, 
    3.9263408145503684e-12, 3.9051071993004028e-12, 3.8798649180493443e-12, 
    3.8492569534846986e-12, 3.8118505803210054e-12, 3.7661856389079406e-12, 
    3.7108793387606871e-12, 3.6447567382520151e-12, 3.5669896471574327e-12, 
    3.4772429895238169e-12, 3.3757654788009911e-12, 3.2634875332679166e-12, 
    3.1420563227151138e-12, 3.0138529171943778e-12, 2.8819929468332222e-12, 
    2.7502924917576479e-12, 2.6232253598954834e-12, 2.5058772794597171e-12, 
    2.4038554701477634e-12, 2.3231904720215906e-12, 2.2701630875312679e-12, 
    2.2511351979012983e-12, 2.2722706592694816e-12, 2.3392551275236011e-12, 
    2.45692776571688e-12, 2.6289540725910957e-12, 2.857442890155182e-12, 
    3.1426536590312918e-12, 3.4827424298236706e-12, 3.873617699143371e-12, 
    4.3089144741462424e-12, 4.7801096422688054e-12, 5.2767789700058739e-12, 
    5.7869683438235431e-12, 6.2976958706002099e-12, 6.7955181081836688e-12, 
    7.2671466319471009e-12, 7.7000545379667798e-12, 8.0830686361761465e-12, 
    8.4068378532701617e-12, 8.6642284895207837e-12, 8.8505520055978325e-12, 
    8.9636559347013538e-12, 9.0038428695752742e-12, 8.9736581573924882e-12, 
    8.8775358549121024e-12, 8.7213559192359971e-12, 8.5119455135332824e-12, 
    8.2565739745235905e-12, 7.9624481610725108e-12, 7.6363138304818548e-12, 
    7.2841342602625762e-12, 6.9109145637044665e-12, 6.5206581203301461e-12, 
    6.1164610550641554e-12, 5.7007275454306328e-12, 5.2754939365363964e-12, 
    4.8427599002392271e-12, 4.4048878137693928e-12, 3.964906234083159e-12, 
    3.5267890971220941e-12, 3.0955552219494789e-12, 2.6772992906271881e-12, 
    2.2790234337073083e-12, 1.9083863564126127e-12, 1.573290806257426e-12, 
    1.2814527684545046e-12, 1.0398830844733641e-12, 8.5441622734940857e-13, 
    7.2928067096609187e-13, 6.6679163889644482e-13, 6.6710019506329197e-13, 
    7.2817765638901571e-13, 8.4583461025686912e-13, 1.0139957882251415e-12, 
    1.2249684233860009e-12, 1.4699370099734945e-12, 1.7393792629110197e-12, 
    2.0236524487955745e-12, 2.3134238754118465e-12, 2.6002103054380231e-12, 
    2.8766901868935979e-12, 3.1370717482655887e-12, 3.3772125258291586e-12, 
    3.5947480819921342e-12, 3.7889876857625579e-12, 3.9608141031787185e-12, 
    4.1123668660443679e-12, 4.2467958377706775e-12, 4.3678191248004982e-12, 
    4.479418215262524e-12, 4.5854097243514155e-12, 4.689159633230338e-12, 
    4.7932952513433287e-12, 4.8995470079683285e-12, 5.0086132109447852e-12, 
    5.1201905623716042e-12, 5.2330211798634877e-12, 5.3450828745525192e-12, 
    5.453776924778888e-12, 5.5562231424588195e-12, 5.649509126931817e-12, 
    5.7310164965124696e-12, 5.7986385235487007e-12, 5.8510339680396865e-12, 
    5.8877509566512575e-12, 5.9093315445243195e-12, 5.9172731184197209e-12, 
    5.9139760712644006e-12, 5.9025256209344802e-12, 5.8864784278556364e-12, 
    5.8695526252421911e-12, 5.8553329439581156e-12, 5.8469268305287526e-12, 
    5.8467190653372023e-12, 5.8561120283466622e-12, 5.8754064958386033e-12, 
    5.9037135749721248e-12, 5.9390395369171748e-12, 5.9783751544091867e-12, 
    6.0179617609931085e-12, 6.0535476703169271e-12, 6.0807593684181324e-12, 
    6.095430471729478e-12, 6.0939727400979801e-12, 6.0736804771192261e-12, 
    6.0330003051096918e-12, 5.9716846291581987e-12, 5.8908991068565249e-12, 
    5.7931559886382506e-12, 5.6821993436600708e-12, 5.5627343300082843e-12, 
    5.440110977485755e-12, 5.3198907170544381e-12, 5.2074415731337581e-12, 
    5.1074514295445307e-12, 5.0235536448696768e-12, 4.957989074659695e-12, 
    4.9114026149060509e-12, 4.8827453859120456e-12, 4.8693651087368039e-12, 
    4.8672030052849226e-12, 4.8711689928736326e-12, 4.8755727571604546e-12, 
    4.8746509139859437e-12, 4.8630847981568884e-12, 4.8365027217242931e-12, 
    4.7918594913719515e-12, 4.7277158613345667e-12, 4.644351968976472e-12, 
    4.5437135046108698e-12, 4.4291933021436336e-12, 4.3052841756807826e-12, 
    4.1771371294428586e-12, 4.0500695323919805e-12, 3.9290847104965968e-12, 
    3.8184528684296e-12, 3.7214007139495846e-12, 3.6399296319832078e-12, 
    3.5747998193055138e-12, 3.5256538197156554e-12, 3.4912466390846492e-12, 
    3.4697809121821764e-12, 3.4592722148770684e-12, 3.4579088927442648e-12, 
    3.4643324947020248e-12, 3.4778557825805847e-12, 3.4985360863069825e-12, 
    3.5271409461356355e-12, 3.5650102096027321e-12, 3.6137772626315399e-12, 
    3.6751130721472401e-12, 3.7504012839562647e-12, 3.840440183725027e-12, 
    3.9452177619444892e-12, 4.0637384227299608e-12, 4.1939647518196236e-12, 
    4.3328281867787591e-12, 4.4763563715064379e-12, 4.6198234786267047e-12, 
    4.7579914813590928e-12, 4.8853567642145958e-12, 4.9964189607046045e-12, 
    5.0859265108345194e-12, 5.1491113930071238e-12, 5.1818927961276976e-12, 
    5.1810420875671683e-12, 5.1443185134049049e-12, 5.0705440905338096e-12, 
    4.9596652931750787e-12, 4.8127605579051774e-12, 4.6319890286652952e-12, 
    4.4205280157766579e-12, 4.1824414551240593e-12, 3.9225351688534802e-12, 
    3.6461547993448286e-12, 3.358975582642338e-12, 3.0667790575234494e-12, 
    2.7752134397972444e-12, 2.489590808073331e-12, 2.2147083732915568e-12, 
    1.9546903913016137e-12, 1.7129049502692965e-12, 1.4919179847126294e-12, 
    1.2935013754294136e-12, 1.1186962755539638e-12, 9.6789618472612713e-13, 
    8.409657068411254e-13, 7.3737227008091847e-13, 6.563083656019463e-13, 
    5.9681436529999764e-13, 5.5788688557435189e-13, 5.3855579448345442e-13, 
    5.3798257909582435e-13, 5.555059775744253e-13, 5.9068958972030165e-13, 
    6.4336810936703206e-13, 7.1365869193463326e-13, 8.0196820585649815e-13, 
    9.0896830938345795e-13, 1.0355462199804263e-12, 1.1827086752537984e-12, 
    1.3514702682231696e-12, 1.5426903726265441e-12, 1.7569219607353581e-12, 
    1.9942165036933553e-12, 2.2539834027585072e-12, 2.5348460307279272e-12, 
    2.8345780538711018e-12, 3.1500704313708182e-12, 3.4774038107796209e-12, 
    3.8119302817617496e-12, 4.1484698649669231e-12, 4.481498886364378e-12, 
    4.8053933009460958e-12, 5.1146386569938053e-12, 5.4040456668268575e-12, 
    5.6689089790832948e-12, 5.9051462584669981e-12, 6.1093490216197881e-12, 
    6.278836464779158e-12, 6.4116235914045915e-12, 6.5064168009884879e-12, 
    6.5625653489350095e-12, 6.5800447520857341e-12, 6.5594249103537821e-12, 
    6.5019007398946935e-12, 6.4092920967640028e-12, 6.2840875946163668e-12, 
    6.1294693475000499e-12, 5.9493400313110995e-12, 5.7482813558904826e-12, 
    5.5315025126285485e-12, 5.3047153016132818e-12, 5.07397084408102e-12, 
    4.8454198877250724e-12, 4.6250962006603341e-12, 4.4186094327521997e-12, 
    4.2308920356038665e-12, 4.065996820971126e-12, 3.9269086254677225e-12, 
    3.8154391413952634e-12, 3.7321945966879453e-12, 3.6766545959312479e-12, 
    3.6472846755955333e-12, 3.6417167543297942e-12, 3.65697934902698e-12, 
    3.6897262214962125e-12, 3.7364462368462944e-12, 3.7936881673620076e-12, 
    3.8582028232615611e-12, 3.9270582914375024e-12, 3.9976982415717065e-12, 
    4.0679804384029335e-12, 4.136162115589928e-12, 4.2008638498104837e-12, 
    4.2610232278232726e-12, 4.3158522460993282e-12, 4.364771334039192e-12, 
    4.4073660947286734e-12, 4.4433228092038457e-12, 4.4723879419913404e-12, 
    4.494314852493284e-12, 4.5088186576092819e-12, 4.5155364848715285e-12, 
    4.5140081483093012e-12, 4.5036548691040186e-12, 4.4838117798852676e-12, 
    4.4537717916503663e-12, 4.4128397815755457e-12, 4.36043787357475e-12, 
    4.2961970390411123e-12, 4.2200701642437508e-12, 4.1324119098540856e-12, 
    4.0340374054852824e-12, 3.9262345593820244e-12, 3.8107486842493488e-12, 
    3.6896769127027299e-12, 3.5653593276839847e-12, 3.4402150162872036e-12, 
    3.3165861850579281e-12, 3.1965661393929279e-12, 3.0818698737289821e-12, 
    2.973752698855375e-12, 2.8729883321968244e-12, 2.7799074672347008e-12, 
    2.6944924445844812e-12, 2.6165267179684584e-12, 2.5457720912403588e-12, 
    2.4821150198447332e-12, 2.4257156404770018e-12, 2.3770757321546601e-12, 
    2.3370452329372557e-12, 2.3067204783562764e-12, 2.2872765840709777e-12, 
    2.2797166370071033e-12, 2.2845899777559922e-12, 2.3016974382905176e-12, 
    2.3298491201593073e-12, 2.366679952091864e-12, 2.4085967670888501e-12, 
    2.4508510235977867e-12, 2.487755061078826e-12, 2.5130078933376886e-12, 
    2.5201517584635833e-12, 2.5030498098914131e-12, 2.4564040447255465e-12, 
    2.3762009876157387e-12, 2.2601062918890587e-12, 2.1076825165607968e-12, 
    1.9204998715284172e-12, 1.7020818248091642e-12, 1.4577156124647859e-12, 
    1.1941014853047654e-12, 9.1896242242611498e-13, 6.4056917214882182e-13, 
    3.6726740871206737e-13, 1.0700982615419456e-13, -1.3302953050851942e-13, 
    -3.4681235111837081e-13, -5.2964767486581523e-13, 
    -6.7836897793417491e-13, -7.9136814671407392e-13, 
    -8.6858988767059658e-13, -9.1139286693862052e-13, 
    -9.2241154697345013e-13, -9.0531288405394765e-13, 
    -8.6454749966652611e-13, -8.0504580867260693e-13, 
    -7.3194740152456479e-13, -6.5027720081127569e-13, 
    -5.6468356074063148e-13, -4.7917456694253108e-13, 
    -3.9690791807028264e-13, -3.2002016621277527e-13, 
    -2.4955053032118253e-13, -1.8540285550179707e-13, 
    -1.2640066426903557e-13, -7.0409004618080625e-14, 
    -1.4522614704604938e-14, 4.4672874910760937e-14, 1.1084648533869221e-13, 
    1.8760676951064e-13, 2.7821754615896375e-13, 3.8533119158111195e-13, 
    5.1079777612662003e-13, 6.5549487463196436e-13, 8.1929964085746971e-13, 
    1.0010710425406324e-12, 1.1987804884984271e-12, 1.4096470902500578e-12, 
    1.6303731826497187e-12, 1.8573458789339054e-12, 2.0869113240469643e-12, 
    2.3155558397274761e-12, 2.5400875649445567e-12, 2.7577319468594773e-12, 
    2.9661773769608029e-12, 3.1635367061556162e-12, 3.3482708891432116e-12, 
    3.5190328859913618e-12, 3.6745530713401904e-12, 3.8134739611146665e-12, 
    3.9342463107685878e-12, 4.0350691770263114e-12, 4.1138869764255034e-12, 
    4.1684575936230902e-12, 4.1965041525323606e-12, 4.1959056359632821e-12, 
    4.1649315697913311e-12, 4.1024904824970777e-12, 4.0083805652072671e-12, 
    3.8834748515198658e-12, 3.7298822654307647e-12, 3.5509986404595219e-12, 
    3.3514841135500599e-12, 3.1371415278138614e-12, 2.9146888419489187e-12, 
    2.6914745770859163e-12, 2.4751122716391967e-12, 2.273092641440618e-12, 
    2.0923840627692436e-12, 1.9390491481990531e-12, 1.8179299358120686e-12, 
    1.7323880176571378e-12, 1.6841600648411703e-12, 1.6733121621346419e-12, 
    1.6983038023358637e-12, 1.7561378629995133e-12, 1.8426458278623111e-12, 
    1.9528106566587026e-12, 2.0811092126670498e-12, 2.2219059845713294e-12, 
    2.3698178261028095e-12, 2.5200143101704255e-12, 2.6684751487803339e-12, 
    2.8121332363771337e-12, 2.9489424242771047e-12, 3.0778328156609039e-12, 
    3.1985887389239257e-12, 3.3116446222544891e-12, 3.4178588154814678e-12, 
    3.5182340221242795e-12, 3.6136976315621588e-12, 3.7048732739548714e-12, 
    3.7919860272494813e-12, 3.874794941257238e-12, 3.9526419765541519e-12, 
    4.02456163231668e-12, 4.0894874126523853e-12, 4.1464246799954801e-12, 
    4.1947069065324887e-12, 4.234154999691005e-12, 4.2651855396094432e-12, 
    4.2888432064663374e-12, 4.306750056907125e-12, 4.3209212260360078e-12, 
    4.3335682013728753e-12, 4.3468098605250962e-12, 4.3624044091475143e-12, 
    4.3814903012587616e-12, 4.4043999997746984e-12, 4.430549879311138e-12, 
    4.4584588381072105e-12, 4.4858308166113935e-12, 4.5097834685036363e-12, 
    4.527110518213998e-12, 4.534597772629037e-12, 4.5293552293735726e-12, 
    4.5090976346885978e-12, 4.4723824181265683e-12, 4.4187601690658396e-12, 
    4.3488190084804663e-12, 4.2641212198987005e-12, 4.1670500821964602e-12, 
    4.0605988494891853e-12, 3.9480650100626862e-12, 3.8327755253241845e-12, 
    3.7178053247476227e-12, 3.6057085080947211e-12, 3.4983602116349785e-12, 
    3.3968455900700391e-12, 3.3014471800740844e-12, 3.2117179788547037e-12, 
    3.1266154717318398e-12, 3.0446978692353574e-12, 2.964329571620877e-12, 
    2.8839141917983136e-12, 2.8020855879586992e-12, 2.7178581026492321e-12, 
    2.6307230074891087e-12, 2.5406909718505319e-12, 2.4482624204911484e-12, 
    2.3543500384513768e-12, 2.2601461629403105e-12, 2.1670122992710436e-12, 
    2.0763023883181932e-12, 1.9892489430774119e-12, 1.9068582023254781e-12, 
    1.829833074473791e-12, 1.7585374608089472e-12, 1.6930384407380497e-12, 
    1.6331358827324798e-12, 1.5784680351477242e-12, 1.5285961620097921e-12, 
    1.483150998286501e-12, 1.4419258915761434e-12, 1.404984140658419e-12, 
    1.3727240715116963e-12, 1.3459077837517066e-12, 1.325626910563439e-12, 
    1.3132606536779287e-12, 1.3103288421396735e-12, 1.3183483679169298e-12, 
    1.3386356083506893e-12, 1.3721060721586369e-12, 1.4190802192621859e-12, 
    1.4791204509187157e-12, 1.5508958784578593e-12, 1.6321545776162106e-12, 
    1.7197262133444266e-12, 1.8096250357755786e-12, 1.8972352458363518e-12, 
    1.9775329093179457e-12, 2.0453868103523396e-12, 2.0958452019667482e-12, 
    2.1244401441608459e-12, 2.1274466101502188e-12, 2.1020942195244937e-12, 
    2.0467037979835913e-12, 1.9607602108053472e-12, 1.8448780941259403e-12, 
    1.7007426750379326e-12, 1.5309517406780467e-12, 1.3388669576396093e-12, 
    1.1284158914995594e-12, 9.0392308064513701e-13, 6.6994735739145086e-13, 
    4.3115530269576856e-13, 1.9220211053028817e-13, -4.233481981284868e-14, 
    -2.6805411064757148e-13, -4.8076894394335011e-13, 
    -6.7660497301862163e-13, -8.5206613608103509e-13, 
    -1.0041374039427597e-12, -1.1303748631284088e-12, 
    -1.2289990239609448e-12, -1.2989655785390984e-12, 
    -1.3400111221620991e-12, -1.3526664549478595e-12, 
    -1.3381964682128541e-12, -1.2985150452097346e-12, 
    -1.2360681838439303e-12, -1.1536516690075052e-12, 
    -1.0542479962718797e-12, -9.4083463893907595e-13, 
    -8.1621365702046977e-13, -6.8287293079975765e-13, 
    -5.4287600868658219e-13, -3.9778880979546295e-13, 
    -2.4866041310868397e-13, -9.6056609694603634e-14, 5.990595665125388e-14, 
    2.1947394007353514e-13, 3.8311523474344102e-13, 5.5140429533538546e-13, 
    7.2488037000162014e-13, 9.0390268085949285e-13, 1.0885113620556828e-12, 
    1.2783159543333497e-12, 1.4723835573952585e-12, 1.6692130914265281e-12, 
    1.8666904322645698e-12, 2.0621382769436428e-12, 2.2523869840180217e-12, 
    2.4339124031723865e-12, 2.6029978834318887e-12, 2.7559468746760287e-12, 
    2.88929653702659e-12, 3.0000545095339077e-12, 3.0858977658049334e-12, 
    3.1453705594218496e-12, 3.1779915050605193e-12, 3.1843446831261723e-12, 
    3.1660625766455424e-12, 3.1257442484987896e-12, 3.0668092074308509e-12, 
    2.9932618861369675e-12, 2.9094196921140177e-12, 2.8195957432728097e-12, 
    2.7277764993543273e-12, 2.6372907295223458e-12, 2.5505675844113451e-12, 
    2.4689174375913805e-12, 2.3924329050377725e-12, 2.3199818812465996e-12, 
    2.2493295273558837e-12, 2.1773707134209396e-12, 2.1004603429605479e-12, 
    2.014823315089768e-12, 1.9170068114394186e-12, 1.804325880885163e-12, 
    1.6752766547834928e-12, 1.5298343904949706e-12, 1.3696613426882406e-12, 
    1.1981236923221078e-12, 1.0201658389417224e-12, 8.4201001216226754e-13, 
    6.707307203893377e-13, 5.13706636229544e-13, 3.7804809788070577e-13, 
    2.6998491148954409e-13, 1.943782659977722e-13, 1.5430955683420865e-13, 
    1.5079864465154535e-13, 1.8274891682619919e-13, 2.470523758065742e-13, 
    3.3886177125442576e-13, 4.5200681142560733e-13, 5.7949664729414145e-13, 
    7.1407142125768195e-13, 8.4872969533161536e-13, 9.7718700674883402e-13, 
    1.0942373635491117e-12, 1.1959601422652332e-12, 1.2797904032834027e-12, 
    1.3444513004791122e-12, 1.3897525947253179e-12, 1.4163259683982628e-12, 
    1.4253057815222613e-12, 1.4180137828973925e-12, 1.3957057138584839e-12, 
    1.3593754939838563e-12, 1.3096667975233649e-12, 1.2468965303069576e-12, 
    1.1711891456432711e-12, 1.082636491692784e-12, 9.815530251412194e-13, 
    8.6872384975838759e-13, 7.4563190987323315e-13, 6.1459872957225285e-13, 
    4.7886930774749838e-13, 3.4258940262277158e-13, 2.1068200101255137e-13, 
    8.8611058636466698e-14, -1.7891738728329913e-14, -1.031922053972182e-13, 
    -1.6210655419201827e-13, -1.9026010219962413e-13, -1.843903323676918e-13, 
    -1.4260001738796965e-13, -6.4496142482860829e-14, 4.8740580770070843e-14, 
    1.9441549485002535e-13, 3.6845742096427915e-13, 5.6567812479438311e-13, 
    7.80038347901151e-13, 1.0050219590259757e-12, 1.2339833341542799e-12, 
    1.4605062442818279e-12, 1.6787161720832337e-12, 1.8835466377426035e-12, 
    2.0709217834577493e-12, 2.2378701552619848e-12, 2.3825468958539103e-12, 
    2.5041833862379307e-12, 2.6029542802249598e-12, 2.6798295920680997e-12, 
    2.7363220170564478e-12, 2.7742685584529341e-12, 2.7955906765093176e-12, 
    2.802061338137414e-12, 2.7950990535504053e-12, 2.7756050327258088e-12, 
    2.7438484255851549e-12, 2.699415816946924e-12, 2.6412266032695934e-12, 
    2.5676264157324324e-12, 2.4765485423325478e-12, 2.365753857262476e-12, 
    2.2331303914580916e-12, 2.0770367743501329e-12, 1.8966598249820521e-12, 
    1.6923684204659323e-12, 1.4660116858649964e-12, 1.2211406463891876e-12, 
    9.6311552979466768e-13, 6.9907176877144044e-13, 4.3772238460786572e-13, 
    1.8899760880706787e-13, -3.6424337497942155e-14, -2.2772674370342517e-13, 
    -3.7462525406289092e-13, -4.6803808978987646e-13, 
    -5.0071535686753855e-13, -4.6775639443386385e-13, 
    -3.6698987089824572e-13, -1.9915713733777629e-13, 3.210673392898812e-14, 
    3.2047311185454171e-13, 6.573192408238775e-13, 1.0322467025793288e-12, 
    1.4336788965972435e-12, 1.8495162455362243e-12, 2.2677483185914293e-12, 
    2.6770147103778003e-12, 3.0670513775889048e-12, 3.4290207137955291e-12, 
    3.7557224206888771e-12, 4.0416648157803963e-12, 4.2830579550887074e-12, 
    4.4777201297658973e-12, 4.624940408454994e-12, 4.7253229017019435e-12, 
    4.7806587524454327e-12, 4.7937885902085572e-12, 4.7685080730283091e-12, 
    4.7094829464277692e-12, 4.6221827469483982e-12, 4.5127813523335238e-12, 
    4.3880420493480011e-12, 4.2551462679128074e-12, 4.1214486574274312e-12, 
    3.9941797875383429e-12, 3.8800845726269666e-12, 3.7850266216582248e-12, 
    3.7135754065271031e-12, 3.668616641107389e-12, 3.6510583274832166e-12, 
    3.6596113208800439e-12, 3.6907244810721766e-12, 3.7386730688762507e-12, 
    3.7958271633700732e-12, 3.8530876938596691e-12, 3.9004220923911707e-12, 
    3.927534781557269e-12, 3.9245775127888177e-12, 3.8828245109420081e-12, 
    3.7953061577145236e-12, 3.6573020542874606e-12, 3.4666695459205851e-12, 
    3.2239956109713362e-12, 2.9325258701365511e-12, 2.5979086878617674e-12, 
    2.2278184889820177e-12, 1.8314110932588585e-12, 1.4187406985410465e-12, 
    1.0001452680846445e-12, 5.856967102390221e-13, 1.8468625330059494e-13, 
    -1.9474892556728791e-13, -5.4590193731834715e-13, 
    -8.6363979252723351e-13, -1.1444493873244766e-12, 
    -1.3863690688998249e-12, -1.5888779124239808e-12, 
    -1.7526944841681654e-12, -1.8795908758903345e-12, 
    -1.9721371270354949e-12, -2.0334977995788759e-12, 
    -2.0671546367903655e-12, -2.0767060519514783e-12, 
    -2.0656097503616427e-12, -2.0369918053502907e-12, 
    -1.9934361055210786e-12, -1.9368564257747341e-12, 
    -1.8683823400974646e-12, -1.7883649646852647e-12, 
    -1.6964088001751752e-12, -1.5915466670297215e-12, 
    -1.4724453212270242e-12, -1.3377370809453726e-12, 
    -1.1863026024486469e-12, -1.0176748868421637e-12, 
    -8.3228113114727411e-13, -6.3169329015423769e-13, 
    -4.1875234819359935e-13, -1.9755301196117089e-13, 2.6735535657641906e-14, 
    2.4813714272384318e-13, 4.603042750672459e-13, 6.5697576233831726e-13, 
    8.3250622773884186e-13, 9.8233188216970124e-13, 1.103384980254664e-12, 
    1.1943439004754408e-12, 1.2557832895592482e-12, 1.290087828151336e-12, 
    1.3012489210110818e-12, 1.2944678889972208e-12, 1.2757021382087138e-12, 
    1.2511203384475891e-12, 1.226589875274474e-12, 1.2072094753863559e-12, 
    1.196961790038881e-12, 1.1985036158816426e-12, 1.2131289345117863e-12, 
    1.2408738905258727e-12, 1.2807690838811802e-12, 1.3311778123857143e-12, 
    1.3901798477714092e-12, 1.4559549221545953e-12, 1.5270908654440659e-12, 
    1.6028091788270747e-12, 1.6830514680979416e-12, 1.7684395610279633e-12, 
    1.8601045738265429e-12, 1.959401227690845e-12, 2.0675814556717694e-12, 
    2.1854377731591446e-12, 2.3129479246531255e-12, 2.4490233237432674e-12, 
    2.5913475117767679e-12, 2.7363525561323758e-12, 2.879318501185779e-12, 
    3.0146195543469126e-12, 3.1360786970902082e-12, 3.2374063648989619e-12, 
    3.3126705691448737e-12, 3.3567761214843798e-12, 3.3658752113142776e-12, 
    3.3377015785889455e-12, 3.2717798669715921e-12, 3.1694864083070065e-12, 
    3.0339766805783534e-12, 2.8699557351069418e-12, 2.6833458244208062e-12, 
    2.4808518583109927e-12, 2.2694885891348205e-12, 2.0560930012932732e-12, 
    1.8468685443034331e-12, 1.6469903895164669e-12, 1.4603227562860029e-12, 
    1.2892369211055948e-12, 1.1345580751279109e-12, 9.9563512107788657e-13, 
    8.705385956924258e-13, 7.563393688147463e-13, 6.4946986328370959e-13, 
    5.4612760847811756e-13, 4.4269262342221403e-13, 3.3611196733274102e-13, 
    2.2425206458795619e-13, 1.0615033124868801e-13, -1.7841400326105026e-14, 
    -1.4601787897310015e-13, -2.7541585713681616e-13, 
    -4.0202917297531978e-13, -5.2113627829825285e-13, 
    -6.2767910781990731e-13, -7.1671728966147045e-13, 
    -7.8384925313407517e-13, -8.2561066003284661e-13, -8.3978998980509679e-13,
  // Sqw-Na(2, 0-1999)
    0.08425175866251558, 0.084017297477583963, 0.083320128631458781, 
    0.082178571386948826, 0.080622100538810831, 0.078689847237389726, 
    0.076428664366906873, 0.073890900140289206, 0.071132038272865461, 
    0.068208362819812948, 0.065174791551205619, 0.062082996149978753, 
    0.058979894168902536, 0.05590656069220018, 0.052897571068445115, 
    0.049980753406712153, 0.047177303338821523, 0.044502195338572602, 
    0.041964815052484554, 0.039569735083011683, 0.03731756121191869, 
    0.035205785472758697, 0.033229594949644128, 0.031382598962696136, 
    0.029657450931856708, 0.028046353583417966, 0.026541446557334154, 
    0.025135083526835814, 0.023820011591040954, 0.022589469101896163, 
    0.021437219536428007, 0.020357538895274328, 0.019345172790905887, 
    0.018395277259870051, 0.017503354729973851, 0.016665193782134977, 
    0.015876818599188134, 0.015134451466910144, 0.014434489510374626, 
    0.013773495087872799, 0.013148197958418421, 0.012555506483725909, 
    0.011992524687788043, 0.011456571920660307, 0.010945202087230028, 
    0.010456219829758273, 0.0099876916188213465, 0.0095379503418466117, 
    0.0091055926235316925, 0.0086894687228895734, 0.0082886653953040002, 
    0.0079024825641444488, 0.0075304050034338188, 0.0071720704852408779, 
    0.0068272359912525706, 0.0064957436283768792, 0.0061774878267546636, 
    0.0058723852420950115, 0.0055803485443222511, 0.0053012649684021137, 
    0.0050349801541018395, 0.0047812874373811317, 0.0045399224074850223, 
    0.0043105622398260553, 0.0040928290794980436, 0.0038862965993632847, 
    0.0036904987950280594, 0.0035049401006310306, 0.0033291059987764866, 
    0.0031624734335523094, 0.0030045204936752687, 0.0028547349917249451, 
    0.0027126217086828057, 0.0025777081910884863, 0.002449549078547554, 
    0.0023277290051176842, 0.002211864165435127, 0.0021016026720073332, 
    0.0019966238589233134, 0.0018966367115256539, 0.0018013776206494015, 
    0.0017106076712108127, 0.0016241096750720266, 0.0015416851451131878, 
    0.0014631513813074789, 0.0013883388027844841, 0.0013170886168579815, 
    0.0012492508722744004, 0.0011846829047129285, 0.0011232481516744303, 
    0.0010648152931085244, 0.0010092576631254308, 0.00095645287497327742, 
    0.00090628260342798857, 0.00085863247327054083, 0.00081339200789839257, 
    0.00077045459775462212, 0.00072971745458864186, 0.00069108152551043483, 
    0.00065445135114417462, 0.00061973486495597765, 0.00058684314500845661, 
    0.00055569014295221133, 0.00052619242540242095, 0.00049826896743545332, 
    0.00047184103505166255, 0.00044683218272329947, 0.00042316837485615954, 
    0.00040077821891533163, 0.00037959327689288054, 0.00035954840477340556, 
    0.00034058206016011363, 0.00032263651842235372, 0.00030565794802006727, 
    0.00028959631458091252, 0.00027440510780408144, 0.00026004091128695509, 
    0.00024646285863671286, 0.00023363203600011229, 0.00022151089888036699, 
    0.00021006276884227829, 0.00019925146413511154, 0.00018904109951569336, 
    0.00017939606775327859, 0.00017028119195666586, 0.00016166201731375413, 
    0.00015350519570385076, 0.00014577890855223646, 0.00013845327270145479, 
    0.00013150068035619074, 0.000124896035826645, 0.00011861686681744247, 
    0.00011264330414661864, 0.00010695793892625047, 0.00010154557866131859, 
    9.6392932253923738e-05, 9.1488257979468099e-05, 8.6821008190759839e-05, 
    8.2381500383254196e-05, 7.816063729305425e-05, 7.414969009171634e-05, 
    7.0340149741500999e-05, 6.6723643325421354e-05, 6.3291905584463633e-05, 
    6.003679156610395e-05, 5.6950314444232264e-05, 5.4024693079661591e-05, 
    5.1252396331714067e-05, 4.8626174871086353e-05, 4.6139075561679025e-05, 
    4.3784437667465664e-05, 4.1555873619438487e-05, 3.9447239450954348e-05, 
    3.7452601111070757e-05, 3.5566202740083942e-05, 3.3782441871509898e-05, 
    3.2095854752672677e-05, 3.05011129469361e-05, 2.8993030460897143e-05, 
    2.7566579122809647e-05, 2.6216909002132413e-05, 2.4939370363257047e-05, 
    2.3729533933045867e-05, 2.2583206993997382e-05, 2.1496443800806118e-05, 
    2.0465549859592968e-05, 1.948708052360165e-05, 1.8557835018322782e-05, 
    1.767484733929296e-05, 1.6835375465799708e-05, 1.6036890054252177e-05, 
    1.5277063315340268e-05, 1.4553758256385319e-05, 1.3865018007001037e-05, 
    1.3209054637806845e-05, 1.2584236792140919e-05, 1.1989075589221466e-05, 
    1.1422208591143048e-05, 1.0882382075648828e-05, 1.0368432323591182e-05, 
    9.8792670050283587e-06, 9.4138479464607017e-06, 8.9711765275376887e-06, 
    8.5502826874457677e-06, 8.1502180588513439e-06, 7.7700531788224247e-06, 
    7.4088781554768473e-06, 7.0658057088615766e-06, 6.7399752399102194e-06, 
    6.4305565646853838e-06, 6.1367521805043666e-06, 5.8577973613112619e-06, 
    5.5929579228767521e-06, 5.3415260513248517e-06, 5.1028150423730924e-06, 
    4.8761540732605962e-06, 4.6608841749783799e-06, 4.4563563895766891e-06, 
    4.2619327243081179e-06, 4.0769900269287133e-06, 3.9009263937900527e-06, 
    3.7331692767265514e-06, 3.573184147963609e-06, 3.4204824615389903e-06, 
    3.2746277227265009e-06, 3.1352387243935666e-06, 3.0019893794215623e-06, 
    2.8746050112083164e-06, 2.7528553907322931e-06, 2.6365451745508847e-06, 
    2.5255026592729989e-06, 2.4195679070759444e-06, 2.3185813104159316e-06, 
    2.222373570470319e-06, 2.130757886865953e-06, 2.0435249280216322e-06, 
    1.9604408982920064e-06, 1.8812487655609176e-06, 1.8056724749213934e-06, 
    1.7334237635780827e-06, 1.664211012777601e-06, 1.5977494312361102e-06, 
    1.5337717637208792e-06, 1.4720386663896054e-06, 1.4123478917567327e-06, 
    1.3545414892874579e-06, 1.2985103533694253e-06, 1.2441956382799903e-06, 
    1.1915867984948135e-06, 1.1407162865745485e-06, 1.0916512245770613e-06, 
    1.0444826323953603e-06, 9.9931301816626146e-07, 9.5624328868659512e-07, 
    9.153600032202126e-07, 8.7672396577619909e-07, 8.4036103071763947e-07, 
    8.0625579891631429e-07, 7.7434862690546704e-07, 7.4453608710173614e-07, 
    7.1667473028315526e-07, 6.9058773975981904e-07, 6.6607385118344052e-07, 
    6.4291776011379693e-07, 6.2090115939967433e-07, 5.9981354380430105e-07, 
    5.7946198513075137e-07, 5.596792091979772e-07, 5.403294817823112e-07, 
    5.2131201821452831e-07, 5.0256185064493338e-07, 4.8404829994149885e-07, 
    4.6577138491635334e-07, 4.4775664612300564e-07, 4.3004895020192643e-07, 
    4.1270586983230219e-07, 3.9579120182385467e-07, 3.793691015567644e-07, 
    3.6349918676728655e-07, 3.4823281819773168e-07, 3.3361061589904383e-07, 
    3.1966113909330089e-07, 3.0640055717292305e-07, 2.9383308076320229e-07, 
    2.8195190476683018e-07, 2.7074043765681026e-07, 2.6017364060398283e-07, 
    2.5021936488485858e-07, 2.4083964087514761e-07, 2.3199192557367924e-07, 
    2.2363034803144606e-07, 2.1570700137980848e-07, 2.0817331540555397e-07, 
    2.0098151273797989e-07, 1.940861109533033e-07, 1.8744539381918295e-07, 
    1.8102274461457862e-07, 1.7478772125459082e-07, 1.6871675905700793e-07, 
    1.6279341354293288e-07, 1.5700809838000482e-07, 1.5135732749147056e-07, 
    1.4584252670880759e-07, 1.4046853242043757e-07, 1.3524193330333024e-07, 
    1.3016943268309749e-07, 1.252564074932511e-07, 1.2050581749581063e-07, 
    1.159175749011061e-07, 1.1148842774739789e-07, 1.0721234525791261e-07, 
    1.0308133037409243e-07, 9.9086530448342369e-08, 9.5219481061469378e-08, 
    9.1473303008894046e-08, 8.7843683360284475e-08, 8.4329504157723135e-08, 
    8.0933034405083334e-08, 7.7659663056131832e-08, 7.4517215383010105e-08, 
    7.1514951183424333e-08, 6.8662384594156157e-08, 6.5968084169260568e-08, 
    6.3438608047034109e-08, 6.1077701946609399e-08, 5.8885844296933764e-08, 
    5.6860168412001975e-08, 5.4994736779433735e-08, 5.3281094237282002e-08, 
    5.1708993434785126e-08, 5.0267170576762075e-08, 4.8944054589386478e-08, 
    4.7728315260777172e-08, 4.6609192087263464e-08, 4.5576587688242787e-08, 
    4.4620951943024558e-08, 4.3733017322461314e-08, 4.2903468569427568e-08, 
    4.2122636804125682e-08, 4.1380300227879656e-08, 4.0665651784040847e-08, 
    3.9967464164906084e-08, 3.9274447710343586e-08, 3.8575764638954121e-08, 
    3.7861636744771329e-08, 3.7123968375353153e-08, 3.6356902563061619e-08, 
    3.5557236621521411e-08, 3.4724641619335737e-08, 3.3861655506353055e-08, 
    3.2973447185183651e-08, 3.2067376101949745e-08, 3.1152393469705388e-08, 
    3.0238346755881753e-08, 2.9335254900851101e-08, 2.8452620236873999e-08, 
    2.7598833387394457e-08, 2.6780713181914686e-08, 2.6003205912013236e-08, 
    2.5269250705784611e-08, 2.4579801516578986e-08, 2.3933983814984052e-08, 
    2.3329355380180694e-08, 2.2762236847208337e-08, 2.2228077563981294e-08, 
    2.172182582917663e-08, 2.123827786834206e-08, 2.0772386758270611e-08, 
    2.0319518918870405e-08, 1.9875652046362028e-08, 1.943751288703319e-08, 
    1.9002656885945652e-08, 1.8569493524453245e-08, 1.8137262337552999e-08, 
    1.7705964653914387e-08, 1.727625640268042e-08, 1.6849307360316837e-08, 
    1.6426633407959815e-08, 1.6009909512208691e-08, 1.560077358086255e-08, 
    1.5200633318379734e-08, 1.4810490457063074e-08, 1.4430797607114501e-08, 
    1.4061362900232879e-08, 1.3701315082383803e-08, 1.3349137831207528e-08, 
    1.3002775923905729e-08, 1.2659808833421274e-08, 1.2317679571175691e-08, 
    1.1973959753389935e-08, 1.1626626097930846e-08, 1.1274320659308657e-08, 
    1.0916566738362892e-08, 1.0553915572737255e-08, 1.0188004525174057e-08, 
    9.8215161777548583e-09, 9.4580369777431634e-09, 9.1018246485215012e-09, 
    8.7575026018295564e-09, 8.4297074822736265e-09, 8.1227208044408396e-09, 
    7.8401177915876416e-09, 7.5844649756743995e-09, 7.3570939045215738e-09, 
    7.1579709952521365e-09, 6.9856750060815314e-09, 6.8374834096305021e-09, 
    6.7095595851085549e-09, 6.5972237320814585e-09, 6.4952837868483038e-09, 
    6.3983979090490911e-09, 6.3014388224225418e-09, 6.1998310653323857e-09, 
    6.0898361960968351e-09, 5.9687665636482456e-09, 5.8351154835034016e-09, 
    5.6885991954825824e-09, 5.5301136163282702e-09, 5.3616152251499501e-09, 
    5.1859405782555626e-09, 5.0065820407014631e-09, 4.8274387323231884e-09, 
    4.6525609619698157e-09, 4.4859047333379461e-09, 4.3311096311674974e-09, 
    4.1913102078191114e-09, 4.0689872961036956e-09, 3.9658626431770171e-09, 
    3.8828375487336438e-09, 3.819974378729674e-09, 3.7765181476129378e-09, 
    3.7509546641579526e-09, 3.7411006035207611e-09, 3.7442203782012823e-09, 
    3.7571637469834628e-09, 3.776517512238103e-09, 3.7987639265832727e-09, 
    3.8204382120421445e-09, 3.8382775162433921e-09, 3.8493545417992908e-09, 
    3.8511899314683677e-09, 3.8418393401544859e-09, 3.8199528020267285e-09, 
    3.7848059182212253e-09, 3.736303871476386e-09, 3.6749605830950435e-09, 
    3.6018557504532744e-09, 3.5185730555800007e-09, 3.4271223419733408e-09, 
    3.3298488060706426e-09, 3.2293317447989317e-09, 3.1282759947081185e-09, 
    3.0293993283996103e-09, 2.9353200604190696e-09, 2.8484496471382288e-09, 
    2.7708958601512878e-09, 2.7043819773268598e-09, 2.650187245408087e-09, 
    2.6091123760119374e-09, 2.5814722497882183e-09, 2.5671155798584738e-09, 
    2.5654690014909876e-09, 2.5756006823429682e-09, 2.596297048575514e-09, 
    2.6261451332425167e-09, 2.663613201725961e-09, 2.7071230626597819e-09, 
    2.7551093157326425e-09, 2.8060627212458037e-09, 2.8585574181738753e-09, 
    2.91126363998424e-09, 2.9629494497912252e-09, 3.0124758127124936e-09, 
    3.0587897724829728e-09, 3.1009197493184441e-09, 3.1379760845027641e-09, 
    3.1691582649658675e-09, 3.1937689239977697e-09, 3.2112329563791441e-09, 
    3.2211193972552352e-09, 3.2231627119163353e-09, 3.2172804712180244e-09, 
    3.2035845026906845e-09, 3.1823836362511753e-09, 3.1541769409823841e-09, 
    3.1196375806316469e-09, 3.0795881229659516e-09, 3.0349690216827593e-09, 
    2.9868022546687934e-09, 2.9361524714931347e-09, 2.8840877122880201e-09, 
    2.8316418762761305e-09, 2.7797804676454324e-09, 2.7293711112555822e-09, 
    2.6811597326386219e-09, 2.6357531518417117e-09, 2.5936082857342872e-09, 
    2.5550280975539908e-09, 2.5201638104519942e-09, 2.4890230067059225e-09, 
    2.4614825912483568e-09, 2.4373058058410354e-09, 2.4161620876344835e-09, 
    2.3976487496742388e-09, 2.3813133236384005e-09, 2.3666757705415381e-09, 
    2.3532496117122788e-09, 2.3405614690572562e-09, 2.3281684706030852e-09, 
    2.3156732077039064e-09, 2.3027358640100637e-09, 2.2890834476425117e-09, 
    2.2745157563170456e-09, 2.2589080715452667e-09, 2.2422103360088756e-09, 
    2.2244429069403856e-09, 2.2056888621549221e-09, 2.1860832592516017e-09, 
    2.1657996773334765e-09, 2.1450348570904556e-09, 2.1239921898724474e-09, 
    2.1028652387175149e-09, 2.0818223064637825e-09, 2.0609933375703178e-09, 
    2.040460033455079e-09, 2.0202501518062158e-09, 2.000336387619868e-09, 
    1.980639979887643e-09, 1.9610387208305032e-09, 1.9413786433811706e-09, 
    1.9214882594851734e-09, 1.9011941272089281e-09, 1.8803362058694397e-09, 
    1.8587817647021407e-09, 1.8364365767106323e-09, 1.8132526409444687e-09, 
    1.7892319045000946e-09, 1.7644260253310867e-09, 1.7389324804871312e-09, 
    1.712887719116708e-09, 1.6864582279153692e-09, 1.6598305117449102e-09, 
    1.6332008663622237e-09, 1.6067658290508349e-09, 1.5807138231416879e-09, 
    1.555218415601484e-09, 1.5304332885852625e-09, 1.5064888660764509e-09, 
    1.4834903254110959e-09, 1.4615167697489073e-09, 1.4406212017941718e-09, 
    1.4208310562063439e-09, 1.402149074428751e-09, 1.3845544785595417e-09, 
    1.3680043696633957e-09, 1.3524354877453978e-09, 1.3377663173910837e-09, 
    1.3238997216999583e-09, 1.3107260770054443e-09, 1.2981269436407759e-09, 
    1.285979142705184e-09, 1.2741591615833853e-09, 1.2625476004201645e-09, 
    1.2510335093118774e-09, 1.2395182933256266e-09, 1.2279190451612609e-09, 
    1.2161710025328649e-09, 1.2042291083146388e-09, 1.1920685281380271e-09, 
    1.1796841815794853e-09, 1.1670893021120979e-09, 1.1543132436294397e-09, 
    1.1413986348583207e-09, 1.1283981719736909e-09, 1.1153712303401108e-09, 
    1.1023805488845683e-09, 1.0894891438446114e-09, 1.0767576502746074e-09, 
    1.0642420977206179e-09, 1.0519922862798702e-09, 1.0400505774171393e-09, 
    1.028451208782334e-09, 1.0172199066500061e-09, 1.0063738381100396e-09, 
    9.9592167125589344e-10, 9.8586385504784708e-10, 9.7619295531790365e-10, 
    9.6689416445207453e-10, 9.5794593200760297e-10, 9.4932087164022195e-10, 
    9.4098687023553036e-10, 9.3290857477609896e-10, 9.2504912324200272e-10, 
    9.1737219194397726e-10, 9.0984417552357102e-10, 9.0243644301068369e-10, 
    8.9512740192456886e-10, 8.8790429011484884e-10, 8.8076435336646546e-10, 
    8.7371539695209612e-10, 8.6677545649344978e-10, 8.5997167133176882e-10, 
    8.5333828191456801e-10, 8.4691403459034739e-10, 8.4073903735181839e-10, 
    8.3485152925979542e-10, 8.2928468501517177e-10, 8.2406389848686399e-10, 
    8.1920460843054254e-10, 8.1471101602230409e-10, 8.1057552282976834e-10, 
    8.0677905443046238e-10, 8.0329192075355978e-10, 8.000751977873993e-10, 
    7.9708223396985349e-10, 7.9426021901184224e-10, 7.9155152577090947e-10, 
    7.8889489932285595e-10, 7.8622633606236698e-10, 7.8347992928869898e-10, 
    7.8058868760614959e-10, 7.7748564197342307e-10, 7.7410528144168243e-10, 
    7.7038557869217733e-10, 7.6627049876679854e-10, 7.6171306111559609e-10, 
    7.5667865414822992e-10, 7.511484663038445e-10, 7.451226113477886e-10, 
    7.3862267351911954e-10, 7.3169325567828511e-10, 7.2440235035587753e-10, 
    7.1684022285343658e-10, 7.0911684196142309e-10, 7.0135781013233423e-10, 
    6.9369907024412601e-10, 6.8628058236561788e-10, 6.792394697249629e-10, 
    6.727029872265044e-10, 6.6678186831517558e-10, 6.6156442148982578e-10, 
    6.5711183633424163e-10, 6.5345494822068599e-10, 6.5059269571926253e-10, 
    6.4849228129912357e-10, 6.4709104743059908e-10, 6.4629983534100564e-10, 
    6.4600763038576665e-10, 6.4608711095923787e-10, 6.4640083760812576e-10, 
    6.4680762180176989e-10, 6.4716885100216612e-10, 6.4735434182148897e-10, 
    6.4724756086739586e-10, 6.4674996715515851e-10, 6.4578432654742275e-10, 
    6.4429686905661887e-10, 6.4225833101336844e-10, 6.3966374550517406e-10, 
    6.3653118118005334e-10, 6.328993977894303e-10, 6.2882464710175997e-10, 
    6.2437674405838086e-10, 6.1963469524090952e-10, 6.1468205324010453e-10, 
    6.0960236725104551e-10, 6.0447492084356197e-10, 5.9937107743958393e-10, 
    5.9435140126400286e-10, 5.8946376894800647e-10, 5.8474252570982361e-10, 
    5.8020872898962849e-10, 5.7587131597477627e-10, 5.7172913409423115e-10, 
    5.6777348152870658e-10, 5.6399096354780419e-10, 5.6036623187292422e-10, 
    5.5688444722678458e-10, 5.5353309327280737e-10, 5.5030307047851476e-10, 
    5.471888811082898e-10, 5.4418807587142285e-10, 5.4129993006573778e-10, 
    5.3852374509026852e-10, 5.3585685481034971e-10, 5.3329280420657922e-10, 
    5.3081983581206422e-10, 5.2842001502237305e-10, 5.2606906052066374e-10, 
    5.2373699820905137e-10, 5.2138953791730389e-10, 5.1899011323630109e-10, 
    5.1650227754793097e-10, 5.1389232491309908e-10, 5.1113177198503691e-10, 
    5.0819954568933676e-10, 5.0508358181245116e-10, 5.0178182103056286e-10, 
    4.9830240051767854e-10, 4.9466317908164302e-10, 4.9089056886712745e-10, 
    4.8701790309972068e-10, 4.8308337608664503e-10, 4.7912787449291225e-10, 
    4.7519273986099033e-10, 4.7131769962673296e-10, 4.6753899149165797e-10, 
    4.6388787738249816e-10, 4.6038941624735003e-10, 4.5706168659608948e-10, 
    4.5391526890603812e-10, 4.5095311024094761e-10, 4.4817058764979046e-10, 
    4.4555588132693937e-10, 4.4309050003236202e-10, 4.4075008366521847e-10, 
    4.3850530812347565e-10, 4.3632306392477595e-10, 4.3416773589484497e-10, 
    4.3200269337823808e-10, 4.2979183325570979e-10, 4.2750123793348535e-10, 
    4.2510074796961363e-10, 4.2256548676271818e-10, 4.1987711386418829e-10, 
    4.1702485045736948e-10, 4.1400605292467111e-10, 4.1082642083314344e-10, 
    4.0749970060487448e-10, 4.0404698968170007e-10, 4.004955850739943e-10, 
    3.9687757843197338e-10, 3.9322817198310634e-10, 3.8958395743758629e-10, 
    3.8598113921515548e-10, 3.824539369428108e-10, 3.7903317705843773e-10, 
    3.7574517175942646e-10, 3.7261089385932292e-10, 3.6964551362677181e-10, 
    3.6685819733609897e-10, 3.6425225219986016e-10, 3.6182543349012258e-10, 
    3.5957050911320151e-10, 3.5747590618506687e-10, 3.555265196744421e-10, 
    3.5370450908859375e-10, 3.5199020371002225e-10, 3.5036295975427687e-10, 
    3.4880206337326099e-10, 3.4728756138882424e-10, 3.4580109409602973e-10, 
    3.4432661144544718e-10, 3.4285103143046778e-10, 3.4136469959638244e-10, 
    3.3986173849862267e-10, 3.3834012092395357e-10, 3.3680157446105802e-10, 
    3.3525118179213383e-10, 3.3369681673726026e-10, 3.3214832688224904e-10, 
    3.3061662625374711e-10, 3.2911267291790682e-10, 3.2764651228735603e-10, 
    3.2622634532021312e-10, 3.2485784213576105e-10, 3.2354362226323393e-10, 
    3.2228306124896154e-10, 3.2107234370768225e-10, 3.1990485277727116e-10, 
    3.1877173054118812e-10, 3.176627020591433e-10, 3.1656698854833861e-10, 
    3.1547428896584053e-10, 3.1437569304025259e-10, 3.1326452353877594e-10, 
    3.1213693622061575e-10, 3.1099232498369575e-10, 3.0983338432881292e-10, 
    3.0866590827218189e-10, 3.0749823304478013e-10, 3.0634044831127675e-10, 
    3.0520335907625067e-10, 3.0409732809960823e-10, 3.0303106302221801e-10, 
    3.0201050691467848e-10, 3.0103784546766087e-10, 3.0011083693706742e-10, 
    2.9922246137191598e-10, 2.9836098518756872e-10, 2.9751038306174108e-10, 
    2.9665119956449951e-10, 2.957616777797682e-10, 2.9481915535947272e-10, 
    2.9380156886601631e-10, 2.9268897792803448e-10, 2.9146494032626514e-10, 
    2.9011770672583086e-10, 2.8864103815408202e-10, 2.8703468654196198e-10, 
    2.8530442855427701e-10, 2.8346169631895078e-10, 2.8152280111081944e-10, 
    2.7950786082112806e-10, 2.7743945941382151e-10, 2.7534119947956574e-10, 
    2.7323620528249999e-10, 2.7114573048549706e-10, 2.690879227097273e-10, 
    2.6707688788117833e-10, 2.6512204965304374e-10, 2.6322788566652551e-10, 
    2.6139404387837172e-10, 2.5961579744286485e-10, 2.5788479748962288e-10, 
    2.5619010484935968e-10, 2.5451934848943675e-10, 2.5285999217866661e-10, 
    2.5120056310382519e-10, 2.4953179819391816e-10, 2.4784757968325326e-10, 
    2.4614563124837715e-10, 2.4442788374434277e-10, 2.4270051207741468e-10, 
    2.4097359908501009e-10, 2.3926046982460879e-10, 2.3757672030079621e-10, 
    2.3593903213074424e-10, 2.3436381866288313e-10, 2.3286585114345587e-10, 
    2.3145697945377644e-10, 2.3014500889978997e-10, 2.28932887858208e-10, 
    2.2781826562498959e-10, 2.2679342055049923e-10, 2.2584564835285446e-10, 
    2.2495799882132783e-10, 2.2411036082367116e-10, 2.2328074141421422e-10, 
    2.2244668579235267e-10, 2.2158667683081114e-10, 2.2068143895124103e-10, 
    2.1971500912544075e-10, 2.1867557058792832e-10, 2.1755594387035041e-10, 
    2.1635378560714394e-10, 2.1507148005378312e-10, 2.1371577539233813e-10, 
    2.1229723559341988e-10, 2.1082952855762483e-10, 2.0932866652395875e-10, 
    2.0781221089139692e-10, 2.0629846494543541e-10, 2.0480577358216196e-10, 
    2.0335183134832855e-10, 2.0195311575610244e-10, 2.0062437433706256e-10, 
    1.9937823000148015e-10, 1.982248687784459e-10, 1.9717182007817391e-10, 
    1.9622384900125859e-10, 1.9538294146851046e-10, 1.9464839153820235e-10, 
    1.940169691085879e-10, 1.9348316462932992e-10, 1.9303947347417763e-10, 
    1.9267670360245238e-10, 1.9238428117788229e-10, 1.9215049629323949e-10, 
    1.9196271828903878e-10, 1.9180754167497111e-10, 1.9167087739874291e-10, 
    1.9153800513705728e-10, 1.9139364719956424e-10, 1.9122205697625896e-10, 
    1.9100721385389437e-10, 1.9073311243096181e-10, 1.9038420892587403e-10, 
    1.8994597594033999e-10, 1.894055870087581e-10, 1.8875265911105818e-10, 
    1.8798000488640833e-10, 1.8708429751759662e-10, 1.8606660848343355e-10, 
    1.8493271648517099e-10, 1.8369317018454875e-10, 1.8236302046962654e-10, 
    1.8096130925649417e-10, 1.7951023988817924e-10, 1.7803417416679962e-10, 
    1.7655844639858034e-10, 1.7510814555830296e-10, 1.7370688456500432e-10, 
    1.723757143491974e-10, 1.7113214437752857e-10, 1.6998944376695749e-10, 
    1.689561643520206e-10, 1.6803594939072742e-10, 1.6722758156528936e-10, 
    1.6652530695799952e-10, 1.6591932452103164e-10, 1.6539648019355592e-10, 
    1.6494103119633833e-10, 1.645355044504908e-10, 1.6416153965306033e-10, 
    1.638007354760073e-10, 1.6343537764464431e-10, 1.6304911502210269e-10, 
    1.6262748921329871e-10, 1.6215835895025116e-10, 1.6163216469058179e-10, 
    1.6104209354455025e-10, 1.6038410596802391e-10, 1.5965687611011953e-10, 
    1.5886162146006876e-10, 1.5800188552581599e-10, 1.5708323626451142e-10, 
    1.5611296759217535e-10, 1.5509973769756468e-10, 1.5405324378646029e-10, 
    1.5298388119800244e-10, 1.5190243556165274e-10, 1.5081977733550794e-10, 
    1.4974661474520238e-10, 1.486932386199279e-10, 1.4766932055050611e-10, 
    1.4668369783438599e-10, 1.4574420763164883e-10, 1.4485749351958089e-10, 
    1.4402886092786057e-10, 1.4326212353700402e-10, 1.4255948611192157e-10, 
    1.4192146208809708e-10, 1.4134684511725737e-10, 1.4083272391073557e-10, 
    1.4037458787115053e-10, 1.3996649098545843e-10, 1.3960130473921892e-10, 
    1.3927102297916201e-10, 1.389671323793795e-10, 1.3868099099666875e-10, 
    1.3840423135233004e-10, 1.3812911641571187e-10, 1.3784886388307139e-10, 
    1.3755785837855914e-10, 1.3725178933099959e-10, 1.3692767183171355e-10, 
    1.3658375997592192e-10, 1.3621935470155491e-10, 1.358345663685673e-10, 
    1.3542999279794444e-10, 1.3500642671402621e-10, 1.345645688501205e-10, 
    1.341048162665789e-10, 1.3362709983457751e-10, 1.3313085053223631e-10, 
    1.3261502532156845e-10, 1.3207825230786052e-10, 1.315190019989629e-10, 
    1.3093582874227397e-10, 1.3032759499105129e-10, 1.2969373374750363e-10, 
    1.290343958500092e-10, 1.2835062825251014e-10, 1.2764444250971873e-10, 
    1.2691885738767491e-10, 1.261778491058194e-10, 1.2542629431111624e-10, 
    1.2466981782444351e-10, 1.2391464793481782e-10, 1.2316739374203691e-10, 
    1.2243485507648084e-10, 1.2172372101616824e-10, 1.2104034328337339e-10, 
    1.2039043779598626e-10, 1.1977884383353402e-10, 1.1920925730722592e-10, 
    1.1868404717774745e-10, 1.1820409122541197e-10, 1.1776873982509061e-10, 
    1.1737579703383614e-10, 1.1702167975870334e-10, 1.1670160062931148e-10, 
    1.1640990236779959e-10, 1.1614040650371945e-10, 1.1588686824163395e-10, 
    1.1564337513831956e-10, 1.1540479466579904e-10, 1.151670805067174e-10, 
    1.1492754454141724e-10, 1.1468493366480372e-10, 1.1443940956412152e-10, 
    1.1419230694407903e-10, 1.1394578518095182e-10, 1.1370233024984727e-10, 
    1.134642098759874e-10, 1.132328326213413e-10, 1.1300822889986176e-10, 
    1.1278855239970331e-10, 1.1256980819844759e-10, 1.1234571130970218e-10, 
    1.1210783329429863e-10, 1.118459091283717e-10, 1.1154840306107725e-10, 
    1.112031972955167e-10, 1.1079842566782769e-10, 1.1032328394411774e-10, 
    1.0976888852370272e-10, 1.091289528028812e-10, 1.0840038160069505e-10, 
    1.0758362200405811e-10, 1.0668284398171954e-10, 1.057058468966907e-10, 
    1.0466381258833113e-10, 1.0357084015216408e-10, 1.0244337109469868e-10, 
    1.0129947457125307e-10, 1.0015812485485001e-10, 9.9038431873764446e-11, 
    9.7958938845656736e-11, 9.6936957028909443e-11, 9.5988019168711018e-11, 
    9.5125409891426805e-11, 9.4359851720852589e-11, 9.3699259733572579e-11, 
    9.3148652951731815e-11, 9.2710099511621337e-11, 9.2382799477352285e-11, 
    9.2163182673133807e-11, 9.2045093566784672e-11, 9.2020000686612443e-11, 
    9.2077270402184475e-11, 9.2204445150564271e-11, 9.2387617653096114e-11, 
    9.2611799009434488e-11, 9.2861386438535064e-11, 9.3120634302878102e-11, 
    9.3374184163019729e-11, 9.3607590371791893e-11, 9.3807836066877192e-11, 
    9.3963805340137777e-11, 9.4066680386965405e-11, 9.4110219221995168e-11, 
    9.4090920576241075e-11, 9.4008021090399527e-11, 9.3863374880665111e-11, 
    9.3661165533021987e-11, 9.3407534019145537e-11, 9.3110103922434354e-11, 
    9.2777488017846602e-11, 9.2418760384440575e-11, 9.2042992406293004e-11, 
    9.1658823859227899e-11, 9.1274138432109791e-11, 9.089581805875303e-11, 
    9.0529610422803073e-11, 9.0180045828742264e-11, 8.9850476341672828e-11, 
    8.9543110132149141e-11, 8.9259128416428917e-11, 8.8998763400340327e-11, 
    8.876142281394693e-11, 8.8545761258487101e-11, 8.8349771130757313e-11, 
    8.8170830733302417e-11, 8.8005775652874735e-11, 8.7850951725006836e-11, 
    8.770230024914401e-11, 8.7555457381791041e-11, 8.7405881621150542e-11, 
    8.7249016566019204e-11, 8.7080496375453325e-11, 8.6896313216881564e-11, 
    8.6693046881299538e-11, 8.6468039621043092e-11, 8.6219555049367104e-11, 
    8.5946862033273711e-11, 8.5650274590123069e-11, 8.5331102650608811e-11, 
    8.4991538647960667e-11, 8.4634452217650859e-11, 8.4263167266041914e-11, 
    8.3881157123755966e-11, 8.3491779784673003e-11, 8.3097982657323766e-11, 
    8.2702097676961316e-11, 8.230565241356347e-11, 8.1909297740176004e-11, 
    8.1512797594699424e-11, 8.111511256795363e-11, 8.0714553113825568e-11, 
    8.0308982922047061e-11, 7.9896058426201672e-11, 7.9473470159210927e-11, 
    7.9039162101246881e-11, 7.859152368280415e-11, 7.8129500774506089e-11, 
    7.7652673332537938e-11, 7.716126137548793e-11, 7.6656078250475557e-11, 
    7.6138452963458134e-11, 7.5610138917703575e-11, 7.5073210633762673e-11, 
    7.4529999201224809e-11, 7.3983038335257047e-11, 7.3435053160256926e-11, 
    7.2888974742478903e-11, 7.2347989258751114e-11, 7.1815549451073362e-11, 
    7.1295413545128564e-11, 7.0791604113583185e-11, 7.030834113877938e-11, 
    6.9849887172744201e-11, 6.9420336889984305e-11, 6.9023349184239035e-11, 
    6.866185936425527e-11, 6.8337777114781413e-11, 6.8051754500512815e-11, 
    6.7802997091782338e-11, 6.7589237145843731e-11, 6.7406804737058167e-11, 
    6.7250884272950855e-11, 6.7115882286583739e-11, 6.6995922458344344e-11, 
    6.6885389536202237e-11, 6.6779496283450414e-11, 6.6674760327481653e-11, 
    6.6569386651036369e-11, 6.6463455210094873e-11, 6.6358924018424404e-11, 
    6.6259388997413163e-11, 6.6169676422677877e-11, 6.6095251967912807e-11, 
    6.6041558679756962e-11, 6.6013314416457663e-11, 6.6013901216336265e-11, 
    6.6044832251776637e-11, 6.6105443468546756e-11, 6.6192785571128384e-11, 
    6.6301742368569907e-11, 6.6425335445491004e-11, 6.6555192902845645e-11, 
    6.668211913997585e-11, 6.6796699659677513e-11, 6.6889843833104526e-11, 
    6.6953260033233616e-11, 6.6979798799562807e-11, 6.6963637900009232e-11, 
    6.6900322226535936e-11, 6.6786678679320027e-11, 6.6620645059225863e-11, 
    6.6401046622806805e-11, 6.6127378077450013e-11, 6.5799622153006877e-11, 
    6.5418148304918881e-11, 6.4983696271922022e-11, 6.4497443312549407e-11, 
    6.3961177482425788e-11, 6.3377473117810462e-11, 6.2749913800381755e-11, 
    6.2083284656716605e-11, 6.1383688925456308e-11, 6.0658571304736164e-11, 
    5.9916633243512589e-11, 5.9167602277461645e-11, 5.8421902356962597e-11, 
    5.7690237675135308e-11, 5.6983111694900447e-11, 5.6310336326372109e-11, 
    5.5680574660849814e-11, 5.5100970022980758e-11, 5.457687772254162e-11, 
    5.4111725057140579e-11, 5.3707023251510322e-11, 5.3362484926314696e-11, 
    5.307624644649611e-11, 5.2845163524996914e-11, 5.2665104330882806e-11, 
    5.2531237331004809e-11, 5.2438251172249106e-11, 5.2380511354910335e-11, 
    5.2352131270847717e-11, 5.2346957057429205e-11, 5.2358529588706165e-11, 
    5.2380024537817737e-11, 5.2404229495713166e-11, 5.242357232911464e-11, 
    5.2430253349230456e-11, 5.2416493550479447e-11, 5.237484643813834e-11, 
    5.2298625967639672e-11, 5.2182338176116918e-11, 5.2022108908737242e-11, 
    5.1816047108504869e-11, 5.1564489352337854e-11, 5.1270094145381152e-11, 
    5.0937785325034911e-11, 5.0574501744761997e-11, 5.0188845167032279e-11, 
    4.9790606230305731e-11, 4.9390245747872722e-11, 4.8998382461847094e-11, 
    4.8625343784993184e-11, 4.8280789831377168e-11, 4.7973455198589044e-11, 
    4.7710979750277436e-11, 4.7499864003592164e-11, 4.7345430796229558e-11, 
    4.725184675242636e-11, 4.7222081527390789e-11, 4.7257869942481917e-11, 
    4.7359553624855555e-11, 4.7525904934434722e-11, 4.7753886219748948e-11, 
    4.8038423292980119e-11, 4.837221233958249e-11, 4.8745639505682763e-11, 
    4.9146831162858213e-11, 4.9561882534467458e-11, 4.9975269138532061e-11, 
    5.0370451630167095e-11, 5.0730602431861014e-11, 5.1039452113135146e-11, 
    5.1282144399420605e-11, 5.1446058614075855e-11, 5.1521499647110379e-11, 
    5.150222613277862e-11, 5.1385721103742325e-11, 5.1173234765430845e-11, 
    5.0869560494948663e-11, 5.0482567936701082e-11, 5.0022557607548329e-11, 
    4.9501488129593162e-11, 4.8932140057036023e-11, 4.8327289548998643e-11, 
    4.7698976527650264e-11, 4.7057904868588281e-11, 4.6413034927369663e-11, 
    4.5771382551581362e-11, 4.5138021546500214e-11, 4.4516285241832255e-11, 
    4.3908135559227928e-11, 4.3314614422227963e-11, 4.2736375880985855e-11, 
    4.2174196619791027e-11, 4.1629441283198779e-11, 4.1104387615198906e-11, 
    4.0602447509891027e-11, 4.0128186520487323e-11, 3.9687217152593766e-11, 
    3.9285895842248512e-11, 3.8930948381018434e-11, 3.8628965694665209e-11, 
    3.8385891981437475e-11, 3.8206520269478678e-11, 3.8094065478870019e-11, 
    3.8049788113608825e-11, 3.807283053838951e-11, 3.8160114962904164e-11, 
    3.8306489836312471e-11, 3.8504932301572745e-11, 3.8746971779729873e-11, 
    3.9023116081542147e-11, 3.9323423783843003e-11, 3.9638010083451331e-11, 
    3.9957614934764992e-11, 4.027399306876086e-11, 4.0580316424154132e-11, 
    4.0871336916281961e-11, 4.1143500448324755e-11, 4.1394835336639256e-11, 
    4.1624789484146925e-11, 4.1833874768943213e-11, 4.2023340854714233e-11, 
    4.2194724793601479e-11, 4.2349527790028848e-11, 4.2488847793240701e-11, 
    4.2613214817553965e-11, 4.2722452473770206e-11, 4.2815766413528002e-11, 
    4.2891828247532004e-11, 4.2949072924924059e-11, 4.2985945996212305e-11, 
    4.3001251379300373e-11, 4.2994385413113543e-11, 4.2965588269418995e-11, 
    4.2916005282076343e-11, 4.284774090589227e-11, 4.2763694708397292e-11, 
    4.2667391470257257e-11, 4.2562671573028319e-11, 4.2453392799231872e-11, 
    4.2343074704495449e-11, 4.2234653618595799e-11, 4.2130183702116911e-11, 
    4.2030739541049283e-11, 4.1936321963626738e-11, 4.1845932420458413e-11, 
    4.1757670622572143e-11, 4.166897403215892e-11, 4.157685241865318e-11, 
    4.1478215407765332e-11, 4.1370138193234881e-11, 4.1250190217559525e-11, 
    4.1116633665159677e-11, 4.0968646095519077e-11, 4.0806409673489757e-11, 
    4.063117902582281e-11, 4.0445202922105891e-11, 4.0251648680914651e-11, 
    4.0054371585062155e-11, 3.9857708875377189e-11, 3.966616938495939e-11, 
    3.9484151808048928e-11, 3.9315596746884753e-11, 3.9163705866227929e-11, 
    3.9030643998672126e-11, 3.8917325109502867e-11, 3.8823217153432236e-11, 
    3.874628003056095e-11, 3.8682917636349483e-11, 3.8628105755132514e-11, 
    3.8575560474034462e-11, 3.8518073266070773e-11, 3.8447878347043326e-11, 
    3.8357166047341488e-11, 3.8238601627664696e-11, 3.8085912680590695e-11, 
    3.7894414279491068e-11, 3.7661508971369748e-11, 3.7387033786514416e-11, 
    3.707348346447486e-11, 3.672599875932178e-11, 3.6352172116358265e-11, 
    3.596161846225671e-11, 3.5565377407951468e-11, 3.5175115241934819e-11, 
    3.4802315005243237e-11, 3.4457391084722284e-11, 3.414893752351448e-11, 
    3.3883085770969839e-11, 3.3663128546103147e-11, 3.3489374463350887e-11, 
    3.3359309808576296e-11, 3.3268016932720216e-11, 3.3208833418826462e-11, 
    3.3174127684108531e-11, 3.3156189967920775e-11, 3.3148049580434078e-11, 
    3.3144217925680297e-11, 3.3141191153265327e-11, 3.3137761132258265e-11, 
    3.3135006216752515e-11, 3.313606110701935e-11, 3.3145628695719557e-11, 
    3.316932812588697e-11, 3.3212953445475928e-11, 3.3281711031837696e-11, 
    3.3379495048383563e-11, 3.3508321092692712e-11, 3.3667898734322047e-11, 
    3.3855446158629203e-11, 3.4065689866159694e-11, 3.4291103281922329e-11, 
    3.4522289962362214e-11, 3.4748531179057165e-11, 3.4958403603827511e-11, 
    3.5140457414177391e-11, 3.5283833940472519e-11, 3.5378877146150442e-11, 
    3.5417588896868779e-11, 3.5394007636461798e-11, 3.5304397044058821e-11, 
    3.514732028554205e-11, 3.4923567819923775e-11, 3.4635977756501855e-11, 
    3.4289133106481954e-11, 3.3889040763845539e-11, 3.3442762051343632e-11, 
    3.2958065966169473e-11, 3.2443087747370968e-11, 3.190607939675271e-11, 
    3.1355183277416894e-11, 3.0798291920753243e-11, 3.0242955749085609e-11, 
    2.9696343151225218e-11, 2.9165194634778505e-11, 2.8655828387814127e-11, 
    2.8174105289886292e-11, 2.7725389829551595e-11, 2.7314490279940277e-11, 
    2.6945579089617392e-11, 2.6622096853048427e-11, 2.6346666993575013e-11, 
    2.6121006747219003e-11, 2.5945893651244969e-11, 2.5821147350900182e-11, 
    2.5745671039886985e-11, 2.5717547615506501e-11, 2.57341762397277e-11, 
    2.5792436672074984e-11, 2.5888899169316496e-11, 2.6020019643235499e-11, 
    2.6182330477799854e-11, 2.6372601739356553e-11, 2.6587963908239752e-11, 
    2.6825960270035492e-11, 2.7084561150954838e-11, 2.7362105876358836e-11, 
    2.7657212166343014e-11, 2.7968633641136804e-11, 2.8295121558282477e-11, 
    2.8635266740374177e-11, 2.8987365616880853e-11, 2.9349325114072638e-11, 
    2.9718605698683027e-11, 3.0092197420319522e-11, 3.0466664917947741e-11, 
    3.0838209739907791e-11, 3.1202776299008737e-11, 3.1556155854812344e-11, 
    3.1894097529758277e-11, 3.2212417496600288e-11, 3.2507069907497376e-11, 
    3.2774195284595676e-11, 3.3010155420372932e-11, 3.3211524561360134e-11, 
    3.3375081442249939e-11, 3.3497792472692935e-11, 3.357681874417561e-11, 
    3.3609499457108901e-11, 3.3593420941088967e-11, 3.3526477274523094e-11, 
    3.3406986152634587e-11, 3.3233835728243564e-11, 3.3006663956344332e-11, 
    3.2726026772401533e-11, 3.2393603053203129e-11, 3.201233636145346e-11, 
    3.15865741697777e-11, 3.1122103863832091e-11, 3.0626162029468648e-11, 
    3.0107290004387113e-11, 2.957513671211228e-11, 2.9040149548065824e-11, 
    2.851319408663416e-11, 2.8005066183598864e-11, 2.752601006233344e-11, 
    2.7085209611288473e-11, 2.6690324493697013e-11, 2.6347073631021656e-11, 
    2.6058950017018759e-11, 2.5827042868361361e-11, 2.5650010810989883e-11, 
    2.5524229120089766e-11, 2.5444073088018448e-11, 2.5402301644005037e-11, 
    2.5390586801794977e-11, 2.5400072333475971e-11, 2.5421974412559998e-11, 
    2.544812739692277e-11, 2.5471479172596638e-11, 2.548648305081828e-11, 
    2.5489353374010475e-11, 2.5478153140083136e-11, 2.5452762059042344e-11, 
    2.5414679300485011e-11, 2.536671635255713e-11, 2.5312597178114783e-11, 
    2.5256516419349885e-11, 2.5202681047900444e-11, 2.5154885348960143e-11, 
    2.5116166525349383e-11, 2.5088546583485522e-11, 2.5072880774771107e-11, 
    2.5068847863541893e-11, 2.5075023713019521e-11, 2.5089086113559196e-11, 
    2.510806696390536e-11, 2.5128656935037531e-11, 2.5147518001353003e-11, 
    2.5161583931422201e-11, 2.5168280263486898e-11, 2.5165706919800315e-11, 
    2.5152721002947098e-11, 2.5128951809843586e-11, 2.5094706592625074e-11, 
    2.5050859403843096e-11, 2.4998670442781719e-11, 2.493961187303448e-11, 
    2.4875189284469026e-11, 2.4806803877829575e-11, 2.4735644885906102e-11, 
    2.4662651296050433e-11, 2.4588476475232169e-11, 2.4513520778768734e-11, 
    2.443795181295787e-11, 2.4361741236015506e-11, 2.4284652414977782e-11, 
    2.4206234812977485e-11, 2.4125745702067413e-11, 2.4042093386979982e-11, 
    2.3953730057003226e-11, 2.3858599987378143e-11, 2.3754091382554514e-11, 
    2.363708610761402e-11, 2.3504045953625236e-11, 2.3351224481593911e-11, 
    2.3174893360024439e-11, 2.297166766477722e-11, 2.2738813729076007e-11, 
    2.2474557280642014e-11, 2.217831877440529e-11, 2.1850893299005179e-11, 
    2.14944856914761e-11, 2.1112671368736259e-11, 2.0710232773605065e-11, 
    2.0292953355307901e-11, 1.9867296964756825e-11, 1.9440128784613645e-11, 
    1.9018422341832653e-11, 1.8609017606126887e-11, 1.8218407896264008e-11, 
    1.7852618518023404e-11, 1.7517093380418008e-11, 1.7216651767145697e-11, 
    1.6955423977917716e-11, 1.6736810023128841e-11, 1.6563397391854183e-11, 
    1.6436879378096482e-11, 1.6357929424401223e-11, 1.6326096676285186e-11, 
    1.6339704556836969e-11, 1.6395818681127383e-11, 1.6490247515480288e-11, 
    1.6617671153848236e-11, 1.6771845994403386e-11, 1.6945910975965791e-11, 
    1.7132771038460108e-11, 1.7325541920297017e-11, 1.751797903635624e-11, 
    1.770490742900988e-11, 1.7882555694632615e-11, 1.8048802819853713e-11, 
    1.8203264300428731e-11, 1.8347262187205554e-11, 1.8483631287495484e-11, 
    1.8616434119376524e-11, 1.8750541758744819e-11, 1.8891207410822613e-11, 
    1.9043597897121514e-11, 1.921238143023756e-11, 1.9401362693842264e-11, 
    1.9613204065188726e-11, 1.9849261518178711e-11, 2.0109502782097775e-11, 
    2.0392509729706726e-11, 2.0695557849586274e-11, 2.1014740537293147e-11, 
    2.1345126714562163e-11, 2.168092343980175e-11, 2.2015661030439682e-11, 
    2.2342371235165082e-11, 2.2653783845936665e-11, 2.2942528796664804e-11, 
    2.3201353381552539e-11, 2.3423381248735975e-11, 2.360236108374902e-11, 
    2.3732928734414587e-11, 2.3810860728586356e-11, 2.3833279882098122e-11, 
    2.3798810868081598e-11, 2.370767358622118e-11, 2.3561680486438217e-11, 
    2.336414584549124e-11, 2.3119726100091963e-11, 2.2834207796951603e-11, 
    2.2514228930740807e-11, 2.2167030025479241e-11, 2.1800186487135945e-11, 
    2.1421384134964795e-11, 2.1038244850907749e-11, 2.0658181908516012e-11, 
    2.0288301417284973e-11, 1.9935342818435944e-11, 1.9605600110586471e-11, 
    1.930486572771356e-11, 1.9038334592575128e-11, 1.8810497445911891e-11, 
    1.8624996342815956e-11, 1.8484486797463369e-11, 1.8390497446096556e-11, 
    1.8343319157193195e-11, 1.8341933951634203e-11, 1.8384049802621481e-11, 
    1.8466192044537395e-11, 1.8583877289127869e-11, 1.8731884898693438e-11, 
    1.8904588307045511e-11, 1.9096300324562974e-11, 1.9301638068438871e-11, 
    1.9515827670439563e-11, 1.9734948782755174e-11, 1.9956064926942718e-11, 
    2.0177247569057677e-11, 2.0397464818438213e-11, 2.0616376717674683e-11, 
    2.0834047844952169e-11, 2.1050605114864414e-11, 2.1265903612802053e-11, 
    2.1479248800940752e-11, 2.1689198415254333e-11, 2.1893471308020646e-11, 
    2.2089001675645851e-11, 2.227213150579978e-11, 2.2438877687241395e-11, 
    2.2585332504068469e-11, 2.2708057874104437e-11, 2.2804442643364201e-11, 
    2.2873028051845782e-11, 2.291368728195936e-11, 2.2927664553818934e-11, 
    2.2917470337907103e-11, 2.2886610164146415e-11, 2.2839215420018651e-11, 
    2.2779592298077488e-11, 2.2711755753629441e-11, 2.2639014190162275e-11, 
    2.2563653183302419e-11, 2.2486760461384529e-11, 2.2408207102744193e-11, 
    2.232680798260258e-11, 2.2240595346600402e-11, 2.214721613714253e-11, 
    2.2044336904012894e-11, 2.1930043938719447e-11, 2.1803160447032757e-11, 
    2.166343668168529e-11, 2.1511567785697623e-11, 2.1349084369806664e-11, 
    2.117810022362424e-11, 2.1000965994102367e-11, 2.0819895983558622e-11, 
    2.0636631587947507e-11, 2.0452154699741911e-11, 2.0266562858498085e-11, 
    2.0079071576426494e-11, 1.9888164179167148e-11, 1.9691876602514209e-11, 
    1.9488150249487244e-11, 1.9275221948898134e-11, 1.9051972820021053e-11, 
    1.8818205811101007e-11, 1.8574796171803597e-11, 1.832368187688407e-11, 
    1.8067729209659628e-11, 1.7810466256111288e-11, 1.7555744372624304e-11, 
    1.7307340588983569e-11, 1.7068604689490655e-11, 1.684216788226353e-11, 
    1.6629761625033965e-11, 1.6432145295474559e-11, 1.6249203749465971e-11, 
    1.6080115780468812e-11, 1.5923635200559668e-11, 1.5778404740120411e-11, 
    1.5643267183887827e-11, 1.5517521139830358e-11, 1.5401090989725957e-11, 
    1.5294596880127536e-11, 1.5199306864322499e-11, 1.5116957666638491e-11, 
    1.504951786561012e-11, 1.4998862536800076e-11, 1.4966438055873365e-11, 
    1.4952954759612584e-11, 1.4958125736796189e-11, 1.4980484987175503e-11, 
    1.5017333769244455e-11, 1.5064779786823488e-11, 1.5117917347802695e-11, 
    1.5171094190034454e-11, 1.5218251296469705e-11, 1.525334354394915e-11, 
    1.5270752339126933e-11, 1.5265678540641871e-11, 1.52344937873e-11, 
    1.5175007621875108e-11, 1.5086625973790101e-11, 1.4970384531535657e-11, 
    1.4828855250107946e-11, 1.4665941417237803e-11, 1.4486547605027294e-11, 
    1.4296183853753832e-11, 1.4100515160064234e-11, 1.3904903494915985e-11, 
    1.3713995644722938e-11, 1.3531376757126842e-11, 1.3359351740984921e-11, 
    1.3198869003003627e-11, 1.3049587023670221e-11, 1.2910115698955774e-11, 
    1.2778353357179417e-11, 1.2651942700454187e-11, 1.2528748086295489e-11, 
    1.240731043496814e-11, 1.2287245070392832e-11, 1.2169493605565394e-11, 
    1.2056427767989386e-11, 1.1951782749415731e-11, 1.1860420145065344e-11, 
    1.1787950586140918e-11, 1.174028287799917e-11, 1.1723115895396237e-11, 
    1.1741450735617611e-11, 1.1799208598261833e-11, 1.1898932211237979e-11, 
    1.2041626178791501e-11, 1.2226759419758076e-11, 1.2452369066235995e-11, 
    1.2715278644207859e-11, 1.3011372542414758e-11, 1.3335878988548517e-11, 
    1.3683644527475415e-11, 1.404936301186926e-11, 1.442773526000779e-11, 
    1.4813545425041587e-11, 1.5201729238575807e-11, 1.5587361672107441e-11, 
    1.5965629224884564e-11, 1.6331818877832206e-11, 1.6681333149865211e-11, 
    1.7009724964878784e-11, 1.7312771407180151e-11, 1.7586572145528612e-11, 
    1.7827668529943405e-11, 1.8033154239079282e-11, 1.8200762860302527e-11, 
    1.8328910447009964e-11, 1.8416708468348292e-11, 1.8463908973146442e-11, 
    1.8470820625152527e-11, 1.8438188569870022e-11, 1.8367078816543215e-11, 
    1.825876940216365e-11, 1.8114677127067041e-11, 1.7936348117176538e-11, 
    1.7725481809785132e-11, 1.7484040482438849e-11, 1.7214367485056025e-11, 
    1.6919337805615009e-11, 1.6602493745515938e-11, 1.6268123325858769e-11, 
    1.5921281931756803e-11, 1.5567705488033909e-11, 1.5213632944985612e-11, 
    1.4865515836992272e-11, 1.4529687530274627e-11, 1.4211963935385578e-11, 
    1.3917260267088941e-11, 1.3649268736989666e-11, 1.3410213944672273e-11, 
    1.3200764867501052e-11, 1.3020081805294836e-11, 1.2866026541530007e-11, 
    1.2735513178691224e-11, 1.2624951522763991e-11, 1.2530760316483773e-11, 
    1.2449847730348503e-11, 1.2380056083271764e-11, 1.2320455697061483e-11, 
    1.2271492900896324e-11, 1.2234945783439632e-11, 1.2213690722119524e-11, 
    1.2211309187024356e-11, 1.2231562679956417e-11, 1.2277789094356783e-11, 
    1.2352330398164579e-11, 1.2456015272322005e-11, 1.2587742487517076e-11, 
    1.2744289265441404e-11, 1.2920312876503995e-11, 1.3108570833994869e-11, 
    1.3300347745165476e-11, 1.3486043053899734e-11, 1.3655859103638575e-11, 
    1.3800536717665046e-11, 1.3912027769728501e-11, 1.3984085184621098e-11, 
    1.4012649380974064e-11, 1.3996055727094187e-11, 1.3935005743152725e-11, 
    1.3832322710865257e-11, 1.3692539701990879e-11, 1.3521365896459897e-11, 
    1.3325077735663199e-11, 1.3109950301461217e-11, 1.2881751362744425e-11, 
    1.2645384150180199e-11, 1.2404680944149973e-11, 1.2162421682670516e-11, 
    1.1920472194463446e-11, 1.1680094899967339e-11, 1.1442363693328941e-11, 
    1.120860277506806e-11, 1.0980787622380214e-11, 1.0761890937675138e-11, 
    1.0556097262100737e-11, 1.0368853950994384e-11, 1.0206751241018998e-11, 
    1.0077250500765399e-11, 9.9882425343780052e-12, 9.9475117152278232e-12, 
    9.9621336624612782e-12, 1.0037857076735683e-11, 1.017852108494598e-11, 
    1.038557598648119e-11, 1.0657732188244351e-11, 1.0990771900169778e-11, 
    1.1377573132061694e-11, 1.1808321322816185e-11, 1.2270888179667189e-11, 
    1.2751417208744272e-11, 1.3235006284062641e-11, 1.3706494506762442e-11, 
    1.4151264995557812e-11, 1.4556038598043301e-11, 1.4909568341971726e-11, 
    1.5203228437416577e-11, 1.543141290429161e-11, 1.5591760841184208e-11, 
    1.5685150524221695e-11, 1.5715539817030019e-11, 1.5689552461468828e-11, 
    1.5615957595620543e-11, 1.5505031552543434e-11, 1.5367835916042475e-11, 
    1.5215472821765039e-11, 1.5058384859746253e-11, 1.4905718298216486e-11, 
    1.4764809288682919e-11, 1.4640811749291331e-11, 1.4536507719026822e-11, 
    1.4452286197084258e-11, 1.4386314086042821e-11, 1.4334885723569555e-11, 
    1.4292911220269814e-11, 1.4254514793460714e-11, 1.4213704294839184e-11, 
    1.4165050312843067e-11, 1.4104307460968044e-11, 1.4028954833046211e-11, 
    1.3938570013368278e-11, 1.3835012776271036e-11, 1.3722401695416197e-11, 
    1.3606892071138552e-11, 1.3496251330170391e-11, 1.3399282309204376e-11, 
    1.3325145071347883e-11, 1.3282651220921364e-11, 1.3279577956573501e-11, 
    1.3322063836868593e-11, 1.3414152428864505e-11, 1.3557491420280429e-11, 
    1.3751222281524161e-11, 1.3992041686231471e-11, 1.4274421319593919e-11, 
    1.4590939853543913e-11, 1.4932703678824884e-11, 1.528979981588667e-11, 
    1.5651764706784771e-11, 1.6008010351330631e-11, 1.6348221758753555e-11, 
    1.6662705072187087e-11, 1.6942688495737357e-11, 1.7180586358540565e-11, 
    1.7370236564024863e-11, 1.7507115363918577e-11, 1.758851545958517e-11, 
    1.7613726063867384e-11, 1.7584129098886661e-11, 1.750325591630002e-11, 
    1.7376740205589296e-11, 1.7212166876639852e-11, 1.7018795376502858e-11, 
    1.68071558696224e-11, 1.6588527666332971e-11, 1.637431913486678e-11, 
    1.6175391504985532e-11, 1.6001371178315544e-11, 1.5860008109771264e-11, 
    1.5756612473941476e-11, 1.5693639138714738e-11, 1.5670467453824976e-11, 
    1.5683372618185533e-11, 1.5725713652122525e-11, 1.5788318450436107e-11, 
    1.5860070279203868e-11, 1.5928620915692051e-11, 1.5981168813739007e-11, 
    1.6005284296190381e-11, 1.5989703041400465e-11, 1.5924999845768991e-11, 
    1.5804152713608807e-11, 1.5622904047952952e-11, 1.5379934041491674e-11, 
    1.5076848105159004e-11, 1.4717956063162269e-11, 1.4309895559069678e-11, 
    1.386116969403345e-11, 1.338158105095856e-11, 1.2881647516452782e-11, 
    1.2372049037081173e-11, 1.1863127883007803e-11, 1.1364473365087966e-11, 
    1.0884615672578338e-11, 1.0430805782579461e-11, 1.0008921501615478e-11, 
    9.6234305869815999e-12, 9.2774479426165433e-12, 8.9728185642462014e-12, 
    8.7102545089893705e-12, 8.4894718296789092e-12, 8.3093657696837471e-12, 
    8.1681658635019596e-12, 8.0636235625278026e-12, 7.9931823747578871e-12, 
    7.9541782022040556e-12, 7.9440006726497752e-12, 7.9602790772896969e-12, 
    8.0010025142707544e-12, 8.0646269894234114e-12, 8.1500910890956979e-12, 
    8.2567874946587261e-12, 8.384437192381363e-12, 8.5329100226954319e-12, 
    8.7019619733745002e-12, 8.8910059198946309e-12, 9.0988061000292585e-12, 
    9.3233117108695769e-12, 9.5615203307511477e-12, 9.8094489853441591e-12, 
    1.0062268738897407e-11, 1.0314545432076222e-11, 1.0560588585411986e-11, 
    1.0794885485676419e-11, 1.1012543436777153e-11, 1.1209723045732651e-11, 
    1.138396694428844e-11, 1.1534425116355703e-11, 1.1661883786593273e-11, 
    1.1768671142600241e-11, 1.1858360898809608e-11, 1.1935360903545048e-11, 
    1.2004415250128089e-11, 1.2070075218717116e-11, 1.2136205303428175e-11, 
    1.2205580474188498e-11, 1.2279623571278859e-11, 1.2358298114202823e-11, 
    1.2440195116662624e-11, 1.2522777464387251e-11, 1.2602763501695251e-11, 
    1.267662256318761e-11, 1.274108391727646e-11, 1.2793657712866171e-11, 
    1.2833061284456931e-11, 1.2859522639526689e-11, 1.2874937050414203e-11, 
    1.2882823341103186e-11, 1.2888107503618726e-11, 1.2896736318887424e-11, 
    1.2915137278232871e-11, 1.2949615160529475e-11, 1.3005703752533047e-11, 
    1.3087532564411217e-11, 1.319730243083851e-11, 1.3334906467325748e-11, 
    1.3497735102211832e-11, 1.3680688148835053e-11, 1.3876422117932567e-11, 
    1.407579497799157e-11, 1.4268482757489213e-11, 1.4443715784119207e-11, 
    1.4591075272534355e-11, 1.4701252476089508e-11, 1.4766751494909731e-11, 
    1.4782414897567696e-11, 1.474578107893618e-11, 1.4657204030189959e-11, 
    1.4519758468977404e-11, 1.4338916927680895e-11, 1.4122069274898535e-11, 
    1.3877899197051598e-11, 1.3615706097204769e-11, 1.3344704581685392e-11, 
    1.3073395797310201e-11, 1.2809025756851381e-11, 1.2557205744776331e-11, 
    1.232167694863983e-11, 1.2104270879930972e-11, 1.1905024905174139e-11, 
    1.1722455832187708e-11, 1.1553930957029719e-11, 1.1396133083798202e-11, 
    1.1245545653699889e-11, 1.1098924791369439e-11, 1.0953718659852456e-11, 
    1.0808402919447808e-11, 1.0662677211194818e-11, 1.0517550883217366e-11, 
    1.0375279232306084e-11, 1.0239177993092585e-11, 1.011331664494939e-11, 
    1.0002156586739767e-11, 9.9101166444035939e-12, 9.8411678724349159e-12, 
    9.7984492492126397e-12, 9.7839764785264209e-12,
  // Sqw-Na(3, 0-1999)
    0.059405377288691802, 0.05931005751740076, 0.059026135860628076, 
    0.058559625953951353, 0.057920227051748062, 0.057120864780751006, 
    0.056177097325443952, 0.0551064300396771, 0.053927585906342501, 
    0.052659779236272186, 0.051322035828941855, 0.049932595282952914, 
    0.048508421329666811, 0.047064835199158571, 0.045615276315099283, 
    0.044171185077130928, 0.042741994865018708, 0.041335215094119034, 
    0.039956584243804417, 0.03861027106966796, 0.037299103301300554, 
    0.036024805523222722, 0.034788231126490599, 0.033589576747514338, 
    0.032428571121488212, 0.0313046335256493, 0.030216999830662266, 
    0.029164816553881673, 0.028147205201967396, 0.0271633006103153, 
    0.026212267945811354, 0.025293303549616904, 0.024405624874228888, 
    0.023548454444978682, 0.022721002107218224, 0.021922448894948224, 
    0.021151934791170408, 0.020408551577403983, 0.019691341018704556, 
    0.018999297905018378, 0.018331377029740154, 0.017686503037628743, 
    0.017063582169080566, 0.016461515177513208, 0.015879210992771269, 
    0.015315600942781574, 0.014769653453200214, 0.014240389089588235, 
    0.013726895606699862, 0.013228342384888896, 0.012743993350202409, 
    0.012273217281967704, 0.011815494380801482, 0.011370418136873138, 
    0.010937691895170579, 0.010517120011973838, 0.010108594054710198, 
    0.0097120750227721684, 0.0093275729730655683, 0.0089551256579714651, 
    0.0085947777967918578, 0.0082465624145452079, 0.0079104853376339365, 
    0.0075865135004903094, 0.0072745672650394132, 0.0069745165535550846, 
    0.0066861802950104856, 0.006409328510386861, 0.0061436863129315242, 
    0.0058889391530084984, 0.0056447387584516425, 0.0054107093706858411, 
    0.0051864540193987986, 0.0049715606900611843, 0.0047656083083226913, 
    0.0045681724950323282, 0.0043788310460685922, 0.0041971690770567947, 
    0.0040227837582192325, 0.0038552885583841043, 0.0036943169228184792, 
    0.0035395253247672447, 0.0033905956496645415, 0.0032472368877039109, 
    0.003109186120650826, 0.0029762087920043897, 0.0028480982492615583, 
    0.0027246745491714729, 0.0026057825280669973, 0.002491289164385476, 
    0.0023810803004097516, 0.0022750568416413089, 0.0021731306075382885, 
    0.0020752200565659221, 0.0019812461412628737, 0.0018911285570334107, 
    0.0018047826272651467, 0.0017221170177153854, 0.0016430324003160446, 
    0.0015674210998313186, 0.0014951676674172468, 0.0014261502443835732, 
    0.001360242516840932, 0.0012973160237979835, 0.0012372425702200014, 
    0.0011798965114314464, 0.0011251567118135749, 0.0010729080327510328, 
    0.0010230422650383229, 0.00097545848244027817, 0.00093006284971842957, 
    0.00088676796553642501, 0.00084549185520023352, 0.00080615674870440309, 
    0.0007686877859287973, 0.00073301178405861588, 0.00069905618421753411, 
    0.0006667482673740683, 0.00063601469669454696, 0.00060678140783136951, 
    0.00057897383338078212, 0.00055251741602405004, 0.00052733833940821575, 
    0.00050336438875229822, 0.00048052584577095364, 0.0004587563251085739, 
    0.00043799347135244521, 0.00041817945517369048, 0.00039926123177883688, 
    0.00038119055172367098, 0.00036392374018745651, 0.0003474212832190418, 
    0.0003316472759922447, 0.00031656879731115051, 0.00030215527598690588, 
    0.00028837790872850464, 0.00027520917714059158, 0.00026262249522315703, 
    0.00025059200067414314, 0.00023909248559995824, 0.0002280994469686211, 
    0.00021758922583842101, 0.00020753919795437776, 0.00019792797693151651, 
    0.0001887355944897635, 0.00017994362911454167, 0.00017153526379910276, 
    0.00016349526378027767, 0.00015580987508864824, 0.0001484666532308277, 
    0.00014145423768224553, 0.00013476209176208683, 0.00012838022890593516, 
    0.00012229894565410273, 0.00011650857931326946, 0.00011099930478338643, 
    0.00010576098099640033, 0.00010078305323163938, 9.6054513568262243e-05, 
    9.1563918104020344e-05, 8.7299456402170335e-05, 8.3249065957623046e-05, 
    7.9400582303512936e-05, 7.574191372593429e-05, 7.2261228451914969e-05, 
    6.8947141685448736e-05, 6.578889005406188e-05, 6.2776481949649958e-05, 
    5.9900813911361267e-05, 5.7153745559931324e-05, 5.4528128527653137e-05, 
    5.2017788147091367e-05, 4.9617460113070165e-05, 4.732268763675564e-05, 
    4.5129687479684191e-05, 4.3035195434981048e-05, 4.1036303109274108e-05, 
    3.9130298134481125e-05, 3.7314519173586516e-05, 3.5586235354590561e-05, 
    3.3942557234972325e-05, 3.2380383315919761e-05, 3.089638279219506e-05, 
    2.9487011975330694e-05, 2.8148558986932665e-05, 2.6877209169986538e-05, 
    2.5669122410387258e-05, 2.4520513302132457e-05, 2.3427725806142704e-05, 
    2.2387295611469661e-05, 2.1395995568199861e-05, 2.0450862021335368e-05, 
    1.954920230107668e-05, 1.8688585713310594e-05, 1.7866821882857749e-05, 
    1.7081931095816446e-05, 1.6332111342363645e-05, 1.5615706171904679e-05, 
    1.4931176417113485e-05, 1.4277077558325768e-05, 1.3652043223278439e-05, 
    1.3054774257926557e-05, 1.2484032097765636e-05, 1.1938634871376456e-05, 
    1.1417454745275089e-05, 1.0919415376204483e-05, 1.0443488835380599e-05, 
    9.9886918706341347e-06, 9.5540817601548364e-06, 9.1387522201315353e-06, 
    8.7418298438157747e-06, 8.3624714112200326e-06, 7.9998621857662453e-06, 
    7.6532150911712544e-06, 7.3217705071714841e-06, 7.0047963800574249e-06, 
    6.7015884156173942e-06, 6.4114702792802559e-06, 6.1337939131281051e-06, 
    5.8679402311599284e-06, 5.6133205163967701e-06, 5.3693787884214238e-06, 
    5.1355952367993387e-06, 4.911490558630529e-06, 4.6966307503656735e-06, 
    4.4906316515716663e-06, 4.2931623797400957e-06, 4.1039467738929743e-06, 
    3.9227620939974859e-06, 3.749434490876674e-06, 3.5838311262356301e-06, 
    3.4258492301787828e-06, 3.2754027707249553e-06, 3.1324077219207602e-06, 
    2.9967671111212579e-06, 2.8683570824049447e-06, 2.747015130093123e-06, 
    2.6325314547609182e-06, 2.5246441039322076e-06, 2.4230382214214171e-06, 
    2.3273493805128485e-06, 2.2371706524380217e-06, 2.1520627878843866e-06, 
    2.0715666844817458e-06, 1.9952171846827903e-06, 1.9225571995342587e-06, 
    1.8531511800934447e-06, 1.7865970537393608e-06, 1.7225358964507685e-06, 
    1.6606588130392109e-06, 1.6007107291020588e-06, 1.5424910447640082e-06, 
    1.4858513403548722e-06, 1.4306905392246617e-06, 1.3769481022157549e-06, 
    1.3245959383846058e-06, 1.2736297564757684e-06, 1.2240605515111073e-06, 
    1.175906826217397e-06, 1.1291880044169789e-06, 1.0839193217390058e-06, 
    1.0401083029016092e-06, 9.9775277463314972e-07, 9.5684023831974027e-07, 
    9.1734834506974059e-07, 8.7924618256960288e-07, 8.4249609021854465e-07, 
    8.0705575686701868e-07, 7.7288040804278482e-07, 7.3992494343960518e-07, 
    7.0814592778388155e-07, 6.775033640125346e-07, 6.4796218465156032e-07, 
    6.1949339220790987e-07, 5.9207476909392173e-07, 5.6569107429520777e-07, 
    5.4033365470086062e-07, 5.1599943108390535e-07, 4.9268927066163247e-07, 
    4.7040582649245303e-07, 4.4915099724760815e-07, 4.2892322785573628e-07, 
    4.0971491780320077e-07, 3.9151022018586189e-07, 3.7428349346075861e-07, 
    3.5799861095374225e-07, 3.4260924485705878e-07, 3.2806013518738148e-07, 
    3.1428924297564314e-07, 3.0123058760224558e-07, 2.8881749318819799e-07, 
    2.7698592851701276e-07, 2.6567762203533417e-07, 2.5484266749860146e-07, 
    2.4444139853093436e-07, 2.3444539352908508e-07, 2.2483756233904708e-07, 
    2.1561135420586582e-07, 2.067692013536213e-07, 1.9832037036756654e-07, 
    1.902784290777811e-07, 1.8265855183931455e-07, 1.754748807109792e-07, 
    1.687381391023014e-07, 1.6245365968151571e-07, 1.5661994526906724e-07, 
    1.5122783213561493e-07, 1.4626027469038614e-07, 1.4169272117045248e-07, 
    1.374940068627665e-07, 1.3362765623738761e-07, 1.3005346283429655e-07, 
    1.2672920585055001e-07, 1.2361236708924682e-07, 1.206617284027686e-07, 
    1.1783875649488787e-07, 1.1510871330916765e-07, 1.1244146300435785e-07, 
    1.098119748452153e-07, 1.0720054343721937e-07, 1.0459276046712659e-07, 
    1.0197927745101925e-07, 9.9355397007374907e-08, 9.6720525710259765e-08, 
    9.4077516164894043e-08, 9.1431923897582808e-08, 8.879120566452524e-08, 
    8.6163891440188218e-08, 8.355876937883171e-08, 8.0984130357448844e-08, 
    7.8447121802062039e-08, 7.595325861016303e-08, 7.3506129164750279e-08, 
    7.1107318718267771e-08, 6.8756551045885109e-08, 6.64520268330583e-08, 
    6.4190915851036122e-08, 6.196994459722783e-08, 5.978601237679421e-08, 
    5.7636769755068202e-08, 5.5521101516972451e-08, 5.3439471730585525e-08, 
    5.1394106705828714e-08, 4.9389011178577587e-08, 4.7429829602414733e-08, 
    4.552357754645582e-08, 4.3678275359400792e-08, 4.1902519282255992e-08, 
    4.0205023135898766e-08, 3.859415982620973e-08, 3.7077525896897182e-08, 
    3.5661547184382744e-08, 3.4351138432420092e-08, 3.3149426472693769e-08, 
    3.2057543663369435e-08, 3.1074496854076976e-08, 3.0197115358783214e-08, 
    2.9420080349935705e-08, 2.8736036011152262e-08, 2.8135781093124388e-08, 
    2.7608536731826474e-08, 2.7142283911734072e-08, 2.6724160588332872e-08, 
    2.6340905598122602e-08, 2.5979332780953545e-08, 2.5626815948962866e-08, 
    2.527176219425671e-08, 2.4904049418824217e-08, 2.4515402887444327e-08, 
    2.4099686963423017e-08, 2.3653090736575694e-08, 2.3174191628579303e-08, 
    2.2663887751524524e-08, 2.2125198587522032e-08, 2.1562942574611631e-08, 
    2.0983309948673287e-08, 2.0393357282507187e-08, 1.9800457302325268e-08, 
    1.9211741561303406e-08, 1.8633575254692259e-08, 1.8071101483818615e-08, 
    1.7527887726683452e-08, 1.7005699508722837e-08, 1.6504416910902464e-08, 
    1.6022098287819315e-08, 1.5555184402665499e-08, 1.5098825077443037e-08, 
    1.4647301339334129e-08, 1.4194508759655916e-08, 1.3734463866708796e-08, 
    1.3261794498517034e-08, 1.2772177928125265e-08, 1.2262695870809042e-08, 
    1.1732083839737228e-08, 1.1180861630075657e-08, 1.0611341878843198e-08, 
    1.0027522906773925e-08, 9.4348802548199323e-09, 8.8400768898811076e-09, 
    8.2506156597421971e-09, 7.6744583656811717e-09, 7.1196349171202296e-09, 
    6.5938632192376928e-09, 6.1041973372505276e-09, 5.6567176941668505e-09, 
    5.2562740689288212e-09, 4.9062893334275057e-09, 4.6086298882418547e-09, 
    4.3635467750598681e-09, 4.1696897175258452e-09, 4.0241937762853488e-09, 
    3.9228355858349368e-09, 3.8602522162938116e-09, 3.8302119431704238e-09, 
    3.8259219342811602e-09, 3.8403548152023676e-09, 3.8665738580953195e-09, 
    3.8980364421968029e-09, 3.928857003212245e-09, 3.9540146085162395e-09, 
    3.9694951489955361e-09, 3.9723644701634798e-09, 3.9607745569901799e-09, 
    3.9339104371550715e-09, 3.8918892236858673e-09, 3.8356251236317684e-09, 
    3.7666743561330921e-09, 3.6870730003019812e-09, 3.5991781255146931e-09, 
    3.5055199564360592e-09, 3.4086696997714846e-09, 3.3111255297190655e-09, 
    3.2152173886263472e-09, 3.1230306790060278e-09, 3.0363485053143431e-09, 
    2.9566125130069798e-09, 2.8849023167348967e-09, 2.8219335799074226e-09, 
    2.7680740053695867e-09, 2.7233757011956706e-09, 2.6876207817394053e-09, 
    2.6603760137785921e-09, 2.641050925293152e-09, 2.628953652900695e-09, 
    2.6233388095756514e-09, 2.6234429825505087e-09, 2.628505048264112e-09, 
    2.6377709408617391e-09, 2.6504845692875498e-09, 2.6658688838407501e-09, 
    2.6831022516774357e-09, 2.7012963394149666e-09, 2.7194810243333517e-09, 
    2.7366013161749129e-09, 2.75152907925591e-09, 2.7630906873950356e-09, 
    2.7701091850415485e-09, 2.7714578568821055e-09, 2.7661202447154922e-09, 
    2.7532510201253602e-09, 2.73223157625538e-09, 2.7027149610548966e-09, 
    2.664655541373371e-09, 2.6183206280622399e-09, 2.5642827572036808e-09, 
    2.5033935061492374e-09, 2.4367410844496116e-09, 2.3655956168167179e-09, 
    2.2913466183552016e-09, 2.2154378320091204e-09, 2.139304136932864e-09, 
    2.0643148977323396e-09, 1.9917267892206628e-09, 1.9226482648184825e-09, 
    1.8580162341940707e-09, 1.7985846250650013e-09, 1.7449232674549649e-09, 
    1.6974251429440169e-09, 1.6563194353947945e-09, 1.6216881234305071e-09, 
    1.5934837948723739e-09, 1.5715472036366553e-09, 1.5556233460077336e-09, 
    1.5453757159516551e-09, 1.5403986869966221e-09, 1.5402285721845863e-09, 
    1.544353937239516e-09, 1.5522259266084553e-09, 1.5632690941158721e-09, 
    1.5768931236563784e-09, 1.5925053090818867e-09, 1.6095236160838884e-09, 
    1.6273895897040918e-09, 1.645580487414192e-09, 1.6636197558265407e-09, 
    1.6810851917602884e-09, 1.6976141844694801e-09, 1.7129058089561644e-09, 
    1.726719626433111e-09, 1.7388715298905748e-09, 1.7492269326831842e-09, 
    1.7576920162496742e-09, 1.7642036155361417e-09, 1.7687185699957887e-09, 
    1.7712031448950514e-09, 1.7716233102490833e-09, 1.7699364385483202e-09, 
    1.7660850165583453e-09, 1.759992836957416e-09, 1.7515641110286957e-09, 
    1.740685733485373e-09, 1.7272328971946713e-09, 1.7110779022594426e-09, 
    1.6921019526355438e-09, 1.6702092659533872e-09, 1.6453427407469032e-09, 
    1.6174999766032521e-09, 1.5867484769524937e-09, 1.5532385014475794e-09, 
    1.5172123196223087e-09, 1.4790085093154307e-09, 1.4390604441004299e-09, 
    1.3978883383105906e-09, 1.3560848685341887e-09, 1.3142947408778779e-09, 
    1.273189325946861e-09, 1.2334377668559062e-09, 1.1956764813824188e-09, 
    1.1604790770903748e-09, 1.1283289147621951e-09, 1.0995962278242455e-09, 
    1.0745215929937511e-09, 1.0532068590507889e-09, 1.0356143085060108e-09, 
    1.0215739541539137e-09, 1.0107984246375042e-09, 1.0029041759114186e-09, 
    9.9743742861961355e-10, 9.9390277997729123e-10, 9.9179244383720862e-10, 
    9.9061400616010541e-10, 9.899148935300092e-10, 9.8930201502819824e-10, 
    9.8845561152657754e-10, 9.8713674682859322e-10, 9.8518853446113337e-10, 
    9.825314702601101e-10, 9.7915393174555851e-10, 9.750989045780606e-10, 
    9.7044843169804084e-10, 9.6530710857124918e-10, 9.5978613175036937e-10, 
    9.539889717380112e-10, 9.4799979103204112e-10, 9.418751565842621e-10, 
    9.3563950724165641e-10, 9.2928432858764708e-10, 9.2277085825884459e-10, 
    9.1603569677528823e-10, 9.0899875055202165e-10, 9.0157249651076316e-10, 
    8.9367184323988107e-10, 8.852235922178734e-10, 8.7617481199456149e-10, 
    8.6649936279422283e-10, 8.5620224467079088e-10, 8.4532138240713971e-10, 
    8.3392685130084187e-10, 8.221175994839487e-10, 8.1001604712976986e-10, 
    7.9776087594910726e-10, 7.8549867562595582e-10, 7.733749239873502e-10, 
    7.6152504220641421e-10, 7.5006607262591292e-10, 7.3908965842865091e-10, 
    7.2865672705360577e-10, 7.1879440699279487e-10, 7.0949527930991325e-10, 
    7.0071923212402964e-10, 6.9239761883961517e-10, 6.8443961750849377e-10, 
    6.7674017275270158e-10, 6.691890524604372e-10, 6.6168015942291209e-10, 
    6.5412050009558927e-10, 6.4643793618819842e-10, 6.3858717691447561e-10, 
    6.3055340721467127e-10, 6.2235332583025726e-10, 6.1403340059338137e-10, 
    6.0566557239035391e-10, 5.9734063956902958e-10, 5.8916000005654871e-10, 
    5.8122631034815853e-10, 5.7363395866983027e-10, 5.6646007268150533e-10, 
    5.5975690254941127e-10, 5.5354617036920846e-10, 5.4781599856671225e-10, 
    5.4252062803613087e-10, 5.3758311212077106e-10, 5.329007262807282e-10, 
    5.2835280302920872e-10, 5.2381027626996301e-10, 5.1914627595403193e-10, 
    5.1424677997570373e-10, 5.0902052810271129e-10, 5.0340725564744005e-10, 
    4.9738360738942258e-10, 4.9096614921751239e-10, 4.8421129956822426e-10, 
    4.7721208831892793e-10, 4.7009217656160103e-10, 4.629975231183619e-10, 
    4.5608655747662733e-10, 4.4951952447858015e-10, 4.4344802103105388e-10, 
    4.380053400379604e-10, 4.3329844077471614e-10, 4.2940191005271215e-10, 
    4.2635432199406248e-10, 4.2415695821735414e-10, 4.2277492472145272e-10, 
    4.2214026971602933e-10, 4.2215686644743363e-10, 4.2270647847017176e-10, 
    4.2365568088195925e-10, 4.2486299863720908e-10, 4.2618601093979331e-10, 
    4.2748786404958539e-10, 4.2864302812457469e-10, 4.2954193276221038e-10, 
    4.3009443336286405e-10, 4.3023193000757112e-10, 4.2990824148778104e-10, 
    4.2909916260356352e-10, 4.2780101062363185e-10, 4.2602815110578684e-10, 
    4.2380991135490062e-10, 4.2118696824805304e-10, 4.1820761313044057e-10, 
    4.1492400371335484e-10, 4.1138879036738731e-10, 4.07652160794441e-10, 
    4.0375962762685539e-10, 3.9975050701254539e-10, 3.9565730822997196e-10, 
    3.9150586257594578e-10, 3.8731627935977491e-10, 3.8310447899781377e-10, 
    3.7888424537397547e-10, 3.7466941802237883e-10, 3.7047618059027644e-10, 
    3.663249883980102e-10, 3.6224207798456316e-10, 3.5826018140961568e-10, 
    3.5441847951199312e-10, 3.5076157745655961e-10, 3.4733767467429494e-10, 
    3.4419589791566589e-10, 3.4138316727337806e-10, 3.389407036288511e-10, 
    3.369006393366422e-10, 3.3528291115826063e-10, 3.3409287090999033e-10, 
    3.3331972156181852e-10, 3.3293608430274643e-10, 3.3289862087332955e-10, 
    3.3314983360962067e-10, 3.3362076182790098e-10, 3.3423451631385434e-10, 
    3.3491023761416303e-10, 3.3556730167441454e-10, 3.3612934512400976e-10, 
    3.3652797017688759e-10, 3.3670573350170081e-10, 3.3661844648268198e-10, 
    3.3623652894971758e-10, 3.3554556040534545e-10, 3.345459601320663e-10, 
    3.3325202980337819e-10, 3.3169034137108499e-10, 3.2989777202738226e-10, 
    3.2791918794525978e-10, 3.2580499737780509e-10, 3.2360855758633979e-10, 
    3.2138363844397066e-10, 3.1918187347821257e-10, 3.1705038450175031e-10, 
    3.1502954036782376e-10, 3.13151036644156e-10, 3.1143627513537593e-10, 
    3.0989526268241082e-10, 3.0852600713528843e-10, 3.0731459244086603e-10, 
    3.0623585207185623e-10, 3.0525477563230583e-10, 3.0432846883770643e-10, 
    3.0340866784784299e-10, 3.0244457864736404e-10, 3.0138593565879918e-10, 
    3.0018601152399982e-10, 2.9880445379164183e-10, 2.9720966758713171e-10, 
    2.9538070429244475e-10, 2.9330841196576737e-10, 2.9099590449512994e-10, 
    2.8845823453431479e-10, 2.85721393478444e-10, 2.828206504901189e-10, 
    2.7979843908410518e-10, 2.7670186920306901e-10, 2.7358013928991606e-10, 
    2.7048191809093058e-10, 2.6745296732607047e-10, 2.6453408600488322e-10, 
    2.6175952130669113e-10, 2.5915586551146211e-10, 2.5674152599393558e-10, 
    2.5452667053740275e-10, 2.5251366347472225e-10, 2.5069780668835842e-10, 
    2.4906839207636247e-10, 2.4760985827803784e-10, 2.4630305266297125e-10, 
    2.4512641274562457e-10, 2.4405713906664642e-10, 2.4307220725818748e-10, 
    2.4214931766042935e-10, 2.4126768068591351e-10, 2.4040875583180097e-10, 
    2.3955681637441107e-10, 2.3869947167440002e-10, 2.3782798377533947e-10, 
    2.369374923159015e-10, 2.3602699061169592e-10, 2.3509912655187244e-10, 
    2.3415972812757709e-10, 2.3321714232795386e-10, 2.3228134194338239e-10, 
    2.3136292771667342e-10, 2.3047204424782631e-10, 2.2961738228555857e-10, 
    2.2880525309713101e-10, 2.2803896486533622e-10, 2.2731843545200722e-10, 
    2.2664018153864996e-10, 2.259976009576118e-10, 2.2538160223604866e-10, 
    2.2478140282939414e-10, 2.2418552331417047e-10, 2.2358278744120633e-10, 
    2.2296327964567825e-10, 2.2231912970749437e-10, 2.2164509938952331e-10, 
    2.2093886253697778e-10, 2.2020104398878726e-10, 2.194349398205055e-10, 
    2.1864603007002026e-10, 2.1784125477595725e-10, 2.1702820490214773e-10, 
    2.162142017261325e-10, 2.1540542605454645e-10, 2.1460608036019844e-10, 
    2.1381772868123439e-10, 2.1303875703011847e-10, 2.1226411581121269e-10, 
    2.1148526779261059e-10, 2.106904453979047e-10, 2.098650912267123e-10, 
    2.0899264390570495e-10, 2.0805543866373135e-10, 2.0703584640206337e-10, 
    2.0591746094637401e-10, 2.0468635340524599e-10, 2.0333220385115951e-10, 
    2.0184935780141804e-10, 2.0023756035390122e-10, 1.9850245193809854e-10, 
    1.9665563474212475e-10, 1.9471438447258216e-10, 1.9270092338288804e-10, 
    1.9064135960077698e-10, 1.8856429285710717e-10, 1.8649924374897649e-10, 
    1.8447496098293146e-10, 1.8251780624962731e-10, 1.8065022785360353e-10, 
    1.7888957690636245e-10, 1.7724722727005657e-10, 1.7572813761938442e-10, 
    1.7433083101653526e-10, 1.7304782394922434e-10, 1.718663940132215e-10, 
    1.7076969677174183e-10, 1.6973804990313369e-10, 1.6875037430669606e-10, 
    1.6778561078899724e-10, 1.6682407540070821e-10, 1.6584862518700031e-10, 
    1.6484561207891288e-10, 1.6380551033762414e-10, 1.6272326695677897e-10, 
    1.6159828266824948e-10, 1.6043410686970911e-10, 1.592378085354333e-10, 
    1.5801915028944505e-10, 1.5678954058080784e-10, 1.5556093750351727e-10, 
    1.5434474049169836e-10, 1.531507820519599e-10, 1.5198650705513178e-10, 
    1.5085642232361428e-10, 1.4976183780732223e-10, 1.4870096542040942e-10, 
    1.4766929936006392e-10, 1.4666030434049681e-10, 1.4566625488768797e-10, 
    1.4467920227032286e-10, 1.4369191340621794e-10, 1.4269872528413937e-10, 
    1.4169619406619751e-10, 1.4068352555675566e-10, 1.396627210913316e-10, 
    1.3863849058923954e-10, 1.3761792860858563e-10, 1.3661003308192481e-10, 
    1.3562511917737969e-10, 1.3467419158829316e-10, 1.337683421098612e-10, 
    1.3291820622255874e-10, 1.3213347576924176e-10, 1.3142253696414312e-10, 
    1.3079215112743007e-10, 1.3024723824683947e-10, 1.2979069021866188e-10, 
    1.2942325690394729e-10, 1.2914346414119538e-10, 1.2894759719895868e-10, 
    1.2882974383511056e-10, 1.2878191791537198e-10, 1.2879427678432484e-10, 
    1.2885541332985012e-10, 1.2895272746805134e-10, 1.2907284699835755e-10, 
    1.2920207105981071e-10, 1.2932679321688152e-10, 1.2943387042762956e-10, 
    1.2951092442430839e-10, 1.2954654754315986e-10, 1.295304343363338e-10, 
    1.2945343052940945e-10, 1.293075699992438e-10, 1.2908609535725508e-10, 
    1.2878353000718213e-10, 1.2839580198120934e-10, 1.2792044850376321e-10, 
    1.2735686941593134e-10, 1.2670661009829001e-10, 1.2597362540753581e-10, 
    1.2516447057351543e-10, 1.2428834695970997e-10, 1.2335697529699656e-10, 
    1.2238427278072111e-10, 1.2138583147486158e-10, 1.2037821524543895e-10, 
    1.1937817546280954e-10, 1.1840180758594266e-10, 1.1746379052067621e-10, 
    1.1657672898268816e-10, 1.1575072703021198e-10, 1.1499315674215578e-10, 
    1.1430870279162865e-10, 1.1369955900061761e-10, 1.1316580442932719e-10, 
    1.1270583419775608e-10, 1.1231676300994754e-10, 1.1199473735032424e-10, 
    1.1173511740463715e-10, 1.1153246303774394e-10, 1.1138040635957351e-10, 
    1.1127136900887693e-10, 1.1119627921119255e-10, 1.1114430127871162e-10, 
    1.11102726592193e-10, 1.1105700292575913e-10, 1.1099105629673954e-10, 
    1.1088781446369385e-10, 1.1072998707550534e-10, 1.1050097115841837e-10, 
    1.101858683166076e-10, 1.0977246134347688e-10, 1.0925211142494683e-10, 
    1.0862041025761081e-10, 1.0787762289360534e-10, 1.0702877094344149e-10, 
    1.0608347133551198e-10, 1.0505544023706763e-10, 1.0396181073240855e-10, 
    1.0282225336647123e-10, 1.016580443765738e-10, 1.0049108547362161e-10, 
    9.9343015739442423e-11, 9.8234390328866998e-11, 9.7184037805948287e-11, 
    9.6208522132185591e-11, 9.532179087614995e-11, 9.4534908139654478e-11, 
    9.3855932834293852e-11, 9.3289835570984718e-11, 9.2838511136068742e-11, 
    9.2500797502443532e-11, 9.2272585763140504e-11, 9.214692589217089e-11, 
    9.2114251731855592e-11, 9.2162635578338884e-11, 9.2278180033400015e-11, 
    9.2445470069181441e-11, 9.264815268245247e-11, 9.2869551263202141e-11, 
    9.309336352280571e-11, 9.330431029138644e-11, 9.3488787643633767e-11, 
    9.3635351148763222e-11, 9.3735117835983969e-11, 9.378193981994357e-11, 
    9.3772430434582945e-11, 9.3705744244103407e-11, 9.358324952070382e-11, 
    9.3408009099010971e-11, 9.3184225735011494e-11, 9.2916625140299148e-11, 
    9.2609908704425526e-11, 9.2268226259416137e-11, 9.189483149037333e-11, 
    9.1491822848930025e-11, 9.1060089681028978e-11, 9.059935675878811e-11, 
    9.010840849890508e-11, 8.958537824399705e-11, 8.9028156328780703e-11, 
    8.8434769716791698e-11, 8.7803821418450805e-11, 8.713484612278574e-11, 
    8.6428640438574569e-11, 8.5687446415377213e-11, 8.49150805188142e-11, 
    8.4116901761486772e-11, 8.3299698684299178e-11, 8.2471418736590149e-11, 
    8.1640885984545161e-11, 8.0817342986844141e-11, 8.001007391375362e-11, 
    7.9227936179414135e-11, 7.8478993127304715e-11, 7.7770154811192444e-11, 
    7.710696251132672e-11, 7.6493439953997831e-11, 7.5932106019165817e-11, 
    7.5424065641425274e-11, 7.4969250948058797e-11, 7.456670769913949e-11, 
    7.4214990507251547e-11, 7.3912530571458508e-11, 7.3658044888408627e-11, 
    7.3450839072754673e-11, 7.3291069935394942e-11, 7.3179828829356179e-11, 
    7.3119127402317381e-11, 7.3111658195754509e-11, 7.3160453233328825e-11, 
    7.3268326498887671e-11, 7.3437250000652745e-11, 7.3667646955633581e-11, 
    7.3957710816631751e-11, 7.4302757094300218e-11, 7.4694785021365331e-11, 
    7.5122196650717962e-11, 7.5569830593025371e-11, 7.601924864533265e-11, 
    7.6449356521658527e-11, 7.6837238908393914e-11, 7.7159244742857457e-11, 
    7.7392181900262643e-11, 7.75145620265759e-11, 7.7507791054140144e-11, 
    7.7357225486010588e-11, 7.7052998134356058e-11, 7.6590587902513179e-11, 
    7.5971074344481315e-11, 7.5201100127862824e-11, 7.4292507817905878e-11, 
    7.3261758394229273e-11, 7.212911593354137e-11, 7.0917723271718992e-11, 
    6.9652571134821849e-11, 6.8359480459859604e-11, 6.7064116644469983e-11, 
    6.5791112611890388e-11, 6.4563300416343822e-11, 6.3401120523825586e-11, 
    6.23221689848756e-11, 6.1340934038106635e-11, 6.0468661345848293e-11, 
    5.9713376218827016e-11, 5.9079981870897521e-11, 5.8570478990715321e-11, 
    5.818419412854855e-11, 5.7918064065267878e-11, 5.7766914722095982e-11, 
    5.772372821391857e-11, 5.7779876483655773e-11, 5.792535883781134e-11, 
    5.8148991281729199e-11, 5.8438621370519031e-11, 5.8781314666137955e-11, 
    5.916358872131846e-11, 5.9571639955618423e-11, 5.99916345585754e-11, 
    6.0409991114820556e-11, 6.0813721633776083e-11, 6.1190753132622953e-11, 
    6.1530285723660558e-11, 6.1823099966149009e-11, 6.2061883440289381e-11, 
    6.22414680036267e-11, 6.2359056756397387e-11, 6.2414348666391626e-11, 
    6.2409604908485512e-11, 6.2349590882949109e-11, 6.224143326856607e-11, 
    6.2094336343962854e-11, 6.1919187273636769e-11, 6.1728039532720265e-11, 
    6.153351500444196e-11, 6.1348104351555642e-11, 6.1183479540416676e-11, 
    6.1049793940132877e-11, 6.0955077718911469e-11, 6.0904729899732482e-11, 
    6.090119484795795e-11, 6.0943792489158066e-11, 6.1028776124815557e-11, 
    6.114955486802443e-11, 6.1297081379935028e-11, 6.1460369636035251e-11, 
    6.1627086357398631e-11, 6.1784177552949165e-11, 6.1918484143868327e-11, 
    6.201730930988361e-11, 6.2068937522149889e-11, 6.2063036363303048e-11, 
    6.1991012794606408e-11, 6.1846268285435643e-11, 6.1624390728248691e-11, 
    6.1323269818723293e-11, 6.0943166236567985e-11, 6.0486701453630014e-11, 
    5.9958811851676142e-11, 5.9366601012440738e-11, 5.871916569137814e-11, 
    5.8027298674518352e-11, 5.7303174033979354e-11, 5.6559931087323016e-11, 
    5.5811235350396888e-11, 5.5070784002643776e-11, 5.4351818391138616e-11, 
    5.3666625795050337e-11, 5.3026083845809105e-11, 5.2439236467345854e-11, 
    5.1912949404218603e-11, 5.1451639015563439e-11, 5.1057104676044703e-11, 
    5.0728456319915471e-11, 5.0462189672891495e-11, 5.0252340996430439e-11, 
    5.0090803388641566e-11, 4.9967746756830822e-11, 4.9872138943646187e-11, 
    4.9792341450098799e-11, 4.9716774570305654e-11, 4.963456738655628e-11, 
    4.9536210388083243e-11, 4.9414112533619799e-11, 4.9263062041657924e-11, 
    4.9080535980852164e-11, 4.8866855091773539e-11, 4.8625105623510886e-11, 
    4.8360920234443849e-11, 4.8082039009025198e-11, 4.779773115356393e-11, 
    4.7518084354217512e-11, 4.725322919404306e-11, 4.7012541742631704e-11, 
    4.6803900952235766e-11, 4.663305267624628e-11, 4.6503154503148369e-11, 
    4.6414510179626733e-11, 4.6364587505076534e-11, 4.6348247493412954e-11, 
    4.6358242501455268e-11, 4.638588585218553e-11, 4.6421870122410879e-11, 
    4.6457124852454264e-11, 4.6483656033135829e-11, 4.6495251308500001e-11, 
    4.6488004219895249e-11, 4.6460599648500925e-11, 4.6414308652744193e-11, 
    4.6352729723129821e-11, 4.6281290159200417e-11, 4.6206552866648464e-11, 
    4.6135437746030244e-11, 4.6074410957397364e-11, 4.6028761999091256e-11, 
    4.6001985099236682e-11, 4.5995383610477865e-11, 4.6007896864629417e-11, 
    4.6036153930045704e-11, 4.607473216162598e-11, 4.6116584279635906e-11, 
    4.6153587149926596e-11, 4.617714086015839e-11, 4.6178729030910478e-11, 
    4.6150446792529509e-11, 4.6085405054387089e-11, 4.5978012923896762e-11, 
    4.5824123820012768e-11, 4.5621060312184055e-11, 4.5367544557612349e-11, 
    4.506355618628074e-11, 4.4710158986364465e-11, 4.4309318720939868e-11, 
    4.3863761187674916e-11, 4.3376847847244569e-11, 4.2852503054174259e-11, 
    4.2295191737950922e-11, 4.1709879486850461e-11, 4.1102034739557264e-11, 
    4.0477589711026415e-11, 3.9842866310216248e-11, 3.9204455800524185e-11, 
    3.8569052282906592e-11, 3.7943234631759464e-11, 3.7333232485892212e-11, 
    3.6744705430255103e-11, 3.6182551528416317e-11, 3.5650773163100301e-11, 
    3.5152436061208108e-11, 3.4689718981222636e-11, 3.4264054175594657e-11, 
    3.3876342693964627e-11, 3.3527216272534481e-11, 3.3217299596810115e-11, 
    3.2947437648936839e-11, 3.2718847006623227e-11, 3.2533145329647536e-11, 
    3.2392258192598804e-11, 3.2298178403841294e-11, 3.2252622141562882e-11, 
    3.2256587821232041e-11, 3.2309883163173492e-11, 3.2410671450256212e-11, 
    3.255512411805539e-11, 3.2737196264955778e-11, 3.2948596378226982e-11, 
    3.3178972665147941e-11, 3.3416325344931987e-11, 3.3647594972696347e-11, 
    3.3859416784863828e-11, 3.4038963190049265e-11, 3.4174773046450339e-11, 
    3.4257542450297877e-11, 3.4280762674381074e-11, 3.4241153115093629e-11, 
    3.4138871651001177e-11, 3.397746556823333e-11, 3.3763590877881239e-11, 
    3.3506538661136455e-11, 3.3217581640300151e-11, 3.2909272514681257e-11, 
    3.259467921669076e-11, 3.2286680573132181e-11, 3.1997317202132738e-11, 
    3.173726643833768e-11, 3.1515439392304851e-11, 3.133869954154242e-11, 
    3.1211694227642577e-11, 3.1136778167657874e-11, 3.1114024846099771e-11, 
    3.1141275299075249e-11, 3.1214241136819874e-11, 3.1326647899543574e-11, 
    3.1470405944451608e-11, 3.163584835709603e-11, 3.1812009632752334e-11, 
    3.1986991274690576e-11, 3.2148374796476345e-11, 3.2283723239984859e-11, 
    3.2381119095723953e-11, 3.2429747560082313e-11, 3.2420454757709164e-11, 
    3.2346283127581232e-11, 3.2202897009447212e-11, 3.1988904320598072e-11, 
    3.170599161358341e-11, 3.1358901376464516e-11, 3.095518556352924e-11, 
    3.0504804401356349e-11, 3.0019530734923017e-11, 2.9512264774146611e-11, 
    2.8996259159191005e-11, 2.8484347342364957e-11, 2.7988213077864476e-11, 
    2.7517787644575521e-11, 2.7080786918463799e-11, 2.668245563961971e-11, 
    2.6325502235095757e-11, 2.6010251412312611e-11, 2.5734939907013903e-11, 
    2.5496185253947647e-11, 2.5289499275787505e-11, 2.5109867860477135e-11, 
    2.4952270636877228e-11, 2.4812174267599966e-11, 2.4685873647757735e-11, 
    2.4570761272340708e-11, 2.4465425633203123e-11, 2.4369665584913757e-11, 
    2.4284365950048262e-11, 2.4211333260417673e-11, 2.4153025801705182e-11, 
    2.41123056087804e-11, 2.4092128969648571e-11, 2.409531142076774e-11, 
    2.4124234589737669e-11, 2.418067852296957e-11, 2.4265617490778572e-11, 
    2.4379150303433612e-11, 2.4520426561747647e-11, 2.4687700269182447e-11, 
    2.4878410054413723e-11, 2.5089372060279252e-11, 2.5316979888464118e-11, 
    2.5557524610010853e-11, 2.5807428523991186e-11, 2.6063582580626314e-11, 
    2.6323538776751737e-11, 2.6585717043392442e-11, 2.684944797999594e-11, 
    2.7114991385412744e-11, 2.7383352319638932e-11, 2.7656124630837445e-11, 
    2.7935151723724434e-11, 2.8222265927879486e-11, 2.8518929477224798e-11, 
    2.882599803904115e-11, 2.9143477534097564e-11, 2.9470427499335322e-11, 
    2.9804865511372451e-11, 3.0143838029637582e-11, 3.0483477186207408e-11, 
    3.0819154617623348e-11, 3.1145619126342075e-11, 3.145717681610423e-11, 
    3.1747815931123029e-11, 3.2011391006427952e-11, 3.2241711554597926e-11, 
    3.2432721677474271e-11, 3.257861990150461e-11, 3.2674054030422749e-11, 
    3.2714289388952638e-11, 3.2695476395389561e-11, 3.2614836965413832e-11, 
    3.2470958612241158e-11, 3.2263988411102239e-11, 3.1995848858806842e-11, 
    3.167033477198122e-11, 3.1293167624243832e-11, 3.0871903846810144e-11, 
    3.0415766121943821e-11, 2.9935317846096727e-11, 2.944207616506298e-11, 
    2.8947982932740568e-11, 2.8464866321394102e-11, 2.8003835282061798e-11, 
    2.7574730412954833e-11, 2.7185588028423426e-11, 2.6842242659892226e-11, 
    2.6548022981811737e-11, 2.6303640305131425e-11, 2.6107208666031937e-11, 
    2.5954477899975929e-11, 2.5839164472572168e-11, 2.5753456762516644e-11, 
    2.568856304459178e-11, 2.5635321043342673e-11, 2.5584773024088539e-11, 
    2.5528712017750392e-11, 2.5460072282418097e-11, 2.5373261369368614e-11, 
    2.5264315877495174e-11, 2.5130959952739779e-11, 2.4972531604240661e-11, 
    2.4789855005148236e-11, 2.4585050563857233e-11, 2.4361356693548629e-11, 
    2.4122926847079333e-11, 2.3874685629850313e-11, 2.3622182895296042e-11, 
    2.3371480123802339e-11, 2.3128991122655964e-11, 2.2901318199331908e-11, 
    2.2695005159797399e-11, 2.2516244404148078e-11, 2.2370472082598925e-11, 
    2.2261958915655969e-11, 2.2193360027922487e-11, 2.2165325479164544e-11, 
    2.2176181710699954e-11, 2.2221798365821184e-11, 2.2295624065295111e-11, 
    2.2388972442390377e-11, 2.249151550085389e-11, 2.2592010173243567e-11, 
    2.2679135723224887e-11, 2.2742444435928147e-11, 2.277327300761722e-11, 
    2.2765579204333593e-11, 2.2716546860251762e-11, 2.2626975137701896e-11, 
    2.2501325056211394e-11, 2.2347474458211222e-11, 2.2176151827567312e-11, 
    2.2000119161336573e-11, 2.1833175338341309e-11, 2.1689065158331373e-11, 
    2.1580374080654243e-11, 2.151754164560457e-11, 2.1508021605750114e-11, 
    2.1555720482214304e-11, 2.1660676887088065e-11, 2.1819082039562034e-11, 
    2.2023538994824831e-11, 2.2263607769066202e-11, 2.2526518067811519e-11, 
    2.2798032764147559e-11, 2.3063330642817404e-11, 2.3307909575173673e-11, 
    2.3518364051617365e-11, 2.3683079131232055e-11, 2.3792691000962595e-11, 
    2.3840406692162086e-11, 2.382211250231573e-11, 2.3736335148010788e-11, 
    2.3584001058046708e-11, 2.3368156025164218e-11, 2.309357916520159e-11, 
    2.276640168593687e-11, 2.2393714199660551e-11, 2.1983247861218731e-11, 
    2.1543096253845181e-11, 2.1081525639834102e-11, 2.060684071590696e-11, 
    2.0127316987104059e-11, 1.9651147368775071e-11, 1.9186424552106748e-11, 
    1.8741093202908124e-11, 1.8322892576285776e-11, 1.7939251204103413e-11, 
    1.7597149014369948e-11, 1.7302938581383474e-11, 1.7062159264935526e-11, 
    1.6879325808122154e-11, 1.6757749978399004e-11, 1.6699372526488137e-11, 
    1.6704654682446487e-11, 1.6772506155743824e-11, 1.6900290802842197e-11, 
    1.7083864208956746e-11, 1.7317696075729767e-11, 1.7595024615945289e-11, 
    1.7908074986211574e-11, 1.8248321430811184e-11, 1.860679922586791e-11, 
    1.8974428926287029e-11, 1.9342403986311469e-11, 1.9702550248384485e-11, 
    2.0047709195909466e-11, 2.0372070529752542e-11, 2.0671460268789119e-11, 
    2.0943523656164829e-11, 2.1187825050233585e-11, 2.1405793101879453e-11, 
    2.1600566026778026e-11, 2.1776662910143717e-11, 2.1939581215889821e-11, 
    2.2095290716782999e-11, 2.2249693353446832e-11, 2.2408063913777757e-11, 
    2.2574551683411671e-11, 2.2751766112208799e-11, 2.2940482848069337e-11, 
    2.3139481207426332e-11, 2.3345556148553672e-11, 2.3553655455072479e-11, 
    2.3757159143261445e-11, 2.3948260268507437e-11, 2.4118424496189478e-11, 
    2.4258853234367748e-11, 2.4360979799403823e-11, 2.4416922135494593e-11, 
    2.4419883512990657e-11, 2.4364488675814199e-11, 2.4247056364216671e-11, 
    2.4065784577205068e-11, 2.3820886864011633e-11, 2.3514632195727819e-11, 
    2.3151354731872234e-11, 2.2737357881834975e-11, 2.2280786843468814e-11, 
    2.1791381500950113e-11, 2.1280185374062886e-11, 2.0759149730717525e-11, 
    2.0240683899376807e-11, 1.9737108589878252e-11, 1.9260107154751883e-11, 
    1.8820156547368684e-11, 1.8426004900023719e-11, 1.8084221161334274e-11, 
    1.7798898604745758e-11, 1.7571493332614028e-11, 1.7400870045768356e-11, 
    1.7283542965929762e-11, 1.7214103054034172e-11, 1.7185770849914998e-11, 
    1.7191068628162983e-11, 1.7222510634195612e-11, 1.7273269927145127e-11, 
    1.7337707632920673e-11, 1.7411759498499842e-11, 1.7493113785489226e-11, 
    1.7581174499884949e-11, 1.7676800404768139e-11, 1.7781889958767158e-11, 
    1.7898846985882642e-11, 1.8030000922993645e-11, 1.8177042083136509e-11, 
    1.8340568373000624e-11, 1.8519754483952407e-11, 1.8712213096619691e-11, 
    1.8914034298418894e-11, 1.9120003394872488e-11, 1.932394374363706e-11, 
    1.9519167800416384e-11, 1.9698949516365014e-11, 1.9856997731757847e-11, 
    1.9987857202583105e-11, 2.008721096900386e-11, 2.0152070933280681e-11, 
    2.0180848664834378e-11, 2.0173284851439719e-11, 2.0130304116158079e-11, 
    2.0053798985245292e-11, 1.9946371307872163e-11, 1.9811053003698083e-11, 
    1.9651075922604609e-11, 1.9469673134179998e-11, 1.9269951003877318e-11, 
    1.9054814046487875e-11, 1.8826972125697013e-11, 1.8588975736975035e-11, 
    1.8343304610680278e-11, 1.8092425795696264e-11, 1.783885131922599e-11, 
    1.7585143629621976e-11, 1.7333867267088784e-11, 1.7087452030478712e-11, 
    1.6848031966659432e-11, 1.6617213330419939e-11, 1.6395863403146834e-11, 
    1.6183898132814165e-11, 1.5980144948511021e-11, 1.5782286684610189e-11, 
    1.5586921555938016e-11, 1.538973578686847e-11, 1.5185795972863107e-11, 
    1.4969907124848191e-11, 1.4737050194567603e-11, 1.448280317771896e-11, 
    1.4203753461785206e-11, 1.3897799659562285e-11, 1.3564378622349283e-11, 
    1.3204535707244155e-11, 1.2820884734289919e-11, 1.2417443367507278e-11, 
    1.1999396068270474e-11, 1.1572767833703644e-11, 1.1144116186045501e-11, 
    1.0720233071893942e-11, 1.0307891260106218e-11, 9.9136438852709356e-12, 
    9.5437126766886507e-12, 9.2038916542612084e-12, 8.899517178291075e-12, 
    8.63541439935987e-12, 8.4158488290762641e-12, 8.2444134990725758e-12, 
    8.1238963548292004e-12, 8.0560798704303737e-12, 8.0415394212748145e-12, 
    8.0794284932652465e-12, 8.1673350553194472e-12, 8.3011796755092296e-12, 
    8.4752805793715572e-12, 8.6825208974093533e-12, 8.9146951209535552e-12, 
    9.1629793871343525e-12, 9.4185331556692613e-12, 9.6731363494438455e-12, 
    9.9198566074294755e-12, 1.015363837869539e-11, 1.0371769615751263e-11, 
    1.057414802867401e-11, 1.0763334087064951e-11, 1.0944351320541815e-11, 
    1.1124262069962425e-11, 1.1311513920757597e-11, 1.1515164671716698e-11, 
    1.1744011526617915e-11, 1.2005727908821742e-11, 1.2306079399797157e-11, 
    1.2648272919976502e-11, 1.3032538429633339e-11, 1.3455915211638238e-11, 
    1.3912294981791427e-11, 1.4392697487728455e-11, 1.4885750236124666e-11, 
    1.5378318007925803e-11, 1.5856238201362386e-11, 1.6305103701729981e-11, 
    1.6711031071352487e-11, 1.7061376619063098e-11, 1.7345345497324696e-11, 
    1.7554478727948097e-11, 1.7683010111228049e-11, 1.7728039743980226e-11, 
    1.7689582258501402e-11, 1.7570462629052793e-11, 1.7376072484018412e-11, 
    1.7114029830415589e-11, 1.6793747400623975e-11, 1.6425949129998111e-11, 
    1.602213714015617e-11, 1.5594087922076031e-11, 1.5153358681994011e-11, 
    1.4710849855876373e-11, 1.4276471868870569e-11, 1.3858883068438765e-11, 
    1.3465344447292916e-11, 1.3101687412409903e-11, 1.2772363814769923e-11, 
    1.2480585063172932e-11, 1.2228514504102179e-11, 1.2017488008574858e-11, 
    1.1848224886243865e-11, 1.1721010909464214e-11, 1.1635829726491207e-11, 
    1.1592423367856768e-11, 1.1590283709619107e-11, 1.1628585029824239e-11, 
    1.1706061912891812e-11, 1.182087358313676e-11, 1.1970475999522185e-11, 
    1.2151545625828574e-11, 1.2359930820331415e-11, 1.2590731759077811e-11, 
    1.2838437994810982e-11, 1.3097157333703575e-11, 1.3360917189296953e-11, 
    1.3623991355107264e-11, 1.3881234267941404e-11, 1.4128386278225701e-11, 
    1.4362294335830964e-11, 1.4581051188840896e-11, 1.4784016107949785e-11, 
    1.4971723916607965e-11, 1.5145683402389537e-11, 1.5308099813028284e-11, 
    1.546155416367919e-11, 1.5608671320454154e-11, 1.5751803508007639e-11, 
    1.5892792564636425e-11, 1.6032809210804185e-11, 1.617227173374209e-11, 
    1.6310890994676793e-11, 1.6447772395439765e-11, 1.6581554485987627e-11, 
    1.671059509131022e-11, 1.6833136116763189e-11, 1.6947422582652331e-11, 
    1.7051777904798918e-11, 1.7144604685034368e-11, 1.7224335175861756e-11, 
    1.7289345559741872e-11, 1.7337861333866533e-11, 1.7367885946097e-11, 
    1.7377191835425897e-11, 1.7363384624065777e-11, 1.7324053857721412e-11, 
    1.7257015571311101e-11, 1.7160590981664082e-11, 1.7033938321727899e-11, 
    1.6877324589627256e-11, 1.6692349265419403e-11, 1.6482046408851281e-11, 
    1.6250848584434701e-11, 1.6004375870219293e-11, 1.5749099647520076e-11, 
    1.5491895409910042e-11, 1.523951109231386e-11, 1.4998061956189645e-11, 
    1.4772569927414732e-11, 1.4566608530952295e-11, 1.4382125311760437e-11, 
    1.4219427843019429e-11, 1.4077355643334393e-11, 1.3953584410077094e-11, 
    1.3845048114032864e-11, 1.3748387890429738e-11, 1.3660388424492861e-11, 
    1.3578341350185447e-11, 1.3500289705966411e-11, 1.342511126437225e-11, 
    1.3352473378398859e-11, 1.3282652603193851e-11, 1.3216265915280576e-11, 
    1.3153939441062076e-11, 1.3096003016880459e-11, 1.3042223597625048e-11, 
    1.2991636680361692e-11, 1.2942473562441127e-11, 1.2892224386377783e-11, 
    1.2837784529176819e-11, 1.2775708052503209e-11, 1.270249306984836e-11, 
    1.2614896065674581e-11, 1.2510221041445058e-11, 1.2386572506155396e-11, 
    1.2243030507323318e-11, 1.2079767904607921e-11, 1.1898067321335712e-11, 
    1.1700288052570681e-11, 1.1489742590034499e-11, 1.1270535790913911e-11, 
    1.1047362252450302e-11, 1.0825275789314106e-11, 1.0609434747666555e-11, 
    1.0404863326127977e-11, 1.0216193182869465e-11, 1.0047451461782762e-11, 
    9.9018484536871561e-12, 9.7816058589026868e-12, 9.6878437210766656e-12, 
    9.6204979302409958e-12, 9.5782893853378315e-12, 9.5587629543867024e-12, 
    9.5583656229719742e-12, 9.5725937130486048e-12, 9.5961576278172354e-12, 
    9.6232044867790638e-12, 9.6475453207463588e-12, 9.6628920791395561e-12, 
    9.6631077655091061e-12, 9.6424195244590919e-12, 9.5956329889257921e-12, 
    9.518318670298489e-12, 9.4069734848495302e-12, 9.2591685918131483e-12, 
    9.073691674934278e-12, 8.8506542006615006e-12, 8.5916100052649707e-12, 
    8.2996239500509451e-12, 7.9793205564008462e-12, 7.6368693379082879e-12, 
    7.2798993805518333e-12, 6.9173226763514485e-12, 6.55904952763121e-12, 
    6.2156125706374699e-12, 5.8977002226461557e-12, 5.615621096803655e-12, 
    5.3787606956222674e-12, 5.195054007224211e-12, 5.070544488064153e-12, 
    5.0090524827675844e-12, 5.0120287178744478e-12, 5.0785630004215772e-12, 
    5.2055734036004776e-12, 5.3881502145408767e-12, 5.6200124225969973e-12, 
    5.8940113044933063e-12, 6.2026485174449806e-12, 6.5385160641655524e-12, 
    6.8946579651188547e-12, 7.2647866243537917e-12, 7.6433664911525315e-12, 
    8.0255619839754718e-12, 8.4071241356492102e-12, 8.7841806941920909e-12, 
    9.1530344505312414e-12, 9.5099755482182611e-12, 9.8511810962133177e-12, 
    1.017266636032603e-11, 1.0470336865073502e-11, 1.0740100777817924e-11, 
    1.0978051233924276e-11, 1.1180657709138902e-11, 1.1344962974210869e-11, 
    1.1468732265205926e-11, 1.1550572619091491e-11, 1.1589963127107832e-11, 
    1.1587242382294937e-11, 1.1543525353742088e-11, 1.146059079176274e-11, 
    1.1340735855030943e-11, 1.1186639209017276e-11, 1.1001238052361093e-11, 
    1.0787628286398239e-11, 1.0549013514055827e-11, 1.0288677275422157e-11, 
    1.0009989055863004e-11, 9.7164358102676174e-12, 9.4116447233935958e-12, 
    9.0994071899746549e-12, 8.7836793079022668e-12, 8.4685481903295862e-12, 
    8.1581699209891015e-12, 7.8566905975983603e-12, 7.5681332620682091e-12, 
    7.2962949536609385e-12, 7.0446448291732184e-12, 6.8162402590597043e-12, 
    6.6136920478254696e-12, 6.4391488200673554e-12, 6.2943335927063099e-12, 
    6.1805954102602557e-12, 6.0989849637005537e-12, 6.0503357348387813e-12, 
    6.0353070684740066e-12, 6.0544254330062293e-12, 6.1080535918941943e-12, 
    6.1963297138364185e-12, 6.3190465419338713e-12, 6.4755033409234105e-12, 
    6.664332643068882e-12, 6.8833249927307391e-12, 7.1292728112667638e-12, 
    7.3978900575716932e-12, 7.6837921850946783e-12, 7.9805515701650716e-12, 
    8.2808804635954408e-12, 8.5768988663857428e-12, 8.8604835074712991e-12, 
    9.1236844744640111e-12, 9.3591544261587923e-12, 9.5605638027860376e-12, 
    9.7229477784759868e-12, 9.8429611724991044e-12, 9.9189843659243689e-12, 
    9.9510869989952058e-12, 9.9408404640175615e-12, 9.8909907161768134e-12, 
    9.8050355600848825e-12, 9.6867584246696461e-12, 9.5397613842545586e-12, 
    9.3670663148937653e-12, 9.1708313439819048e-12, 8.9522260106477494e-12, 
    8.7114795532811227e-12, 8.4481077602820008e-12, 8.1612957808962112e-12, 
    7.8503945264405882e-12, 7.5154661182461005e-12, 7.1578578834087889e-12, 
    6.7806920400195572e-12, 6.3892198051226023e-12, 5.991030253000539e-12, 
    5.5960440354970774e-12, 5.2162902950398017e-12, 4.8654715924086161e-12, 
    4.5583400309583279e-12, 4.3099164368473947e-12, 4.1346007558143682e-12, 
    4.0452521017262702e-12, 4.0522703178486401e-12, 4.1627651958173694e-12, 
    4.37987513093964e-12, 4.7022813031851688e-12, 5.1239622074820542e-12, 
    5.6342427636065968e-12, 6.218126655753941e-12, 6.8569005709985262e-12, 
    7.5290260076991407e-12, 8.2112264329351706e-12, 8.8797246278405474e-12, 
    9.5115477911454594e-12, 1.0085795685429577e-11, 1.0584799255819054e-11, 
    1.0995060861806747e-11, 1.1307924412299907e-11, 1.1519914196755823e-11, 
    1.1632719170357048e-11, 1.1652856642871001e-11, 1.1590998908245327e-11, 
    1.1461078503077444e-11, 1.1279241836508761e-11, 1.1062702976824822e-11, 
    1.0828639179085904e-11, 1.0593172345799397e-11, 1.0370522423406537e-11, 
    1.0172377369787656e-11, 1.0007492104721624e-11, 9.8815379701463505e-12, 
    9.7971554539322975e-12, 9.754198792770531e-12, 9.7501370301374178e-12, 
    9.7805319748775596e-12, 9.8395802809075536e-12, 9.9206661759838544e-12, 
    1.001689554181365e-11, 1.0121581960523775e-11, 1.0228686733775194e-11, 
    1.0333185314496533e-11, 1.0431344333450449e-11, 1.0520927564094715e-11, 
    1.0601313195588216e-11, 1.0673510129491647e-11, 1.0740064170632655e-11, 
    1.0804868810653487e-11, 1.0872865132272392e-11, 1.094964626970508e-11, 
    1.1040987988782182e-11, 1.1152328603222739e-11, 1.1288244136400089e-11, 
    1.1451954433427204e-11, 1.1644906713197701e-11, 1.1866482376620579e-11, 
    1.2113852144611298e-11, 1.2382006136014744e-11, 1.2663953918741611e-11, 
    1.2951091844245677e-11, 1.3233691420232569e-11, 1.3501498847559498e-11, 
    1.3744352523249723e-11, 1.3952817092686875e-11, 1.4118750930033233e-11, 
    1.4235789739888488e-11, 1.4299698364260811e-11, 1.4308581858077264e-11, 
    1.4262972602406279e-11, 1.4165753486663657e-11, 1.4021956847608877e-11, 
    1.3838467681293351e-11, 1.362361372010181e-11, 1.3386715417795342e-11, 
    1.3137566369041373e-11, 1.2885921031758481e-11, 1.2640961163637404e-11, 
    1.2410814509940476e-11, 1.2202105385547327e-11, 1.2019603043191545e-11, 
    1.1865943505556104e-11, 1.1741482827182469e-11, 1.1644287128579287e-11, 
    1.1570242492183127e-11, 1.1513308577459415e-11, 1.1465879492121384e-11, 
    1.1419260129122193e-11, 1.1364205025506467e-11, 1.1291457810484754e-11, 
    1.1192311156763559e-11, 1.1059106930805429e-11, 1.0885634835837782e-11, 
    1.0667439538215514e-11, 1.0401995997929424e-11, 1.0088746630179889e-11, 
    9.7290499747901159e-12, 9.3260014774792038e-12, 8.884202124103022e-12, 
    8.4094967249016812e-12, 7.9086986715608165e-12, 7.389311465668148e-12, 
    6.8593074140979246e-12, 6.3269304764457165e-12, 5.800540374559568e-12, 
    5.2884824046124785e-12, 4.7989641939544249e-12, 4.3399450100105861e-12, 
    3.9190001284061672e-12, 3.5431595036375083e-12, 3.2187329142238481e-12, 
    2.9511015914860908e-12, 2.7445084826013996e-12, 2.6018567225029801e-12, 
    2.5245295345322162e-12, 2.5122549785157288e-12, 2.563028877452542e-12, 
    2.6731189635294954e-12, 2.8371353519676841e-12, 3.04818966319486e-12, 
    3.2981230148910995e-12, 3.5777969792652888e-12, 3.8774402951442255e-12, 
    4.1870158106784559e-12, 4.4966130898266845e-12, 4.7968278379000665e-12, 
    5.0791112835091844e-12, 5.3361063406056539e-12, 5.5618971197779445e-12, 
    5.7522224710853255e-12, 5.9046133726653346e-12, 6.0184311130905351e-12, 
    6.0948599364593572e-12, 6.1368039754565344e-12, 6.1487082683887761e-12, 
    6.1363262882192257e-12, 6.106416821140027e-12, 6.0664062796849471e-12, 
    6.0240120753091417e-12, 5.9868731675883984e-12, 5.9621658958928014e-12, 
    5.9562753789722109e-12, 5.9744985490026379e-12, 6.0208086591011925e-12, 
    6.0977067440875832e-12, 6.2061494455902887e-12, 6.3455578576347056e-12, 
    6.5139160674806139e-12, 6.7079333030735709e-12, 6.923265647024949e-12, 
    7.1547885183194382e-12, 7.3968979859009789e-12, 7.6438130504051098e-12, 
    7.8899027379592425e-12, 8.1299642593797344e-12, 8.3595008074701826e-12, 
    8.5749393921509662e-12, 8.7737895467212104e-12, 8.9547447642782725e-12, 
    9.1176908244475699e-12, 9.2636368215737489e-12, 9.3945528708800168e-12, 
    9.5131212881372091e-12, 9.62242324382909e-12, 9.7255894765968666e-12, 
    9.8254064923854432e-12, 9.9239660480138407e-12, 1.0022371061813527e-11, 
    1.0120528939275138e-11, 1.0217061026296981e-11, 1.0309355374879813e-11, 
    1.0393744670395659e-11, 1.046580894548681e-11, 1.0520767955467108e-11, 
    1.0553913881396265e-11, 1.0561047306757793e-11, 1.0538875616464248e-11, 
    1.0485313868930505e-11, 1.0399674829824371e-11, 1.0282724813977835e-11, 
    1.0136609156007209e-11, 9.964636514024091e-12, 9.7709806742730282e-12, 
    9.5602995934600764e-12, 9.3373268065329076e-12, 9.1064570970089859e-12, 
    8.8713752638153248e-12, 8.6347433146771146e-12, 8.3980007229486502e-12, 
    8.1612518314486359e-12, 7.9233038226395595e-12, 7.6818299442019544e-12, 
    7.4336644135993058e-12, 7.1752051463461979e-12, 6.9029204298782032e-12, 
    6.6138934233418023e-12, 6.3063701433157122e-12, 5.9802717967150575e-12, 
    5.6375885457123836e-12, 5.2826083837961111e-12, 4.9219580193324495e-12, 
    4.5644122960332732e-12, 4.2204795250593267e-12, 3.9017772083990837e-12, 
    3.6202573026518653e-12, 3.3873381309617699e-12, 3.2130272948522678e-12, 
    3.1051266127602644e-12, 3.0685922678780598e-12,
  // Sqw-Na(4, 0-1999)
    0.04301919242650231, 0.042987862512806049, 0.04289430123424124, 
    0.042739774656850936, 0.042526329879378426, 0.04225670527013347, 
    0.041934213871786682, 0.041562608079672478, 0.04114593474589312, 
    0.040688390138966815, 0.040194183700886239, 0.039667418364888664, 
    0.039111993462504838, 0.038531534135409162, 0.037929348877959228, 
    0.037308414575103865, 0.036671386356597897, 0.036020627919048663, 
    0.035358256784950644, 0.034686198334473915, 0.034006242371205135, 
    0.033320096428820667, 0.03262943091288787, 0.031935912391852408, 
    0.031241222776931796, 0.030547063628720127, 0.029855146269246034, 
    0.02916716964497312, 0.028484788881447981, 0.027809578122389846, 
    0.027142991514402262, 0.026486326077917694, 0.025840689728085928, 
    0.025206976946175168, 0.024585853655214832, 0.023977751847716496, 
    0.023382873579380129, 0.022801203198881802, 0.022232526215707083, 
    0.021676453052553321, 0.021132446066304263, 0.020599848577896311, 
    0.020077915111999727, 0.019565842480612633, 0.019062801629695435, 
    0.01856797022227849, 0.018080565730181186, 0.017599878389754419, 
    0.017125302842822206, 0.01665636676730128, 0.016192754445278248, 
    0.015734323137469895, 0.015281110397921295, 0.01483333106941453, 
    0.014391363576723539, 0.01395572615388598, 0.013527044644626427, 
    0.013106014344195326, 0.012693358879660653, 0.012289789282133239, 
    0.011895966182496312, 0.011512467519550883, 0.011139763392565696, 
    0.010778198851023518, 0.010427984623805814, 0.01008919515392338, 
    0.0097617728868878515, 0.0094455375757516516, 0.0091401993832492204, 
    0.0088453747180157992, 0.0085606039589854379, 0.0082853704248315504, 
    0.0080191200782107393, 0.007761281491454948, 0.0075112855468622711, 
    0.0072685842335170172, 0.0070326677829758285, 0.0068030793111743251, 
    0.006579426147265496, 0.0063613871563701569, 0.0061487156026490122, 
    0.0059412374279422028, 0.0057388451969441869, 0.0055414883299501477, 
    0.00534916055621337, 0.0051618857321283412, 0.0049797032526783126, 
    0.0048026542358563353, 0.0046307694917499262, 0.004464060030193351, 
    0.0043025105525441041, 0.0041460760560341481, 0.0039946813909898411, 
    0.003848223380543225, 0.0037065749557390316, 0.0035695906801766091, 
    0.0034371130306918738, 0.003308978849649482, 0.0031850254719482623, 
    0.0030650961375421355, 0.0029490444126587883, 0.0028367374490236314, 
    0.0027280580042885138, 0.002622905226822448, 0.0025211942751619792, 
    0.0024228548989661744, 0.0023278291560454726, 0.0022360684792413548, 
    0.0021475303361489337, 0.0020621747410526593, 0.0019799608786975043, 
    0.0019008440811190751, 0.0018247733610399614, 0.0017516896502537923, 
    0.0016815248236745465, 0.0016142015163545581, 0.0015496336700837247, 
    0.0014877276864404233, 0.0014283840211649643, 0.00137149903463805, 
    0.0013169669159075234, 0.0012646815205770072, 0.0012145380005742091, 
    0.0011664341492315998, 0.0011202714306962943, 0.0010759557018433991, 
    0.0010333976630040303, 0.00099251308896572432, 0.00095322289452374131, 
    0.00091545308218065388, 0.00087913460748815272, 0.0008442031843115174, 
    0.00081059904154006475, 0.00077826663663731514, 0.00074715433041271139, 
    0.00071721403049988222, 0.00068840081622611679, 0.00066067256251518857, 
    0.00063398958317240094, 0.00060831431318550129, 0.00058361104540139894, 
    0.00055984572993932557, 0.00053698583643556114, 0.00051500027134033697, 
    0.00049385933640282804, 0.00047353471103000425, 0.00045399944054687363, 
    0.00043522791408586554, 0.00041719581908730377, 0.00039988006333430099, 
    0.00038325865939554309, 0.00036731056998346763, 0.00035201551607979181, 
    0.00033735375299808574, 0.00032330582312554556, 0.00030985229801015643, 
    0.00029697352648696, 0.00028464940905909898, 0.00027285922088499082, 
    0.00026158150554796502, 0.00025079405858075839, 0.0002404740132325287, 
    0.00023059803155742994, 0.00022114259257345986, 0.00021208435749499167, 
    0.00020340058165820943, 0.00019506953544099818, 0.00018707089355325139, 
    0.00017938605420853341, 0.00017199835677092146, 0.00016489317760045054, 
    0.00015805789747078711, 0.00015148174819993074, 0.00014515555906840317, 
    0.0001390714335015429, 0.00013322239218519749, 0.00012760201974676508, 
    0.00012220414855109791, 0.00011702260582780854, 0.00011205104051270227, 
    0.0001072828353204207, 0.00010271109914125601, 9.8328726134137219e-05, 
    9.4128501786874304e-05, 9.010323321362185e-05, 8.6245881104000157e-05, 
    8.2549673674023669e-05, 7.9008188042985764e-05, 7.5615390822141956e-05, 
    7.2365636431389444e-05, 6.9253627875506791e-05, 6.6274349670128636e-05, 
    6.3422985774855221e-05, 6.0694836497467328e-05, 5.8085247383306328e-05, 
    5.5589560371195219e-05, 5.3203093471053345e-05, 5.0921150541789574e-05, 
    4.8739058116939723e-05, 4.6652222301265008e-05, 4.4656196068211729e-05, 
    4.274674615102296e-05, 4.091990921688574e-05, 3.917202898094185e-05, 
    3.7499768979814912e-05, 3.5900099371970808e-05, 3.4370259796932866e-05, 
    3.2907703481696692e-05, 3.1510030017101789e-05, 3.0174915300641442e-05, 
    2.8900047003333084e-05, 2.7683072700442237e-05, 2.6521565778480366e-05, 
    2.5413011751846751e-05, 2.4354815064221483e-05, 2.3344324150253221e-05, 
    2.2378870743000643e-05, 2.1455818280770336e-05, 2.0572613828700168e-05, 
    1.9726838131796127e-05, 1.8916249131199099e-05, 1.8138815347614371e-05, 
    1.7392736796935043e-05, 1.6676452406142348e-05, 1.5988634119679997e-05, 
    1.5328168943861342e-05, 1.4694131011667017e-05, 1.4085746335680694e-05, 
    1.3502353240123894e-05, 1.2943361530949937e-05, 1.2408213290219293e-05, 
    1.1896347800028082e-05, 1.1407172552666225e-05, 1.0940041645944829e-05, 
    1.0494242159580176e-05, 1.0068988432297985e-05, 9.6634235735087843e-06, 
    9.2766271022292644e-06, 8.9076273379829966e-06, 8.5554170801756285e-06, 
    8.2189711804524067e-06, 7.8972647955942606e-06, 7.5892913501495459e-06, 
    7.2940794845842544e-06, 7.0107084693629153e-06, 6.738321704590827e-06, 
    6.4761379934719835e-06, 6.223460296510415e-06, 5.9796816728301475e-06, 
    5.7442881348177389e-06, 5.5168582115138972e-06, 5.2970591525073555e-06, 
    5.084639901053714e-06, 4.8794212002509132e-06, 4.6812834285079394e-06, 
    4.4901529487159544e-06, 4.3059878595738056e-06, 4.1287640372375818e-06, 
    3.9584622472941452e-06, 3.7950569140864788e-06, 3.6385068918854625e-06, 
    3.4887483387773424e-06, 3.3456895913176929e-06, 3.2092078097633943e-06, 
    3.0791471211619167e-06, 2.9553180248762552e-06, 2.8374979144214813e-06, 
    2.7254326761263609e-06, 2.6188394092406513e-06, 2.5174103453422491e-06, 
    2.4208180102864281e-06, 2.328721574427774e-06, 2.240774194280506e-06, 
    2.1566309949749517e-06, 2.0759572111529619e-06, 1.998435928086871e-06, 
    1.9237748625696252e-06, 1.8517117013910795e-06, 1.7820176609120537e-06, 
    1.7144991219478872e-06, 1.6489973964003123e-06, 1.585386865536225e-06, 
    1.5235718656448581e-06, 1.4634827705916716e-06, 1.4050717266558098e-06, 
    1.3483084425131753e-06, 1.2931763412005302e-06, 1.2396692644856919e-06, 
    1.1877888026500346e-06, 1.1375422232364464e-06, 1.0889409001801832e-06, 
    1.0419991049802527e-06, 9.9673301056069348e-07, 9.5315977099903439e-07, 
    9.1129656676499368e-07, 8.7115953949310912e-07, 8.3276257551583298e-07, 
    7.9611593182161346e-07, 7.612247292073285e-07, 7.2808736672935316e-07, 
    6.9669393705248848e-07, 6.6702474461627227e-07, 6.3904904331874736e-07, 
    6.1272411612421029e-07, 5.8799481093391803e-07, 5.6479362478947233e-07, 
    5.430413912842589e-07, 5.2264857825532232e-07, 5.035171490687798e-07, 
    4.8554288966395047e-07, 4.6861806097272324e-07, 4.5263421020993682e-07, 
    4.3748496662249641e-07, 4.2306865935987857e-07, 4.0929062245507461e-07, 
    3.9606509026727103e-07, 3.8331662757096094e-07, 3.7098107672604058e-07, 
    3.5900603332035585e-07, 3.4735088059134087e-07, 3.3598642072132957e-07, 
    3.2489414217819581e-07, 3.1406515962631143e-07, 3.0349886265834851e-07, 
    2.9320131364669266e-07, 2.831834466632561e-07, 2.734591358249707e-07, 
    2.6404322146187511e-07, 2.5494959944004915e-07, 2.4618948987243939e-07, 
    2.3777000012716465e-07, 2.2969308288873283e-07, 2.2195496174880078e-07, 
    2.14546058252132e-07, 2.0745140915396565e-07, 2.006515179708787e-07, 
    1.9412354566768676e-07, 1.8784271776223873e-07, 1.8178381145640098e-07, 
    1.7592258877245521e-07, 1.7023705752511242e-07, 1.647084694952715e-07, 
    1.5932199858835175e-07, 1.5406707763194554e-07, 1.4893740519872874e-07, 
    1.4393066121752437e-07, 1.3904798884928446e-07, 1.3429331097938008e-07, 
    1.2967255140562675e-07, 1.2519282669985312e-07, 1.2086166463080586e-07, 
    1.1668629292843389e-07, 1.1267302795169969e-07, 1.0882678000034977e-07, 
    1.0515068022846166e-07, 1.0164582563870324e-07, 9.8311132785113874e-08, 
    9.5143288951282989e-08, 9.2136789821976762e-08, 8.9284055885300925e-08, 
    8.6575623137742304e-08, 8.400040726810879e-08, 8.1546041497949028e-08, 
    7.9199287131854551e-08, 7.6946510447164313e-08, 7.4774211903916851e-08, 
    7.2669583251469535e-08, 7.0621058148463057e-08, 6.8618813601152422e-08, 
    6.6655175938860381e-08, 6.4724887020343381e-08, 6.2825195576999295e-08, 
    6.0955753661630178e-08, 5.9118318483311715e-08, 5.7316281639102368e-08, 
    5.5554068995787501e-08, 5.3836470465819063e-08, 5.2167968575417285e-08, 
    5.055213487366245e-08, 4.8991155097830629e-08, 4.7485527460265161e-08, 
    4.6033957183554875e-08, 4.4633446312168841e-08, 4.3279555839626347e-08, 
    4.1966798713449297e-08, 4.0689111294486502e-08, 3.94403466799051e-08, 
    3.821473743492125e-08, 3.7007284918745092e-08, 3.5814046660533485e-08, 
    3.4632308580919337e-08, 3.3460643966268544e-08, 3.2298872663866853e-08, 
    3.1147942259428341e-08, 3.0009756087044947e-08, 2.8886972543042848e-08, 
    2.7782796072820093e-08, 2.6700774824194014e-08, 2.5644613557070939e-08, 
    2.4618005287545455e-08, 2.3624480982847571e-08, 2.2667275047841932e-08, 
    2.1749203979781983e-08, 2.0872557299601594e-08, 2.0039001883456924e-08, 
    1.9249503501802191e-08, 1.8504271055755535e-08, 1.7802730184954125e-08, 
    1.7143532295659346e-08, 1.652460375631288e-08, 1.5943236779587924e-08, 
    1.5396220273295453e-08, 1.4880004570951185e-08, 1.4390890333973804e-08, 
    1.3925228510375148e-08, 1.3479616348778719e-08, 1.3051073736755844e-08, 
    1.2637185431746438e-08, 1.2236197347482764e-08, 1.1847059583561335e-08, 
    1.1469413793273804e-08, 1.110352829577522e-08, 1.0750189265543313e-08, 
    1.0410560632677347e-08, 1.0086027521235768e-08, 9.7780387860090778e-09, 
    9.4879624110429223e-09, 9.2169647685684299e-09, 8.9659200830341402e-09, 
    8.7353523246021166e-09, 8.5254072559196703e-09, 8.3358496849720037e-09, 
    8.166079163788371e-09, 8.0151577325800618e-09, 7.8818444614148707e-09, 
    7.7646341396812746e-09, 7.6617995740924187e-09, 7.5714392282347727e-09, 
    7.4915325659108084e-09, 7.4200052875941276e-09, 7.3548047376032519e-09, 
    7.2939833796938777e-09, 7.2357850195814698e-09, 7.1787261660328081e-09, 
    7.1216629763308969e-09, 7.0638345319156387e-09, 7.0048743903639383e-09, 
    6.9447858315602382e-09, 6.8838801784226187e-09, 6.8226825161506268e-09, 
    6.761813351278428e-09, 6.7018584340174277e-09, 6.6432406591639875e-09, 
    6.5861084209335657e-09, 6.5302529043710299e-09, 6.475063900227333e-09, 
    6.4195292963747365e-09, 6.3622789684788077e-09, 6.3016688816632052e-09, 
    6.2358975361602484e-09, 6.1631436025342686e-09, 6.0817121304387174e-09, 
    5.990176070904755e-09, 5.8875009267287211e-09, 5.7731421002377264e-09, 
    5.6471075482624505e-09, 5.5099813757363765e-09, 5.3629077893127299e-09, 
    5.2075378378993726e-09, 5.0459445801512733e-09, 4.8805141583531757e-09, 
    4.7138218679369636e-09, 4.5485024742248918e-09, 4.3871237870024503e-09, 
    4.2320710943491113e-09, 4.0854485483276316e-09, 3.949001458484504e-09, 
    3.8240616731926834e-09, 3.711516246883399e-09, 3.6117985366122781e-09, 
    3.5248995531059267e-09, 3.4503972201280149e-09, 3.3875006758578867e-09, 
    3.3351069437842476e-09, 3.2918670827492174e-09, 3.2562591640234715e-09, 
    3.2266650003477116e-09, 3.2014475999205274e-09, 3.1790258555528211e-09, 
    3.1579430677714371e-09, 3.1369256344946774e-09, 3.1149289906337212e-09, 
    3.0911680295722747e-09, 3.0651306764796255e-09, 3.0365740534252416e-09, 
    3.0055042962330465e-09, 2.9721420228900135e-09, 2.9368768348801924e-09, 
    2.9002146750610154e-09, 2.8627225119887126e-09, 2.8249745453665935e-09, 
    2.7875039081060674e-09, 2.7507629060340119e-09, 2.7150940971850577e-09, 
    2.6807131677374205e-09, 2.6477038636097931e-09, 2.6160239111184165e-09, 
    2.5855203932595956e-09, 2.5559522057602421e-09, 2.5270171508769985e-09, 
    2.4983808682763688e-09, 2.4697052089922547e-09, 2.44067374510414e-09, 
    2.4110128344357365e-09, 2.3805070302583193e-09, 2.3490084742936799e-09, 
    2.3164403191313475e-09, 2.2827949126974454e-09, 2.2481276973785731e-09, 
    2.212548151019771e-09, 2.1762088911086463e-09, 2.1392941900685334e-09, 
    2.1020086248473718e-09, 2.0645665395027473e-09, 2.0271824608022873e-09, 
    1.9900626501072052e-09, 1.9533976544865503e-09, 1.9173559365969878e-09, 
    1.8820785969357538e-09, 1.8476755613734148e-09, 1.8142235771957212e-09, 
    1.7817665604138251e-09, 1.7503186328721203e-09, 1.7198701557884538e-09, 
    1.6903964803862945e-09, 1.6618689802007112e-09, 1.6342672424053065e-09, 
    1.6075911967257832e-09, 1.5818715328883315e-09, 1.5571770377241238e-09, 
    1.5336174981357367e-09, 1.5113415072826037e-09, 1.4905288924645992e-09, 
    1.4713783619429357e-09, 1.4540913827817418e-09, 1.4388539788644067e-09, 
    1.4258181615901576e-09, 1.4150850658787298e-09, 1.4066913169263744e-09, 
    1.4006000689234315e-09, 1.3966973463004626e-09, 1.3947940401093768e-09, 
    1.3946330647401434e-09, 1.3959009848867816e-09, 1.3982429050480943e-09, 
    1.401279408839478e-09, 1.4046241639603592e-09, 1.407901091277166e-09, 
    1.4107599985403552e-09, 1.4128900194920197e-09, 1.414030209451302e-09, 
    1.4139771670882979e-09, 1.4125894334137267e-09, 1.409788887746821e-09, 
    1.4055591554440427e-09, 1.3999414774932972e-09, 1.393028256387279e-09, 
    1.3849547714043149e-09, 1.3758894296384303e-09, 1.3660231489102602e-09, 
    1.3555582458445156e-09, 1.3446974763396146e-09, 1.3336335862878745e-09, 
    1.3225399359468783e-09, 1.311562501688069e-09, 1.300813676431712e-09, 
    1.2903680205196622e-09, 1.28026027304203e-09, 1.2704855766555553e-09, 
    1.2610020814098103e-09, 1.2517356998379455e-09, 1.2425869369557547e-09, 
    1.2334393428134518e-09, 1.2241692194858218e-09, 1.2146558425236938e-09, 
    1.204791586077937e-09, 1.1944910319496464e-09, 1.1836983649799308e-09, 
    1.1723922704516895e-09, 1.1605878787102876e-09, 1.1483354564154925e-09, 
    1.135715952969078e-09, 1.1228337237050015e-09, 1.1098072180782071e-09, 
    1.0967584401344403e-09, 1.0838023202797092e-09, 1.0710369722930824e-09, 
    1.0585358229056259e-09, 1.0463422487880423e-09, 1.0344672390658353e-09, 
    1.0228900957923082e-09, 1.011562051473822e-09, 1.0004122722446123e-09, 
    9.893556647341272e-10, 9.7830161891973418e-10, 9.6716301069178579e-10, 
    9.5586458218442805e-10, 9.4435016929377934e-10, 9.325881583088324e-10, 
    9.2057491280740551e-10, 9.0833592505803596e-10, 8.9592476018079134e-10, 
    8.8341983008228266e-10, 8.7091939840739085e-10, 8.585351100406112e-10, 
    8.463845953474835e-10, 8.3458361904795009e-10, 8.2323842432683086e-10, 
    8.1243874275449346e-10, 8.0225205105715753e-10, 7.9271944115583489e-10, 
    7.838534629574436e-10, 7.7563801976212466e-10, 7.6803038883878562e-10, 
    7.609650946158056e-10, 7.543593740879985e-10, 7.4811967505314253e-10, 
    7.4214872137287978e-10, 7.3635246089041707e-10, 7.3064640530251046e-10, 
    7.2496078788603825e-10, 7.1924425808266311e-10, 7.1346576560379002e-10, 
    7.0761469065162446e-10, 7.0169922198027453e-10, 6.9574329190351981e-10, 
    6.8978232827410286e-10, 6.8385834701382923e-10, 6.780146940851051e-10, 
    6.722910176984672e-10, 6.6671874463466104e-10, 6.6131748000279441e-10, 
    6.560925209992466e-10, 6.5103369249413253e-10, 6.4611549934747966e-10, 
    6.4129863129412856e-10, 6.365326005145727e-10, 6.3175940653557957e-10, 
    6.2691783682850313e-10, 6.2194818238875954e-10, 6.1679694739058435e-10, 
    6.1142127194949618e-10, 6.0579264887437981e-10, 5.9989977576660121e-10, 
    5.9375020964440317e-10, 5.8737081072213395e-10, 5.808068126750857e-10, 
    5.7411968886653286e-10, 5.6738387729571153e-10, 5.6068266036466405e-10, 
    5.5410340251644413e-10, 5.4773260217766208e-10, 5.4165096537324668e-10, 
    5.3592898100556349e-10, 5.3062314734998396e-10, 5.2577321399258737e-10, 
    5.2140046734198332e-10, 5.1750720858007798e-10, 5.1407731741315652e-10, 
    5.1107785737256763e-10, 5.0846147193907157e-10, 5.0616945251698358e-10, 
    5.0413516175490164e-10, 5.0228767227476374e-10, 5.0055535713326609e-10, 
    4.9886932799907747e-10, 4.9716649272840389e-10, 4.9539224399928946e-10, 
    4.9350255148643352e-10, 4.9146552334634434e-10, 4.892622780900153e-10, 
    4.8688718614161733e-10, 4.843473707473596e-10, 4.8166160224692484e-10, 
    4.7885853354838356e-10, 4.7597444989425471e-10, 4.7305059367970394e-10, 
    4.701302930499768e-10, 4.672559754745421e-10, 4.6446637152599009e-10, 
    4.6179395703220668e-10, 4.5926290184517196e-10, 4.5688753509756636e-10, 
    4.5467150467531297e-10, 4.5260757184144646e-10, 4.5067812287966918e-10, 
    4.4885623547453503e-10, 4.4710735296590174e-10, 4.4539132515258081e-10, 
    4.4366481106694633e-10, 4.4188379986499647e-10, 4.4000620583855457e-10, 
    4.3799430586898038e-10, 4.358169695399209e-10, 4.3345146657100639e-10, 
    4.308848557924158e-10, 4.2811475281014073e-10, 4.2514955865334839e-10, 
    4.2200803539576188e-10, 4.1871833923853829e-10, 4.15316507819677e-10, 
    4.1184459528277696e-10, 4.0834847488942241e-10, 4.0487557224992187e-10, 
    4.0147255787885914e-10, 3.9818324142915326e-10, 3.9504669489828817e-10, 
    3.9209576779082407e-10, 3.8935595003635432e-10, 3.8684470997319658e-10, 
    3.8457119438712342e-10, 3.8253634601983853e-10, 3.8073328947205845e-10, 
    3.7914804812239222e-10, 3.777604305696324e-10, 3.7654513897560528e-10, 
    3.754729583057513e-10, 3.7451209517642977e-10, 3.7362953685271203e-10, 
    3.7279246757536649e-10, 3.7196962905894517e-10, 3.711326364718739e-10, 
    3.7025709953148477e-10, 3.69323592416354e-10, 3.6831827012280533e-10, 
    3.6723322765560274e-10, 3.6606642326879603e-10, 3.6482128379036785e-10, 
    3.6350590960990431e-10, 3.6213202140299016e-10, 3.6071364409116202e-10, 
    3.5926572543145361e-10, 3.5780270072609017e-10, 3.5633723480413456e-10, 
    3.5487912539214818e-10, 3.5343459029252851e-10, 3.5200587282331081e-10, 
    3.5059130825957618e-10, 3.4918573207584921e-10, 3.4778129648920825e-10, 
    3.4636849031029014e-10, 3.4493738962732086e-10, 3.4347888442263919e-10, 
    3.4198587723106804e-10, 3.4045421891825396e-10, 3.38883384473419e-10, 
    3.3727671451034624e-10, 3.3564129577601021e-10, 3.3398736545488177e-10, 
    3.3232741209535744e-10, 3.3067492786778367e-10, 3.2904304810237455e-10, 
    3.274430983776193e-10, 3.2588328419435914e-10, 3.2436756422139133e-10, 
    3.2289491275215895e-10, 3.2145894250621801e-10, 3.2004804415104187e-10, 
    3.1864594226465528e-10, 3.1723271555741561e-10, 3.1578609880744937e-10, 
    3.1428307661510491e-10, 3.1270152871481456e-10, 3.1102188703139769e-10, 
    3.0922861074371389e-10, 3.0731141625046919e-10, 3.0526612309880573e-10, 
    3.030951451732324e-10, 3.008074777412967e-10, 2.9841832693632784e-10, 
    2.9594829864850286e-10, 2.9342229514505495e-10, 2.9086811643080334e-10, 
    2.8831494637711015e-10, 2.8579173764380363e-10, 2.8332566662341352e-10, 
    2.809406959923234e-10, 2.786564080848452e-10, 2.7648706071548949e-10, 
    2.7444106723610445e-10, 2.7252079217997558e-10, 2.7072275274182111e-10, 
    2.6903813565438604e-10, 2.6745364867671887e-10, 2.659525473704107e-10, 
    2.6451585409851595e-10, 2.6312358157409295e-10, 2.617559713944276e-10, 
    2.6039457977112972e-10, 2.5902322874177207e-10, 2.5762870345059185e-10, 
    2.5620124411333809e-10, 2.5473473614287167e-10, 2.5322670725773692e-10, 
    2.5167804725311083e-10, 2.500925865284025e-10, 2.484764783003087e-10, 
    2.4683753479177902e-10, 2.451844597389284e-10, 2.4352613949635698e-10, 
    2.4187097019537007e-10, 2.4022630851095507e-10, 2.385980654887181e-10, 
    2.3699049126148671e-10, 2.3540612827222313e-10, 2.3384597246681509e-10, 
    2.3230975440817729e-10, 2.307963764916037e-10, 2.2930436951497386e-10, 
    2.2783238995429287e-10, 2.2637963291258157e-10, 2.2494618143253902e-10, 
    2.2353319463838573e-10, 2.2214298729147314e-10, 2.2077892842732343e-10, 
    2.1944527503693731e-10, 2.181468764607275e-10, 2.1688885714291434e-10, 
    2.1567627877507788e-10, 2.1451382779939141e-10, 2.134055268753269e-10, 
    2.1235451767791849e-10, 2.113628447651477e-10, 2.1043132058038063e-10, 
    2.095593686372063e-10, 2.0874491932111859e-10, 2.0798428639735267e-10, 
    2.0727210297823541e-10, 2.0660126934088053e-10, 2.05963008513054e-10, 
    2.0534697469619862e-10, 2.0474153018127012e-10, 2.0413411341742397e-10, 
    2.0351177708993474e-10, 2.0286178450211433e-10, 2.0217232097822173e-10, 
    2.0143317421715828e-10, 2.0063639571931102e-10, 1.9977680222215118e-10, 
    1.988523384864556e-10, 1.9786418256032318e-10, 1.9681664900773238e-10, 
    1.9571681917916316e-10, 1.9457401692543382e-10, 1.9339909467739426e-10, 
    1.9220368732911217e-10, 1.9099943398215703e-10, 1.8979730550102182e-10, 
    1.8860703562484772e-10, 1.8743674551230992e-10, 1.8629273119693236e-10, 
    1.8517944806889403e-10, 1.8409959400401271e-10, 1.8305432321764492e-10, 
    1.8204346585334935e-10, 1.8106578366806278e-10, 1.8011914210408453e-10, 
    1.7920069615562705e-10, 1.7830698728502028e-10, 1.7743408472903771e-10, 
    1.7657770088770567e-10, 1.7573341099625301e-10, 1.74896912805724e-10, 
    1.7406441085731986e-10, 1.732330065109683e-10, 1.7240114825434298e-10, 
    1.7156899874204213e-10, 1.7073870116094346e-10, 1.6991440922754223e-10, 
    1.6910212546948408e-10, 1.6830921959396421e-10, 1.6754374769199575e-10, 
    1.6681352397458628e-10, 1.6612513748699703e-10, 1.6548292917184035e-10, 
    1.6488815397102582e-10, 1.6433831750602743e-10, 1.6382691629981631e-10, 
    1.6334352340868637e-10, 1.6287431339925005e-10, 1.6240290999544455e-10, 
    1.619115633298477e-10, 1.6138246890637883e-10, 1.607991605336464e-10, 
    1.6014777641576865e-10, 1.5941817033120141e-10, 1.5860464771154224e-10, 
    1.5770641434539268e-10, 1.5672758709457031e-10, 1.5567689409105772e-10, 
    1.545670311315308e-10, 1.5341384111967631e-10, 1.5223531443429725e-10, 
    1.5105059910102153e-10, 1.498790054318112e-10, 1.4873915587325411e-10, 
    1.4764823757249314e-10, 1.4662143820762507e-10, 1.4567150520651813e-10, 
    1.4480844659534092e-10, 1.4403931229643257e-10, 1.4336806577991187e-10, 
    1.4279548124878285e-10, 1.4231912651874965e-10, 1.4193335678168642e-10, 
    1.4162943912935414e-10, 1.4139574617448146e-10, 1.4121812729632987e-10, 
    1.4108040201392156e-10, 1.4096505795929471e-10, 1.4085403896279512e-10, 
    1.407296873024112e-10, 1.4057565874139561e-10, 1.40377848876252e-10, 
    1.4012511394360021e-10, 1.3980983316830138e-10, 1.3942815153103134e-10, 
    1.3897994078759003e-10, 1.3846841737264895e-10, 1.3789953893593332e-10, 
    1.3728114356482563e-10, 1.3662203705815674e-10, 1.3593105042607361e-10, 
    1.3521622951614177e-10, 1.3448417583308999e-10, 1.3373968360911939e-10, 
    1.3298560854080324e-10, 1.3222303370952161e-10, 1.3145161482508018e-10, 
    1.3067010563783466e-10, 1.2987691149027352e-10, 1.2907066012377783e-10, 
    1.2825062447977667e-10, 1.2741704812006626e-10, 1.2657124750988316e-10, 
    1.2571557673316646e-10, 1.2485320904337275e-10, 1.2398784384094689e-10, 
    1.2312334352413739e-10, 1.2226342050436731e-10, 1.2141134282306809e-10, 
    1.2056981916342562e-10, 1.1974092095986768e-10, 1.189262238617587e-10, 
    1.1812698523380851e-10, 1.1734445015783392e-10, 1.1658014277445632e-10, 
    1.1583618898751266e-10, 1.1511554030352353e-10, 1.1442215772845656e-10, 
    1.1376103947205728e-10, 1.1313819145503242e-10, 1.1256043622917565e-10, 
    1.1203518395399691e-10, 1.1157008930363137e-10, 1.1117271408749409e-10, 
    1.1085012013650418e-10, 1.1060851529813389e-10, 1.10452870864103e-10, 
    1.103865960220068e-10, 1.1041120675064453e-10, 1.1052607602596268e-10, 
    1.1072816044534551e-10, 1.1101181387386337e-10, 1.1136864835406032e-10, 
    1.1178748121655373e-10, 1.1225434183212526e-10, 1.1275266880593744e-10, 
    1.1326357732322178e-10, 1.1376634723978228e-10, 1.1423901331058526e-10, 
    1.1465915322080898e-10, 1.1500473041395391e-10, 1.1525506417255926e-10, 
    1.1539176059279317e-10, 1.1539963923758756e-10, 1.1526749215433798e-10, 
    1.1498871084183651e-10, 1.1456163067976859e-10, 1.1398965409189048e-10, 
    1.1328104760862039e-10, 1.1244851458457643e-10, 1.1150845295400632e-10, 
    1.1048008316619597e-10, 1.0938438318793289e-10, 1.0824301860667388e-10, 
    1.0707724288399707e-10, 1.0590694983859818e-10, 1.0474985844885256e-10, 
    1.0362095721230092e-10, 1.0253217950879344e-10, 1.014923852850318e-10, 
    1.0050755878996039e-10, 9.9581259763541915e-11, 9.8715189533973692e-11, 
    9.7909880212534465e-11, 9.7165319675802416e-11, 9.6481558775907312e-11, 
    9.5859104993910839e-11, 9.5299161106821546e-11, 9.480361567668801e-11, 
    9.4374842951966931e-11, 9.4015281743035121e-11, 9.3726931871725195e-11, 
    9.3510750610679221e-11, 9.3366119836534874e-11, 9.3290355345138047e-11, 
    9.3278436681611302e-11, 9.332288575784093e-11, 9.3413911803851579e-11, 
    9.3539736684124557e-11, 9.3687139470558362e-11, 9.3842107405105996e-11, 
    9.3990594237346187e-11, 9.4119267959278607e-11, 9.4216255541814599e-11, 
    9.4271744156948991e-11, 9.4278502801379374e-11, 9.4232212296073007e-11, 
    9.4131665142392086e-11, 9.3978757886245814e-11, 9.3778363566443658e-11, 
    9.3538009132135694e-11, 9.3267456114168305e-11, 9.2978124689828811e-11, 
    9.2682456623269534e-11, 9.2393170959704806e-11, 9.212253104957987e-11, 
    9.1881582679956415e-11, 9.1679491253755732e-11, 9.1522956312309069e-11, 
    9.1415812190877722e-11, 9.1358787231947828e-11, 9.1349506577815009e-11, 
    9.1382668580820158e-11, 9.1450448727814797e-11, 9.1543005878449937e-11, 
    9.1649123283087216e-11, 9.1756841932087878e-11, 9.1854090573130641e-11, 
    9.1929201321963778e-11, 9.1971326920331447e-11, 9.1970676763392434e-11, 
    9.1918647206417731e-11, 9.1807791303443519e-11, 9.1631744944731815e-11, 
    9.1385061779775789e-11, 9.1063110816942293e-11, 9.0661977374663236e-11, 
    9.0178499580650209e-11, 8.9610360818975009e-11, 8.8956340843924612e-11, 
    8.8216600334736117e-11, 8.7393076691438801e-11, 8.6489841169401803e-11, 
    8.5513458939105597e-11, 8.4473187743829944e-11, 8.33810840348008e-11, 
    8.2251860440522404e-11, 8.110256650380396e-11, 7.9952007168614158e-11, 
    7.8820001116435623e-11, 7.7726441874893831e-11, 7.6690309456592427e-11, 
    7.5728628047724343e-11, 7.4855544612795548e-11, 7.4081519164184736e-11, 
    7.3412786994216115e-11, 7.2851073865528982e-11, 7.2393646890276237e-11, 
    7.2033642287745715e-11, 7.1760701323056594e-11, 7.1561797116339677e-11, 
    7.1422240580088307e-11, 7.1326716002695993e-11, 7.1260332118866738e-11, 
    7.1209537955313426e-11, 7.1162915757862928e-11, 7.1111692777904941e-11, 
    7.1050072492059198e-11, 7.0975241913297762e-11, 7.0887176625741879e-11, 
    7.078818492217377e-11, 7.0682289003120065e-11, 7.0574462991692915e-11, 
    7.0469828713497737e-11, 7.0372843433887578e-11, 7.0286600989494114e-11, 
    7.0212248748676185e-11, 7.0148659261426393e-11, 7.0092309847249548e-11, 
    7.0037468594268327e-11, 6.9976598821162745e-11, 6.9901010287687304e-11, 
    6.9801643248903809e-11, 6.9669946590894091e-11, 6.9498712495887861e-11, 
    6.9282826711890229e-11, 6.9019823733120773e-11, 6.8710198148521493e-11, 
    6.8357445841947016e-11, 6.7967846097430046e-11, 6.7549981175375277e-11, 
    6.7114102512010108e-11, 6.6671371183507263e-11, 6.6233088320609815e-11, 
    6.5809946474884866e-11, 6.5411418801012264e-11, 6.5045289828417337e-11, 
    6.4717371211934696e-11, 6.4431374139931995e-11, 6.4188950805684374e-11, 
    6.3989839563922945e-11, 6.3832093144448974e-11, 6.3712319377748008e-11, 
    6.3625939358564203e-11, 6.3567402829303616e-11, 6.353037974926779e-11, 
    6.3507912077331712e-11, 6.3492568046561158e-11, 6.3476594612451293e-11, 
    6.3452113579762706e-11, 6.3411368830519933e-11, 6.3347023789391745e-11, 
    6.3252526069653725e-11, 6.3122490148516764e-11, 6.295306819174795e-11, 
    6.274229210506198e-11, 6.2490284823128544e-11, 6.219936465005658e-11, 
    6.1873960407777088e-11, 6.1520365341254107e-11, 6.1146301160049478e-11, 
    6.0760366187680324e-11, 6.0371365233470203e-11, 5.9987631703410276e-11, 
    5.9616378142480787e-11, 5.9263149057125429e-11, 5.8931424208903719e-11, 
    5.86224161162337e-11, 5.8335070115529485e-11, 5.8066263021563262e-11, 
    5.7811167042656509e-11, 5.756374447097376e-11, 5.7317305517293116e-11, 
    5.7065088327915731e-11, 5.6800794298158079e-11, 5.6519042938276215e-11, 
    5.6215709608802642e-11, 5.5888136429300848e-11, 5.5535211233939399e-11, 
    5.5157336009755982e-11, 5.4756287266773259e-11, 5.4335019544709546e-11, 
    5.3897422239299242e-11, 5.3448079816543092e-11, 5.2992011469235922e-11, 
    5.2534463881265716e-11, 5.2080726810483392e-11, 5.1635985722979505e-11, 
    5.1205196890969559e-11, 5.0793013087744561e-11, 5.0403687500539517e-11, 
    5.0041014732602287e-11, 4.9708252172786948e-11, 4.9408043472977204e-11, 
    4.9142332115328758e-11, 4.8912269712958783e-11, 4.8718133158950286e-11, 
    4.8559265280078638e-11, 4.8434019231802142e-11, 4.8339769852417764e-11, 
    4.8272954573901306e-11, 4.8229172561851437e-11, 4.8203326563965169e-11, 
    4.8189811017616703e-11, 4.8182725362394894e-11, 4.8176100994965953e-11, 
    4.8164121081977682e-11, 4.8141315945551022e-11, 4.8102734707541237e-11, 
    4.804407242572979e-11, 4.7961742442297382e-11, 4.7852943837820618e-11, 
    4.7715663476132277e-11, 4.7548692339349303e-11, 4.7351621955174342e-11, 
    4.7124853174488772e-11, 4.6869590768021526e-11, 4.6587878065712514e-11, 
    4.6282593680056975e-11, 4.5957472242638921e-11, 4.5617070882602956e-11, 
    4.5266730751815943e-11, 4.4912473058408938e-11, 4.4560867784250846e-11, 
    4.4218828555139332e-11, 4.3893396101934222e-11, 4.3591449608151792e-11, 
    4.3319432560648499e-11, 4.3083032982128098e-11, 4.2886896263614433e-11, 
    4.2734342380028251e-11, 4.2627130746437099e-11, 4.2565263490650414e-11, 
    4.2546868467645699e-11, 4.256813716017606e-11, 4.2623383904422103e-11, 
    4.2705166172025148e-11, 4.2804543273917689e-11, 4.2911395138444367e-11, 
    4.3014879090025615e-11, 4.3103901231145769e-11, 4.3167690426730034e-11, 
    4.319634163912325e-11, 4.3181372094773679e-11, 4.3116180939145138e-11, 
    4.2996449188774958e-11, 4.2820376074323029e-11, 4.2588804617142362e-11, 
    4.230515190390164e-11, 4.1975224617601023e-11, 4.1606852579114179e-11, 
    4.1209443076473637e-11, 4.0793425069443559e-11, 4.0369685191376937e-11, 
    3.9948954783507549e-11, 3.9541302373289532e-11, 3.9155646087800799e-11, 
    3.8799438199892954e-11, 3.8478431915867071e-11, 3.8196648459968422e-11, 
    3.7956445769524625e-11, 3.7758751908517518e-11, 3.7603381983062435e-11, 
    3.7489459486258416e-11, 3.7415807543812757e-11, 3.738139666888973e-11, 
    3.7385659169343957e-11, 3.7428766043615533e-11, 3.7511729063401925e-11, 
    3.763641227779177e-11, 3.7805346468659899e-11, 3.8021482026825613e-11, 
    3.828777147957251e-11, 3.8606762810386424e-11, 3.898009135231902e-11, 
    3.9408060840595363e-11, 3.9889229228072221e-11, 4.0420127527450112e-11, 
    4.099505197703958e-11, 4.1606038671552932e-11, 4.22429180222711e-11, 
    4.289355423041661e-11, 4.354415637556674e-11, 4.4179726605665115e-11, 
    4.478454134789644e-11, 4.5342735230410834e-11, 4.5838841681099479e-11, 
    4.625839144739496e-11, 4.6588441071500952e-11, 4.681808308296275e-11, 
    4.693885232126823e-11, 4.6945099823581289e-11, 4.6834190934922952e-11, 
    4.6606666314943702e-11, 4.6266228963479517e-11, 4.5819658085289655e-11, 
    4.5276552254204394e-11, 4.4649019049476844e-11, 4.3951220997897961e-11, 
    4.3198890200129017e-11, 4.2408751875224705e-11, 4.1597968215988646e-11, 
    4.0783531820329079e-11, 3.9981740528432492e-11, 3.9207685887827609e-11, 
    3.8474845447279837e-11, 3.7794727607962022e-11, 3.71766522149185e-11, 
    3.662758559205176e-11, 3.6152108363574257e-11, 3.5752443141767933e-11, 
    3.5428591241252429e-11, 3.5178484761119008e-11, 3.4998243176084641e-11, 
    3.4882418116476536e-11, 3.4824286821108682e-11, 3.481613524554293e-11, 
    3.4849566234738105e-11, 3.4915755377196233e-11, 3.5005740105999583e-11, 
    3.5110662192073571e-11, 3.5222027501428993e-11, 3.5331919701347486e-11, 
    3.5433237591615163e-11, 3.5519892148097072e-11, 3.5587010419442334e-11, 
    3.5631086838205932e-11, 3.5650124256584047e-11, 3.5643686880771868e-11, 
    3.5612922155670642e-11, 3.5560453861497946e-11, 3.5490213961460317e-11, 
    3.5407156892802889e-11, 3.5316901467166279e-11, 3.5225276049951018e-11, 
    3.5137850014021668e-11, 3.5059436287717131e-11, 3.4993650455477085e-11, 
    3.4942530483162565e-11, 3.4906292458915291e-11, 3.4883214188735345e-11, 
    3.4869700360348793e-11, 3.4860498624675444e-11, 3.4849088341244978e-11, 
    3.4828160774409516e-11, 3.479022181296823e-11, 3.472819890392758e-11, 
    3.4636070034894571e-11, 3.450938526124683e-11, 3.4345725244741143e-11, 
    3.4144981328894292e-11, 3.3909501499166398e-11, 3.3644029190895151e-11, 
    3.3355496766609685e-11, 3.3052640646561639e-11, 3.2745513161129863e-11, 
    3.2444872216061671e-11, 3.2161557780031734e-11, 3.1905826842121896e-11, 
    3.1686768981459908e-11, 3.15117668720449e-11, 3.1386101400454328e-11, 
    3.1312670927465615e-11, 3.1291873617940137e-11, 3.1321632492491032e-11, 
    3.1397572299868621e-11, 3.151329019758499e-11, 3.1660746607429227e-11, 
    3.1830698465951315e-11, 3.2013188989925787e-11, 3.2197997614974144e-11, 
    3.2375100804210425e-11, 3.2535078852693874e-11, 3.266947217572426e-11, 
    3.2771043828327429e-11, 3.2834005660718343e-11, 3.2854157094906397e-11, 
    3.2828969396915551e-11, 3.2757584342926186e-11, 3.2640779020764483e-11, 
    3.2480850124818562e-11, 3.2281464346768895e-11, 3.2047445884070858e-11, 
    3.1784553158975581e-11, 3.1499191722198519e-11, 3.1198158332579451e-11, 
    3.0888353031034087e-11, 3.0576542095364567e-11, 3.0269135153980867e-11, 
    2.9972026028434173e-11, 2.9690468436109337e-11, 2.9429028816857369e-11, 
    2.9191556358087991e-11, 2.898121394515102e-11, 2.8800508190724843e-11, 
    2.8651338952173958e-11, 2.8535027325130356e-11, 2.8452333252794866e-11, 
    2.8403439860559139e-11, 2.8387942322459743e-11, 2.840479539294367e-11, 
    2.845229801830303e-11, 2.8528092443735754e-11, 2.8629211883169201e-11, 
    2.8752170120129618e-11, 2.8893134416756017e-11, 2.9048132798033569e-11, 
    2.9213331965589971e-11, 2.9385313506728165e-11, 2.9561366868552141e-11, 
    2.9739716227349793e-11, 2.9919704806265288e-11, 3.0101852248332442e-11, 
    3.0287816412846327e-11, 3.0480210582797105e-11, 3.0682315560024355e-11, 
    3.0897685464812638e-11, 3.1129695656903136e-11, 3.1381047311287551e-11, 
    3.1653309268471755e-11, 3.1946510218422028e-11, 3.2258851505551021e-11, 
    3.2586526229911444e-11, 3.2923726559211065e-11, 3.3262784182844411e-11, 
    3.359447501372247e-11, 3.390844822286276e-11, 3.4193766964592085e-11, 
    3.4439473212835206e-11, 3.4635203120582285e-11, 3.4771752106417177e-11, 
    3.4841584860438743e-11, 3.4839236893015935e-11, 3.4761607198810619e-11, 
    3.4608099062043734e-11, 3.4380647386972875e-11, 3.4083589937582151e-11, 
    3.3723445688219872e-11, 3.3308571470589333e-11, 3.2848776955910718e-11, 
    3.2354850241306439e-11, 3.1838095641213682e-11, 3.130985972655843e-11, 
    3.0781088722791166e-11, 3.0261915132678951e-11, 2.9761329446447627e-11, 
    2.9286913513395041e-11, 2.8844670976100577e-11, 2.8438936757109245e-11, 
    2.8072401197491361e-11, 2.77461993782648e-11, 2.7460094209337623e-11, 
    2.7212726837499334e-11, 2.7001922178192471e-11, 2.6824973354325238e-11, 
    2.6678978621661059e-11, 2.6561100413104824e-11, 2.6468806219076167e-11, 
    2.6400003359700177e-11, 2.6353118863883051e-11, 2.632708312205809e-11, 
    2.6321257317584239e-11, 2.6335279137636648e-11, 2.6368911495300874e-11, 
    2.6421864836893407e-11, 2.6493660279498998e-11, 2.6583508187157016e-11, 
    2.6690265231702296e-11, 2.68124135456011e-11, 2.694809372662135e-11, 
    2.7095155771605385e-11, 2.7251219874541765e-11, 2.7413698827878182e-11, 
    2.7579824622024442e-11, 2.7746615387768457e-11, 2.7910835080624197e-11, 
    2.8068933504955779e-11, 2.8217002475759704e-11, 2.8350763081120209e-11, 
    2.8465622847463187e-11, 2.855677804513842e-11, 2.8619418151240169e-11, 
    2.8648991139124675e-11, 2.8641527265134215e-11, 2.8593966024831523e-11, 
    2.8504498594122039e-11, 2.8372847715510535e-11, 2.8200474302525327e-11, 
    2.7990650114001669e-11, 2.7748417009406021e-11, 2.7480380083420798e-11, 
    2.7194370416185237e-11, 2.6898961338293454e-11, 2.6602892237372934e-11, 
    2.6314422596464715e-11, 2.6040677215267904e-11, 2.5787011486413054e-11, 
    2.555648576364043e-11, 2.5349466229656606e-11, 2.5163424922160931e-11, 
    2.4992934917073183e-11, 2.4829922552311128e-11, 2.4664109636089208e-11, 
    2.4483680229851996e-11, 2.4276085015947717e-11, 2.4028964236270803e-11, 
    2.3731066007684689e-11, 2.3373153724705885e-11, 2.2948784944394814e-11, 
    2.2454926346260371e-11, 2.1892341321362643e-11, 2.1265745912708478e-11, 
    2.0583700350867548e-11, 1.9858269687345302e-11, 1.9104467070572786e-11, 
    1.8339547091697674e-11, 1.7582150404594335e-11, 1.6851424688642736e-11, 
    1.6166134536335943e-11, 1.554382429889151e-11, 1.500007806151644e-11, 
    1.4547920591348541e-11, 1.4197362858649701e-11, 1.3955130932286898e-11, 
    1.3824545315444417e-11, 1.3805579281039005e-11, 1.3895025580460161e-11, 
    1.4086800005760973e-11, 1.4372317774693679e-11, 1.4740920755156097e-11, 
    1.5180340494990044e-11, 1.5677162186453807e-11, 1.6217264809524424e-11, 
    1.6786260437690249e-11, 1.7369894552382422e-11, 1.7954420896349952e-11, 
    1.8526968223273929e-11, 1.9075888844269713e-11, 1.9591075489482309e-11, 
    2.0064280020502814e-11, 2.0489376953806083e-11, 2.0862590935703241e-11, 
    2.1182625181090436e-11, 2.1450693199948602e-11, 2.1670421968266165e-11, 
    2.1847600102286914e-11, 2.1989770788136181e-11, 2.2105684845742075e-11, 
    2.2204637172270372e-11, 2.2295724780516149e-11, 2.2387103060244312e-11, 
    2.2485266374147697e-11, 2.2594480614960755e-11, 2.2716374683423234e-11, 
    2.2849750130159514e-11, 2.2990663414882599e-11, 2.3132746121532817e-11, 
    2.3267753380483966e-11, 2.3386294786997034e-11, 2.3478661575435213e-11, 
    2.3535690137896753e-11, 2.3549556291158507e-11, 2.3514438604030978e-11, 
    2.3426970475051133e-11, 2.3286473410183745e-11, 2.3094929491797716e-11, 
    2.285672196762523e-11, 2.2578193926057448e-11, 2.2267063213467246e-11, 
    2.1931784000504278e-11, 2.1580921185350605e-11, 2.1222591531334722e-11, 
    2.0864028259961394e-11, 2.0511299149111715e-11, 2.0169189073285954e-11, 
    1.9841211137725821e-11, 1.9529766326796716e-11, 1.9236354683911481e-11, 
    1.8961837470034638e-11, 1.870668932083101e-11, 1.8471211095606724e-11, 
    1.8255681179752239e-11, 1.8060441044464592e-11, 1.7885914670469348e-11, 
    1.773257049662671e-11, 1.7600855858959068e-11, 1.7491121436805938e-11, 
    1.7403541596742875e-11, 1.7338077414002384e-11, 1.7294452725236942e-11, 
    1.7272162384585942e-11, 1.7270507569960104e-11, 1.7288648286651345e-11, 
    1.732566618068044e-11, 1.7380611022252005e-11, 1.7452555175226661e-11, 
    1.7540638027624267e-11, 1.7644095018839286e-11, 1.7762297282647447e-11, 
    1.7894768869052503e-11, 1.8041224970493779e-11, 1.8201582796304546e-11, 
    1.837596982492625e-11, 1.8564700873139401e-11, 1.8768233573909248e-11, 
    1.898707173065565e-11, 1.922162737643181e-11, 1.9472049120983215e-11, 
    1.9738025528000815e-11, 2.0018584904430967e-11, 2.0311901777140658e-11, 
    2.061517069338649e-11, 2.092454725733738e-11, 2.1235161920803975e-11, 
    2.1541272589822433e-11, 2.1836488011534938e-11, 2.2114076669132278e-11, 
    2.2367345876338349e-11, 2.259004390108104e-11, 2.2776746776237389e-11, 
    2.2923199265886763e-11, 2.3026578329960607e-11, 2.3085648928851452e-11, 
    2.3100810860183667e-11, 2.3074024588686577e-11, 2.3008644144310791e-11, 
    2.2909167926208716e-11, 2.2780936512952455e-11, 2.2629813044608731e-11, 
    2.2461878413440397e-11, 2.2283140518422976e-11, 2.2099320429002311e-11, 
    2.1915672022123213e-11, 2.1736865992656195e-11, 2.156693554251913e-11, 
    2.1409256614472062e-11, 2.1266539618872197e-11, 2.1140852113493602e-11, 
    2.1033651913629069e-11, 2.0945797754241167e-11, 2.0877583274500756e-11, 
    2.0828767322272613e-11, 2.0798596640940154e-11, 2.0785863922956576e-11, 
    2.0788967235903666e-11, 2.0805990388105e-11, 2.083479247199121e-11, 
    2.0873109919235051e-11, 2.0918629227941235e-11, 2.0969054305069971e-11, 
    2.1022142517455228e-11, 2.1075702397874007e-11, 2.1127536148384523e-11, 
    2.117536809097207e-11, 2.1216749934097012e-11, 2.1248966085693147e-11, 
    2.1268961255686622e-11, 2.1273317685375431e-11, 2.1258299139835855e-11, 
    2.1219969999323135e-11, 2.1154376393942959e-11, 2.1057803541354786e-11, 
    2.0927061482409984e-11, 2.0759778928332667e-11, 2.0554670960239911e-11, 
    2.0311742504602126e-11, 2.0032415046973909e-11, 1.9719542174791873e-11, 
    1.9377328636977249e-11, 1.9011152064398496e-11, 1.8627318429973834e-11, 
    1.8232771668609092e-11, 1.783478887975743e-11, 1.7440690546445766e-11, 
    1.7057590833117138e-11, 1.669218926290104e-11, 1.6350598874660689e-11, 
    1.6038221465351677e-11, 1.5759621462142506e-11, 1.551841484939124e-11, 
    1.5317131778363932e-11, 1.5157044999968156e-11, 1.5038001634866329e-11, 
    1.4958231411821202e-11, 1.4914172249032596e-11, 1.4900358927401988e-11, 
    1.490940094337506e-11, 1.4932084361154059e-11, 1.4957606889448314e-11, 
    1.4973989158172074e-11, 1.49686163242349e-11, 1.492889542335819e-11, 
    1.4843016221389165e-11, 1.4700705110673052e-11, 1.4493955277652026e-11, 
    1.4217655548754874e-11, 1.3870055013434655e-11, 1.3453037943637863e-11, 
    1.2972178726348222e-11, 1.2436552824368204e-11, 1.1858348322541894e-11, 
    1.125227628062629e-11, 1.0634835690226229e-11, 1.0023490048403494e-11, 
    9.435794150971075e-12, 8.8885519199194757e-12, 8.3970248948706463e-12, 
    7.9742617172547862e-12, 7.6305747090491517e-12, 7.3731755761861848e-12, 
    7.2059998577264943e-12, 7.1297022052623153e-12, 7.1418281676931916e-12, 
    7.2371221531178354e-12, 7.4079787590197387e-12, 7.6449586171541735e-12, 
    7.9373773853451355e-12, 8.273898547059272e-12, 8.643120527926865e-12, 
    9.0341088265174155e-12, 9.4368599701526952e-12, 9.842664292804574e-12, 
    1.0244373547615131e-11, 1.0636548319940112e-11, 1.1015492295062246e-11, 
    1.1379176493484476e-11, 1.1727083561675956e-11, 1.2059958321255312e-11, 
    1.2379482943841382e-11, 1.2687926520136478e-11, 1.2987767121436506e-11, 
    1.3281303111655023e-11, 1.3570291837740973e-11, 1.3855627413992901e-11, 
    1.4137081496755369e-11, 1.4413119107989246e-11, 1.4680810819233188e-11, 
    1.4935845731942402e-11, 1.5172653880058884e-11, 1.5384633354890896e-11, 
    1.5564488323366636e-11, 1.5704640866421442e-11, 1.5797727809611884e-11, 
    1.5837130562351761e-11, 1.5817517557648881e-11, 1.5735364245118096e-11, 
    1.5589409954092028e-11, 1.5381010051091238e-11, 1.5114357125548867e-11, 
    1.4796528963202049e-11, 1.4437354084454903e-11, 1.4049088056429272e-11, 
    1.3645893969745413e-11, 1.3243177238076393e-11, 1.285678002008227e-11, 
    1.2502121413407257e-11, 1.2193326979606487e-11, 1.1942417666170258e-11, 
    1.175862637464557e-11, 1.1647897516813786e-11, 1.1612598700297974e-11, 
    1.1651492521133286e-11, 1.1759930787380171e-11, 1.1930282485036607e-11, 
    1.2152516576704198e-11, 1.241490807747762e-11, 1.2704789956735907e-11, 
    1.3009275316351818e-11, 1.3315913989863944e-11, 1.3613223383219163e-11, 
    1.389107222750314e-11, 1.4140924990331821e-11, 1.435594560294228e-11, 
    1.4531008658337802e-11, 1.4662619750723692e-11, 1.474881409421037e-11, 
    1.4789054270185068e-11, 1.4784142610288127e-11, 1.4736130590113713e-11, 
    1.4648279696999352e-11, 1.4524997320340654e-11, 1.4371766162602629e-11, 
    1.4195020115326175e-11, 1.4001965938373677e-11, 1.3800319888711027e-11, 
    1.3597982979940074e-11, 1.3402628966216324e-11, 1.3221279614300471e-11, 
    1.3059820649899428e-11, 1.2922577228260962e-11, 1.2811914548231288e-11, 
    1.272794631812136e-11, 1.2668362343104188e-11, 1.2628412107971378e-11, 
    1.2601034391910816e-11, 1.2577188523858583e-11, 1.2546323438075377e-11, 
    1.2497022762424803e-11, 1.241773256166495e-11, 1.229760047716717e-11, 
    1.2127309234558916e-11, 1.1899882335411741e-11, 1.1611410175744105e-11, 
    1.1261620463955534e-11, 1.085422541376081e-11, 1.0397065165933234e-11, 
    9.9019683465824241e-12, 9.384361116966348e-12, 8.8626130922617029e-12, 
    8.3571812065453368e-12, 7.8895748525537584e-12, 7.4812172200768766e-12, 
    7.1522807077388335e-12, 6.9205576097798266e-12, 6.8004350802094422e-12, 
    6.8020755486622998e-12, 6.9307944193141724e-12, 7.1867440848565146e-12, 
    7.5648707396015673e-12, 8.0551936000414142e-12, 8.6433190925392593e-12, 
    9.3112409901262685e-12, 1.0038301551483953e-11, 1.0802290201687248e-11, 
    1.1580573771681512e-11, 1.2351223302451468e-11, 1.3094018535978263e-11, 
    1.3791315569075528e-11, 1.4428688744584387e-11, 1.4995353769815837e-11, 
    1.5484320403790698e-11, 1.5892344191364392e-11, 1.6219623625435241e-11, 
    1.6469358061227447e-11, 1.6647185571238642e-11, 1.6760539762346907e-11, 
    1.6817998123669354e-11, 1.6828667633516258e-11, 1.6801627065365559e-11, 
    1.6745467988839173e-11, 1.6667939603952914e-11, 1.6575718806273499e-11, 
    1.6474258753402831e-11, 1.6367766686154051e-11, 1.6259248833292688e-11, 
    1.6150644870020103e-11, 1.6042997696055653e-11, 1.5936692865496852e-11, 
    1.5831714648459836e-11, 1.5727925124393687e-11, 1.5625349095784751e-11, 
    1.5524452262933025e-11, 1.5426371150195808e-11, 1.5333113610649415e-11, 
    1.524767629605457e-11, 1.5174083325035151e-11, 1.5117311871463656e-11, 
    1.5083113749044103e-11, 1.5077709533509614e-11, 1.5107386850282937e-11, 
    1.5178000718746749e-11, 1.529441381336842e-11, 1.5459917591741757e-11, 
    1.567568850619917e-11, 1.5940309952547963e-11, 1.6249448256537772e-11, 
    1.6595688461253834e-11, 1.6968610082434231e-11, 1.735508973686326e-11, 
    1.7739844470045091e-11, 1.8106201730470914e-11, 1.8437040144765128e-11, 
    1.8715841147116687e-11, 1.8927780976798651e-11, 1.9060760922185498e-11, 
    1.9106311043400324e-11, 1.906025766089978e-11, 1.8923110217129708e-11, 
    1.8700142784913592e-11, 1.8401105491810124e-11, 1.8039627525706384e-11, 
    1.763234181435053e-11, 1.7197772199294259e-11, 1.6755111759930694e-11, 
    1.6322954002379903e-11, 1.5918088735910382e-11, 1.5554462631945869e-11, 
    1.5242368358051691e-11, 1.4987935354183822e-11, 1.4792949421005329e-11, 
    1.4654991620511509e-11, 1.4567892092642286e-11, 1.4522446970286625e-11, 
    1.4507307432786901e-11, 1.4509969849216268e-11, 1.4517768922496447e-11, 
    1.4518803820260311e-11, 1.4502708140909621e-11, 1.4461191666211552e-11, 
    1.4388364255277733e-11, 1.4280821145266401e-11, 1.4137494321721136e-11, 
    1.3959355336636786e-11, 1.3748986740026925e-11, 1.351011860879123e-11, 
    1.3247180908849403e-11, 1.2964914229933932e-11, 1.2668077608963374e-11, 
    1.2361289888518841e-11, 1.2048950234038592e-11, 1.1735247444358775e-11, 
    1.1424214362851807e-11, 1.1119794177972145e-11, 1.0825876898388315e-11, 
    1.0546280411847262e-11, 1.0284668381650773e-11, 1.0044426140878803e-11, 
    9.8284825900070908e-12, 9.6391206886524018e-12, 9.4778173657980198e-12, 
    9.3451260912980094e-12, 9.2406251589503293e-12, 9.1629632064776338e-12, 
    9.1099725589749953e-12, 9.0788526281060601e-12, 9.0663951565176314e-12, 
    9.0692376332727893e-12, 9.0840883280055524e-12, 9.1079267665931931e-12, 
    9.1381400347188101e-12, 9.1726073395371396e-12, 9.2097133375599749e-12, 
    9.248317441223344e-12, 9.2876871508463596e-12, 9.3274075840865067e-12, 
    9.3672926977566879e-12, 9.407325183872946e-12, 9.447598375770804e-12, 
    9.4883054301815153e-12, 9.5297508567099744e-12, 9.5723694860699877e-12, 
    9.6167825190034781e-12, 9.6638376701123594e-12, 9.7146541471933144e-12, 
    9.7706541515572759e-12, 9.8335699620108233e-12, 9.9054354549140858e-12, 
    9.9885404328111223e-12, 1.008536796664132e-11, 1.019848064995959e-11, 
    1.0330400939006343e-11, 1.0483442723129851e-11, 1.0659525596969536e-11, 
    1.0859975308344923e-11, 1.1085318470352961e-11, 1.1335096799539422e-11, 
    1.1607719741192276e-11, 1.1900359388594809e-11, 1.2208936248463666e-11, 
    1.252818461729697e-11, 1.285181336686706e-11, 1.317275892652858e-11, 
    1.3483532540649355e-11, 1.377661625157083e-11, 1.4044891527344863e-11, 
    1.4282080137963879e-11, 1.4483123589444322e-11, 1.4644500039862577e-11, 
    1.476443564332166e-11, 1.4842981381518781e-11, 1.4881950902226915e-11, 
    1.4884708582684746e-11, 1.4855849001747105e-11, 1.4800758310861032e-11, 
    1.4725103029063047e-11, 1.4634307480718543e-11, 1.4533051540155904e-11, 
    1.4424831294491429e-11, 1.4311634927304992e-11, 1.4193763488036036e-11, 
    1.406981267945646e-11, 1.3936824896926635e-11, 1.3790603468474174e-11, 
    1.3626160498909848e-11, 1.3438251385765153e-11, 1.3221965043102872e-11, 
    1.297330379041131e-11, 1.2689700111721148e-11, 1.2370431514308743e-11, 
    1.2016883491499231e-11, 1.1632632788594138e-11, 1.1223355467055525e-11, 
    1.0796542963800166e-11, 1.0361064279215393e-11, 9.9265996570197713e-12, 
    9.5029889800448036e-12, 9.0995593995680394e-12, 8.7244841224741842e-12, 
    8.3842217618116644e-12, 8.0830996471247399e-12, 7.8230737260246407e-12, 
    7.6036950114420246e-12, 7.4222716342147086e-12, 7.2742472547937512e-12, 
    7.1537225124158616e-12, 7.0540962513723866e-12, 6.9687609097443007e-12, 
    6.8917599966189886e-12, 6.8183564377665577e-12, 6.7454464319496937e-12, 
    6.6717652164858235e-12, 6.5978728851638365e-12, 6.5259134138271458e-12, 
    6.4591945429430377e-12, 6.4016265398660622e-12, 6.3571066755650127e-12, 
    6.3289253544946279e-12, 6.3192753377813717e-12,
  // Sqw-Na(5, 0-1999)
    0.0340203703631601, 0.034008661015146074, 0.033973578156716845, 
    0.033915257584438585, 0.033833926172579236, 0.033729901872605286, 
    0.033603592285098467, 0.03345549082891295, 0.033286169790340679, 
    0.033096270027805269, 0.032886487744043638, 0.032657559391029968, 
    0.03241024630568673, 0.032145320966586455, 0.031863556735418269, 
    0.031565722582835375, 0.031252583641228564, 0.030924907577996791, 
    0.030583475880409595, 0.030229098336948101, 0.029862628423552796, 
    0.02948497705003721, 0.029097122230574143, 0.028700112692174429, 
    0.028295064154052096, 0.02788314788996506, 0.027465572100165196, 
    0.027043557448866693, 0.026618308767582449, 0.026190985316671699, 
    0.025762672105865598, 0.025334354603729244, 0.02490689875110192, 
    0.024481037593770606, 0.024057365141013025, 0.023636337324495393, 
    0.023218279262892012, 0.022803397510625177, 0.022391795646557383, 
    0.021983491476481994, 0.021578434284576321, 0.021176520939514189, 
    0.020777610172233788, 0.020381534900737016, 0.019988112978998874, 
    0.019597157096952408, 0.019208484688829131, 0.018821928591948076, 
    0.018437348860120228, 0.018054645643621733, 0.017673772502808653, 
    0.017294749039818248, 0.016917671417716065, 0.016542719263198502, 
    0.016170157645890679, 0.01580033327112591, 0.01543366464386132, 
    0.015070626656555522, 0.014711730708533665, 0.014357501973467674, 
    0.014008455718846877, 0.013665074612047098, 0.013327788732626555, 
    0.012996959601034856, 0.01267286900922274, 0.012355712889060472, 
    0.012045599964038454, 0.011742554561476546, 0.011446522749327094, 
    0.011157380904132623, 0.010874945887190787, 0.010598986158175524, 
    0.010329233336327667, 0.010065393880957403, 0.0098071606719055196, 
    0.009554224312749075, 0.0093062839605406438, 0.0090630574269695563, 
    0.0088242902268443908, 0.0085897632010863197, 0.0083592983366528942, 
    0.0081327624570906552, 0.0079100685635096861, 0.0076911747535558907, 
    0.0074760808142564248, 0.0072648227493942851, 0.0070574656415367081, 
    0.0068540953474044196, 0.0066548095755358163, 0.0064597088979535811, 
    0.0062688882099242744, 0.0060824290846318322, 0.005900393383980968, 
    0.0057228183923946968, 0.0055497136439523406, 0.0053810595180804792, 
    0.005216807586666608, 0.005056882606632093, 0.0049011859680371025, 
    0.00474960033161579, 0.004601995125813523, 0.0044582325275341088, 
    0.0043181735283879755, 0.0041816836933032901, 0.0040486382523647994, 
    0.0039189262278680401, 0.0037924533817087825, 0.0036691438655505008, 
    0.0035489405582283967, 0.0034318041716945194, 0.0033177112895384003, 
    0.0032066515638196147, 0.0030986243324881086, 0.0029936349300495623, 
    0.0028916909503992278, 0.0027927986875315291, 0.0026969599335572038, 
    0.0026041692613638263, 0.0025144118683022129, 0.0024276620131681013, 
    0.0023438820451008959, 0.0022630220009797431, 0.0021850197361212892, 
    0.0021098015482615994, 0.002037283252518863, 0.0019673716608993781, 
    0.001899966410676241, 0.0018349620704184101, 0.0017722504317951172, 
    0.0017117228730596161, 0.0016532726614482589, 0.0015967970522174576, 
    0.0015421990464272815, 0.0014893886905656636, 0.0014382838384916941, 
    0.001388810346626552, 0.0013409017307399668, 0.0012944983692042081, 
    0.0012495463849282378, 0.0012059963691344858, 0.0011638021198610736, 
    0.001122919554990369, 0.0010833059256809014, 0.0010449194064731417, 
    0.0010077190804935639, 0.0009716652805686353, 0.00093672019778255318, 
    0.00090284863455853282, 0.00087001876366395734, 0.000838202758628325, 
    0.00080737718301786428, 0.00077752306158000121, 0.00074862559967973203, 
    0.00072067356240610955, 0.00069365836535394923, 0.00066757296070889737, 
    0.00064241062188393795, 0.00061816373644340054, 0.00059482271102318592, 
    0.00057237507545643176, 0.00055080484932995208, 0.00053009220616305442, 
    0.00051021344170816118, 0.00049114122650130052, 0.0004728451010320574, 
    0.00045529215624619235, 0.00043844783319748346, 0.00042227677344685953, 
    0.0004067436555711058, 0.0003918139617652869, 0.00037745463061237752, 
    0.00036363456617162645, 0.00035032498816562404, 0.00033749962194964934, 
    0.00032513473908150718, 0.00031320906892409603, 0.00030170360835717145, 
    0.00029060136020927211, 0.00027988703157527146, 0.00026954672112364334, 
    0.00025956762034611209, 0.00024993774809300778, 0.00024064573133160823, 
    0.00023168063850655766, 0.00022303186574412821, 0.00021468907090733231, 
    0.00020664214653844161, 0.00019888122025977511, 0.00019139667034287323, 
    0.00018417914486339393, 0.00017721957494517147, 0.00017050917573564273, 
    0.00016403943249207304, 0.00015780207296346957, 0.00015178903057143871, 
    0.00014599240523418782, 0.00014040442968450052, 0.00013501744866082404, 
    0.00012982391649355311, 0.00012481641570135, 0.00011998769576913862, 
    0.00011533072791357235, 0.0001108387689438512, 0.00010650542576244025, 
    0.0001023247118695048, 9.8291088431526138e-05, 9.4399484790554111e-05, 
    9.0645296280422312e-05, 8.7024360332033592e-05, 8.3532914557663785e-05, 
    8.016754237607967e-05, 7.6925112535394861e-05, 7.3802718579062771e-05, 
    7.0797623059961921e-05, 6.7907209464866891e-05, 6.5128942775711723e-05, 
    6.2460337764740285e-05, 5.9898932822831743e-05, 5.74422665430856e-05, 
    5.5087854464806774e-05, 5.2833164216555495e-05, 5.0675588562706911e-05, 
    4.8612417272443799e-05, 4.6640810006312662e-05, 4.4757773306877008e-05, 
    4.2960145124899025e-05, 4.1244590046826367e-05, 3.9607607556396254e-05, 
    3.8045554390708226e-05, 3.6554680533777005e-05, 3.5131176847556828e-05, 
    3.37712309913305e-05, 3.2471087304731134e-05, 3.1227105853887509e-05, 
    3.0035815915299828e-05, 2.8893959779044895e-05, 2.7798523802209398e-05, 
    2.6746754997338283e-05, 2.5736162926715334e-05, 2.4764508114933052e-05, 
    2.3829779423715258e-05, 2.2930163726580866e-05, 2.2064011692930435e-05, 
    2.1229803516199086e-05, 2.0426118024402132e-05, 1.9651607870970497e-05, 
    1.8904982527624047e-05, 1.818499972159513e-05, 1.7490464907033444e-05, 
    1.6820237455459184e-05, 1.6173241581030339e-05, 1.5548479639089846e-05, 
    1.4945045362009149e-05, 1.4362134802094467e-05, 1.3799053179040411e-05, 
    1.3255216405720676e-05, 1.2730146706135853e-05, 1.2223462367806317e-05, 
    1.1734862224014193e-05, 1.1264105899896441e-05, 1.0810991160059881e-05, 
    1.0375329866414011e-05, 9.9569241050024937e-06, 9.555543990619929e-06, 
    9.1709085248465126e-06, 8.8026706821774176e-06, 8.4504076370401528e-06, 
    8.1136167285291739e-06, 7.7917173948307679e-06, 7.4840589100631127e-06, 
    7.1899333429796999e-06, 6.9085927641615442e-06, 6.6392693931051375e-06, 
    6.3811971418817322e-06, 6.1336329096216128e-06, 5.8958760343551701e-06, 
    5.6672845136137905e-06, 5.4472869437906291e-06, 5.2353895577291658e-06, 
    5.0311782088539633e-06, 4.8343155984007504e-06, 4.6445344198772083e-06, 
    4.4616273614835027e-06, 4.2854350459273135e-06, 4.1158329979944825e-06, 
    3.9527186351049654e-06, 3.7959991053095391e-06, 3.6455805892606965e-06, 
    3.5013594699321906e-06, 3.3632155835237744e-06, 3.2310076094929635e-06, 
    3.1045705418923074e-06, 2.9837151008459886e-06, 2.8682288842799623e-06, 
    2.7578790143154395e-06, 2.6524159957807856e-06, 2.5515784727829673e-06, 
    2.4550985479653113e-06, 2.3627073217860208e-06, 2.2741403223937161e-06, 
    2.1891425310749681e-06, 2.1074727632441121e-06, 2.028907232506276e-06, 
    1.9532421978451062e-06, 1.8802956603675218e-06, 1.8099081301989281e-06, 
    1.7419425212452707e-06, 1.6762832540825192e-06, 1.6128346588342241e-06, 
    1.5515187790451089e-06, 1.4922726891063384e-06, 1.4350454572360205e-06, 
    1.3797949108587206e-06, 1.3264843885194701e-06, 1.275079682013221e-06, 
    1.2255463769758928e-06, 1.1778477803462316e-06, 1.1319435773033406e-06, 
    1.0877892887077476e-06, 1.0453365125158802e-06, 1.0045338396798787e-06, 
    9.653282532975705e-07, 9.2766676157337095e-07, 8.9149799275623184e-07, 
    8.5677349687404821e-07, 8.2344855423808982e-07, 7.9148237406960109e-07, 
    7.6083766611797393e-07, 7.3147966577057259e-07, 7.0337477494534963e-07, 
    6.7648903270061507e-07, 6.507866459166937e-07, 6.2622878928430467e-07, 
    6.0277283295880434e-07, 5.8037208439216624e-07, 5.5897605324798723e-07, 
    5.3853117642820302e-07, 5.1898188663286635e-07, 5.0027187743325147e-07, 
    4.8234541376737777e-07, 4.6514855432519983e-07, 4.4863018619424811e-07, 
    4.3274281249437372e-07, 4.1744307365137717e-07, 4.0269201450806652e-07, 
    3.8845513049870075e-07, 3.7470223469174904e-07, 3.6140718748159939e-07, 
    3.4854752421578032e-07, 3.361040092712041e-07, 3.2406013972368629e-07, 
    3.1240162139305179e-07, 3.0111584301551277e-07, 2.9019138029315086e-07, 
    2.7961756618174089e-07, 2.6938416541622232e-07, 2.5948118601937721e-07, 
    2.4989884908586599e-07, 2.4062771956768052e-07, 2.3165897929780792e-07, 
    2.2298480096846743e-07, 2.1459876374756731e-07, 2.0649623969186648e-07, 
    1.986746788013987e-07, 1.9113372869604653e-07, 1.8387514294990003e-07, 
    1.7690245598282695e-07, 1.7022043027884907e-07, 1.638343083442427e-07, 
    1.5774892539520256e-07, 1.5196775541234687e-07, 1.4649197279763665e-07, 
    1.4131961286528695e-07, 1.3644490846195365e-07, 1.3185786687798176e-07, 
    1.2754413362525233e-07, 1.2348516748084533e-07, 1.196587273565868e-07, 
    1.1603964618341658e-07, 1.1260084317736771e-07, 1.093145040030815e-07, 
    1.0615334220253055e-07, 1.0309184505142468e-07, 1.0010740615980602e-07, 
    9.7181254747382694e-08, 9.4299109154582058e-08, 9.1451506702649271e-08, 
    8.8633792523968848e-08, 8.584578155840246e-08, 8.3091138052441382e-08, 
    8.0376540709900965e-08, 7.7710717670366709e-08, 7.5103440703377287e-08, 
    7.2564563722039529e-08, 7.0103177074884975e-08, 6.7726929643657943e-08, 
    6.5441547807126561e-08, 6.325055831876776e-08, 6.1155202646954248e-08, 
    5.9154516794270266e-08, 5.7245542550508909e-08, 5.5423634471149844e-08, 
    5.3682829186893459e-08, 5.2016249356567589e-08, 5.04165202769583e-08, 
    4.8876182715577463e-08, 4.738808834369405e-08, 4.5945765335006296e-08, 
    4.4543740388412452e-08, 4.3177802101487869e-08, 4.1845188874838804e-08, 
    4.0544685484978798e-08, 3.9276615054884004e-08, 3.8042719395542024e-08, 
    3.684592870820857e-08, 3.5690031918285938e-08, 3.4579268751122302e-08, 
    3.3517873947250344e-08, 3.2509610130303697e-08, 3.1557329081536263e-08, 
    3.0662599623925762e-08, 2.9825435419031951e-08, 2.9044146897650748e-08, 
    2.8315330498853898e-08, 2.7633995431569639e-08, 2.6993815838267934e-08, 
    2.6387484637615481e-08, 2.5807136929492224e-08, 2.5244805187225002e-08, 
    2.4692867293476381e-08, 2.4144450715628827e-08, 2.3593762559589805e-08, 
    2.3036323869954038e-08, 2.2469097587136642e-08, 2.1890510434692425e-08, 
    2.1300379660727915e-08, 2.0699763386922011e-08, 2.0090758936573611e-08, 
    1.9476274864036088e-08, 1.8859800969923783e-08, 1.8245195563238004e-08, 
    1.7636502767493481e-08, 1.7037804722567551e-08, 1.6453106742806508e-08, 
    1.5886247425977482e-08, 1.5340822918701974e-08, 1.4820113592619906e-08, 
    1.4327003931087177e-08, 1.3863890376310867e-08, 1.3432577662619354e-08, 
    1.303416968886986e-08, 1.2668966163252634e-08, 1.23363792388003e-08, 
    1.2034885696800065e-08, 1.1762028427581316e-08, 1.1514477452618378e-08, 
    1.128815474130759e-08, 1.1078420558997362e-08, 1.0880311642418903e-08, 
    1.068881547889537e-08, 1.0499159678628495e-08, 1.0307093012637775e-08, 
    1.0109134244438534e-08, 9.9027675227524594e-09, 9.6865676866592829e-09, 
    9.4602455895355719e-09, 9.2246109005829406e-09, 8.9814577424170573e-09, 
    8.7333850648344642e-09, 8.4835692624598589e-09, 8.2355093544935661e-09, 
    7.9927662070160243e-09, 7.7587155676332933e-09, 7.5363317355987552e-09, 
    7.3280139493312839e-09, 7.1354628255867454e-09, 6.9596090563275398e-09, 
    6.8005927119193219e-09, 6.6577880996406573e-09, 6.529867591819046e-09, 
    6.4148966551848748e-09, 6.3104527302326402e-09, 6.2137607973314352e-09, 
    6.1218394183818204e-09, 6.0316512876709436e-09, 5.9402528588079003e-09, 
    5.8449372799293751e-09, 5.7433649519179781e-09, 5.6336756026880493e-09, 
    5.5145761861107953e-09, 5.3853992177256233e-09, 5.2461276869036014e-09, 
    5.0973840921432939e-09, 4.940383766125502e-09, 4.7768547503573052e-09, 
    4.6089292454516207e-09, 4.4390135241071758e-09, 4.2696450398409868e-09, 
    4.1033460717449081e-09, 3.9424835948636941e-09, 3.7891441346424023e-09, 
    3.6450312665339696e-09, 3.5113913299196511e-09, 3.3889710622914676e-09, 
    3.2780082539646372e-09, 3.1782546544984928e-09, 3.0890280275506001e-09, 
    3.0092887382613692e-09, 2.9377346932541653e-09, 2.8729076901819152e-09, 
    2.8133035048844259e-09, 2.7574782048482099e-09, 2.7041433970174605e-09, 
    2.6522442324838269e-09, 2.6010150735779784e-09, 2.5500096796748074e-09, 
    2.4991044279331344e-09, 2.4484754525969158e-09, 2.3985522963654685e-09, 
    2.3499527711028053e-09, 2.3034048669435318e-09, 2.2596626948354301e-09, 
    2.2194235585399124e-09, 2.183253111468961e-09, 2.151524454897522e-09, 
    2.1243758580121554e-09, 2.1016898105086749e-09, 2.0830944126600856e-09, 
    2.0679860059872412e-09, 2.0555704478050414e-09, 2.0449188470631205e-09, 
    2.0350328400096739e-09, 2.0249138086957285e-09, 2.0136307243783391e-09, 
    2.00038149322691e-09, 1.9845437494241882e-09, 1.9657118504073397e-09, 
    1.9437182699523427e-09, 1.9186385377920432e-09, 1.8907803123432661e-09, 
    1.8606579136550659e-09, 1.8289547602189323e-09, 1.7964765278594276e-09, 
    1.7640985086795452e-09, 1.7327105795680304e-09, 1.7031634106884279e-09, 
    1.6762189978207101e-09, 1.6525084702064011e-09, 1.6324992650480127e-09, 
    1.6164732212976098e-09, 1.6045162307533214e-09, 1.5965194526466849e-09, 
    1.5921911817120214e-09, 1.5910780341816651e-09, 1.5925934928158771e-09, 
    1.5960517291552769e-09, 1.600704404843901e-09, 1.6057783978721605e-09, 
    1.6105124635651876e-09, 1.6141913218853809e-09, 1.6161757890080832e-09, 
    1.6159281311191491e-09, 1.6130318449815626e-09, 1.607205512632556e-09, 
    1.5983102786590346e-09, 1.5863509833482417e-09, 1.5714708028037254e-09, 
    1.5539397332487177e-09, 1.5341372828123081e-09, 1.5125302568034584e-09, 
    1.4896466138459416e-09, 1.4660469204286742e-09, 1.4422948932137452e-09, 
    1.418928928034142e-09, 1.3964362229906751e-09, 1.3752311346485767e-09, 
    1.3556389089715192e-09, 1.3378856436452777e-09, 1.3220946691911047e-09, 
    1.3082892324094767e-09, 1.2964007016614032e-09, 1.2862813609671368e-09, 
    1.2777204488147285e-09, 1.2704621960903292e-09, 1.2642244507546406e-09, 
    1.2587168241243015e-09, 1.2536573071862304e-09, 1.248786738889388e-09, 
    1.243880522407142e-09, 1.2387574523760089e-09, 1.2332854119793421e-09, 
    1.2273840707787418e-09, 1.2210245499876489e-09, 1.2142263236182553e-09, 
    1.2070514462151846e-09, 1.1995964818449601e-09, 1.1919824057174813e-09, 
    1.1843430618852781e-09, 1.1768126933121279e-09, 1.1695134073226504e-09, 
    1.1625433143620311e-09, 1.1559663432440056e-09, 1.149804497059921e-09, 
    1.1440333615159128e-09, 1.1385812928576499e-09, 1.133332570621054e-09, 
    1.1281342849673484e-09, 1.12280653378898e-09, 1.1171549834059901e-09, 
    1.1109848046075432e-09, 1.1041146438280043e-09, 1.0963894753847194e-09, 
    1.0876910956382172e-09, 1.077945513235747e-09, 1.0671265795956761e-09, 
    1.0552558262623579e-09, 1.042398630082457e-09, 1.0286574279323735e-09, 
    1.0141627090430341e-09, 9.9906289561294004e-10, 9.8351404339323286e-10, 
    9.676704129516172e-10, 9.5167656721211119e-10, 9.3566163902697785e-10, 
    9.1973589047925993e-10, 9.0398966111852038e-10, 8.8849428014299434e-10, 
    8.7330467023232711e-10, 8.5846290250247007e-10, 8.4400226937150586e-10, 
    8.2995116177898758e-10, 8.1633643346121559e-10, 8.0318576504583754e-10, 
    7.9052897339011229e-10, 7.7839811130823161e-10, 7.6682657131867319e-10, 
    7.5584726493697375e-10, 7.4549030586159535e-10, 7.357803655725316e-10, 
    7.2673414146860031e-10, 7.1835810824246221e-10, 7.1064686537413133e-10, 
    7.035821507667705e-10, 6.9713265516180634e-10, 6.9125456138308942e-10, 
    6.8589283503981056e-10, 6.8098304962498764e-10, 6.764537266669618e-10, 
    6.7222894442900179e-10, 6.6823118798668137e-10, 6.643842354617352e-10, 
    6.6061606296799969e-10, 6.5686155528754571e-10, 6.5306503554358289e-10, 
    6.4918238526397153e-10, 6.4518269885613998e-10, 6.4104922409251508e-10, 
    6.367795656880061e-10, 6.3238492857354894e-10, 6.2788844657308762e-10, 
    6.2332252789851568e-10, 6.1872547985993859e-10, 6.1413752491322001e-10, 
    6.0959666105279604e-10, 6.0513464532045139e-10, 6.0077362410593636e-10, 
    5.9652366044159636e-10, 5.9238155512865706e-10, 5.883310254859138e-10, 
    5.8434433326923318e-10, 5.8038511982370359e-10, 5.7641224973760587e-10, 
    5.7238419951051953e-10, 5.6826357624796135e-10, 5.6402128841057115e-10, 
    5.596399818055698e-10, 5.5511636394916886e-10, 5.5046228260727505e-10, 
    5.4570438125375989e-10, 5.4088247493151871e-10, 5.3604670582729945e-10, 
    5.3125383130496644e-10, 5.2656283030703877e-10, 5.2203031676327368e-10, 
    5.1770600093107505e-10, 5.1362863237571546e-10, 5.0982265435292994e-10, 
    5.062959138298124e-10, 5.0303850104195308e-10, 5.0002293056019806e-10, 
    4.972055687713056e-10, 4.9452930859566381e-10, 4.9192722979768511e-10, 
    4.8932706817585301e-10, 4.8665608809694186e-10, 4.8384607638044494e-10, 
    4.8083798678658644e-10, 4.7758598197323882e-10, 4.7406046045355522e-10, 
    4.7024993413850114e-10, 4.6616152468710812e-10, 4.6182015486422795e-10, 
    4.5726643135298493e-10, 4.5255350178554962e-10, 4.4774308522701133e-10, 
    4.4290111332977143e-10, 4.3809326002959929e-10, 4.333808155891973e-10, 
    4.2881714772728295e-10, 4.244450797198674e-10, 4.2029527264219056e-10, 
    4.1638574947471786e-10, 4.1272243753187649e-10, 4.093006950821998e-10, 
    4.0610751557775149e-10, 4.0312425807086422e-10, 4.0032954769309875e-10, 
    3.9770216113435521e-10, 3.9522355252674121e-10, 3.9287991964427325e-10, 
    3.9066357037067184e-10, 3.8857357848460611e-10, 3.8661559428624351e-10, 
    3.8480095869003345e-10, 3.8314510918675671e-10, 3.8166549614583419e-10, 
    3.8037912474917264e-10, 3.793000193583511e-10, 3.7843677239890647e-10, 
    3.7779047573283869e-10, 3.7735318542069301e-10, 3.771071488067451e-10, 
    3.7702481219802649e-10, 3.7706971935771578e-10, 3.7719814159090891e-10, 
    3.7736139008755739e-10, 3.7750851327186235e-10, 3.7758920417816614e-10, 
    3.7755660250844236e-10, 3.7736979163704384e-10, 3.7699574439220884e-10, 
    3.7641065421826042e-10, 3.7560052522286928e-10, 3.7456111827469214e-10, 
    3.7329727039688036e-10, 3.7182179136902732e-10, 3.7015404192302775e-10, 
    3.6831840030577851e-10, 3.6634269531023358e-10, 3.6425677984849346e-10, 
    3.6209123037503194e-10, 3.5987626799375979e-10, 3.5764081653531999e-10, 
    3.5541174181144377e-10, 3.5321317436265562e-10, 3.5106595737226438e-10, 
    3.4898713348839728e-10, 3.4698956390489299e-10, 3.4508162318428765e-10, 
    3.4326707878782644e-10, 3.4154511281903055e-10, 3.39910593556895e-10, 
    3.3835451460167942e-10, 3.3686467674563668e-10, 3.3542649755880438e-10, 
    3.340239622329703e-10, 3.3264057679778481e-10, 3.3126033160401356e-10, 
    3.2986852893092141e-10, 3.2845251011910755e-10, 3.2700213056474111e-10, 
    3.2551009815497212e-10, 3.2397206912874187e-10, 3.2238660355283561e-10, 
    3.2075496047808043e-10, 3.1908082272428991e-10, 3.1736993800606501e-10, 
    3.1562979332778831e-10, 3.1386923286331723e-10, 3.1209816823663948e-10, 
    3.1032724499563262e-10, 3.085675775882484e-10, 3.068304124114638e-10, 
    3.0512680472921751e-10, 3.03467200267077e-10, 3.0186097997995188e-10, 
    3.0031591403638293e-10, 2.9883761615733264e-10, 2.9742893507261662e-10, 
    2.960894597959307e-10, 2.9481509435038817e-10, 2.9359784390857164e-10, 
    2.9242580446819718e-10, 2.9128346891791629e-10, 2.9015228952616566e-10, 
    2.8901155797454326e-10, 2.8783947753739493e-10, 2.8661444273899005e-10, 
    2.8531633651128536e-10, 2.8392781268429625e-10, 2.8243538375617666e-10, 
    2.8083026960655342e-10, 2.791088686239101e-10, 2.7727286755477964e-10, 
    2.7532891163498775e-10, 2.7328795020461125e-10, 2.7116422030107482e-10, 
    2.6897408958603283e-10, 2.6673474676104872e-10, 2.644629769719398e-10, 
    2.6217405705407326e-10, 2.5988092186990588e-10, 2.5759363144494373e-10, 
    2.553192248553984e-10, 2.5306189932434894e-10, 2.5082354809605384e-10, 
    2.4860451215133612e-10, 2.4640453194070041e-10, 2.4422370898491972e-10, 
    2.4206344553453407e-10, 2.3992718725947159e-10, 2.3782093986032669e-10, 
    2.35753450001266e-10, 2.3373607812737556e-10, 2.3178229630824506e-10, 
    2.2990694446062349e-10, 2.2812522280635933e-10, 2.2645159314428533e-10, 
    2.2489863920937075e-10, 2.2347603692301936e-10, 2.22189697244091e-10, 
    2.2104120874177935e-10, 2.200275692959706e-10, 2.1914130349750193e-10, 
    2.1837087126521753e-10, 2.1770139685814897e-10, 2.1711556788954111e-10, 
    2.165946845091446e-10, 2.1611969609678332e-10, 2.156721884116961e-10, 
    2.152351811682604e-10, 2.147937462127807e-10, 2.1433535366599584e-10, 
    2.1385001644365098e-10, 2.1333018362465e-10, 2.1277051692816057e-10, 
    2.1216753519756874e-10, 2.1151926043154059e-10, 2.1082483850440762e-10, 
    2.1008427383000424e-10, 2.0929820355372682e-10, 2.0846780518572761e-10, 
    2.0759473717118828e-10, 2.0668118150428131e-10, 2.0572985714615218e-10, 
    2.0474407602742105e-10, 2.0372773453437514e-10, 2.0268529317278311e-10, 
    2.0162167359921106e-10, 2.005421529848908e-10, 1.9945219952624603e-10, 
    1.9835732678882424e-10, 1.9726291529237299e-10, 1.9617409057150206e-10, 
    1.9509559338625414e-10, 1.9403171635706185e-10, 1.9298622953363431e-10, 
    1.9196238232783165e-10, 1.9096288525771382e-10, 1.8998995582769728e-10, 
    1.8904533155379676e-10, 1.8813033442978782e-10, 1.8724589851882693e-10, 
    1.8639263561977556e-10, 1.8557083334905972e-10, 1.847804750895636e-10, 
    1.8402120637941047e-10, 1.8329227658248083e-10, 1.8259242596588646e-10, 
    1.8191976276738549e-10, 1.8127157899533728e-10, 1.8064419926710214e-10, 
    1.8003279105364451e-10, 1.7943123937090721e-10, 1.788320589248929e-10, 
    1.7822640786468285e-10, 1.7760415702434938e-10, 1.7695411581457334e-10, 
    1.7626434195379517e-10, 1.7552258634024362e-10, 1.747168051134175e-10, 
    1.738357738652834e-10, 1.7286972515420165e-10, 1.718109950363478e-10, 
    1.7065461807172239e-10, 1.6939886809071384e-10, 1.6804562978623748e-10, 
    1.6660066102612356e-10, 1.6507363986894588e-10, 1.6347804895298007e-10, 
    1.6183083885480581e-10, 1.6015194332739406e-10, 1.5846360828705908e-10, 
    1.5678961950559293e-10, 1.5515441284577425e-10, 1.5358215234224381e-10, 
    1.5209575734465142e-10, 1.5071598245744005e-10, 1.4946050849665568e-10, 
    1.4834316136907076e-10, 1.4737323461397491e-10, 1.4655500676284334e-10, 
    1.4588745858004644e-10, 1.4536426623937818e-10, 1.4497405314366069e-10, 
    1.4470097258069779e-10, 1.44525550148808e-10, 1.4442580619808764e-10, 
    1.4437853396054086e-10, 1.4436071073790866e-10, 1.4435084539046628e-10, 
    1.4433023202236134e-10, 1.44283916813458e-10, 1.4420135209626279e-10, 
    1.4407659974768327e-10, 1.4390814982721585e-10, 1.4369830622245939e-10, 
    1.4345226822614252e-10, 1.4317696206548112e-10, 1.4287982143765066e-10, 
    1.4256757308421101e-10, 1.4224523888910132e-10, 1.4191540149141543e-10, 
    1.41577833125084e-10, 1.4122947261092351e-10, 1.4086478247684227e-10, 
    1.4047636656781875e-10, 1.4005579993757473e-10, 1.3959452334734328e-10, 
    1.3908473293040584e-10, 1.3852011635236598e-10, 1.3789642031741219e-10, 
    1.3721172299134356e-10, 1.364664947093478e-10, 1.3566338763601948e-10, 
    1.3480686787652727e-10, 1.339026972487025e-10, 1.3295740622281928e-10, 
    1.3197777339054988e-10, 1.3097043477272265e-10, 1.2994158756314439e-10, 
    1.2889692882509979e-10, 1.2784167550139999e-10, 1.2678079981995075e-10, 
    1.257193053105301e-10, 1.2466259371654366e-10, 1.2361677369599949e-10, 
    1.2258894182747133e-10, 1.2158731131969954e-10, 1.2062123602579822e-10, 
    1.1970102566093649e-10, 1.1883765532923784e-10, 1.1804229496435694e-10, 
    1.1732577701585261e-10, 1.1669796884330827e-10, 1.161671768841355e-10, 
    1.1573955112755805e-10, 1.1541861895521685e-10, 1.1520488945168838e-10, 
    1.1509565296812174e-10, 1.1508489334970273e-10, 1.1516341454754198e-10, 
    1.1531906035125387e-10, 1.1553711808906424e-10, 1.1580081337798159e-10, 
    1.1609190942895468e-10, 1.1639132661546412e-10, 1.1667984835574158e-10, 
    1.1693876629571718e-10, 1.1715056129100158e-10, 1.1729948829434877e-10, 
    1.1737214904445677e-10, 1.1735792385608646e-10, 1.1724935563711734e-10, 
    1.1704237422125396e-10, 1.1673642534628014e-10, 1.1633440977213079e-10, 
    1.1584252055600085e-10, 1.1526986335355535e-10, 1.1462797395343501e-10, 
    1.1393016057915391e-10, 1.1319077502466158e-10, 1.124243675327845e-10, 
    1.1164487429329166e-10, 1.1086480558499133e-10, 1.1009457261296851e-10, 
    1.0934194678895877e-10, 1.0861175934513568e-10, 1.0790582218553167e-10, 
    1.0722313698429953e-10, 1.06560325009283e-10, 1.0591230714970901e-10, 
    1.0527309724150271e-10, 1.0463672587916591e-10, 1.0399810632941329e-10, 
    1.0335386224569497e-10, 1.0270291116114152e-10, 1.0204687219703215e-10, 
    1.0139013183115911e-10, 1.0073965125867007e-10, 1.0010447409168688e-10, 
    9.9495026436139925e-11, 9.8922226488391769e-11, 9.8396566850100649e-11, 
    9.7927176618427707e-11, 9.7521050215448226e-11, 9.718241303110606e-11, 
    9.6912381696926578e-11, 9.6708846342587967e-11, 9.6566659599201454e-11, 
    9.6478027273843471e-11, 9.643311361293855e-11, 9.6420738139397719e-11, 
    9.6429157217798912e-11, 9.6446784487994031e-11, 9.6462892193497473e-11, 
    9.6468128215457992e-11, 9.6454947266547766e-11, 9.6417844919295792e-11, 
    9.6353477400946676e-11, 9.6260610106503642e-11, 9.6139999362878664e-11, 
    9.5994149977204402e-11, 9.5827060513539796e-11, 9.5643890891330423e-11, 
    9.5450661165585652e-11, 9.5253900640021431e-11, 9.5060354662288416e-11, 
    9.4876658369075449e-11, 9.4709071026931788e-11, 9.4563193164510607e-11, 
    9.4443742622086454e-11, 9.435431446998523e-11, 9.4297208070434873e-11, 
    9.4273241414884745e-11, 9.4281633925762385e-11, 9.4319878901067834e-11, 
    9.4383702463073588e-11, 9.446701932246353e-11, 9.4561989797173278e-11, 
    9.4659101930153798e-11, 9.4747373707925762e-11, 9.4814595316310845e-11, 
    9.484771380574387e-11, 9.483325846839648e-11, 9.4757899067545772e-11, 
    9.4609008764481142e-11, 9.4375314795627366e-11, 9.4047498077928302e-11, 
    9.3618792573262398e-11, 9.3085465493631622e-11, 9.2447216637900605e-11, 
    9.1707392684521625e-11, 9.0873067083032737e-11, 8.9954914616490385e-11, 
    8.8966945547360977e-11, 8.792602880063686e-11, 8.6851321984706338e-11, 
    8.5763540665543858e-11, 8.4684174108839977e-11, 8.363461861606347e-11, 
    8.2635323269838885e-11, 8.1704935892640815e-11, 8.0859535389025267e-11, 
    8.0111946993609721e-11, 7.9471235968994402e-11, 7.8942342366280702e-11, 
    7.8525960252032724e-11, 7.8218615539344427e-11, 7.8012982492031365e-11, 
    7.7898389636870294e-11, 7.7861519751720927e-11, 7.7887202209091784e-11, 
    7.7959294151883002e-11, 7.8061538594044328e-11, 7.8178362579204292e-11, 
    7.8295545732790979e-11, 7.8400742431381097e-11, 7.8483779189279113e-11, 
    7.8536806012533737e-11, 7.8554244785347772e-11, 7.8532613814292171e-11, 
    7.8470245714516475e-11, 7.8366948014312918e-11, 7.8223652084686406e-11, 
    7.8042086848194941e-11, 7.7824483885260962e-11, 7.7573356915644421e-11, 
    7.7291310704396396e-11, 7.6980927282192072e-11, 7.6644663816751859e-11, 
    7.6284798784486795e-11, 7.5903373997417245e-11, 7.5502163528554775e-11, 
    7.5082648705800173e-11, 7.4646014987846173e-11, 7.4193167255700737e-11, 
    7.3724786996234101e-11, 7.3241425649769072e-11, 7.2743627470825924e-11, 
    7.223208984544572e-11, 7.1707836741519502e-11, 7.1172376796320042e-11, 
    7.062784629645568e-11, 7.0077099094271788e-11, 6.9523744845287841e-11, 
    6.897209170297008e-11, 6.8427035611337762e-11, 6.7893874540026464e-11, 
    6.7378072436964171e-11, 6.6884978092793028e-11, 6.6419546520918966e-11, 
    6.5986050260105991e-11, 6.558783242669452e-11, 6.5227079408625301e-11, 
    6.4904660800104721e-11, 6.4620007997625575e-11, 6.4371066723954677e-11, 
    6.4154309460898994e-11, 6.3964817866829189e-11, 6.379644792266852e-11, 
    6.3642077040608962e-11, 6.3493923597529052e-11, 6.3343962636885216e-11, 
    6.3184395927935146e-11, 6.3008167097979485e-11, 6.2809479144030967e-11, 
    6.2584289029708831e-11, 6.2330688569266308e-11, 6.2049175759751205e-11, 
    6.1742734840961816e-11, 6.1416720572034348e-11, 6.107852466083543e-11, 
    6.073705524179336e-11, 6.0402041561458756e-11, 6.0083248341170167e-11, 
    5.9789659413577044e-11, 5.9528705348362109e-11, 5.9305604258285384e-11, 
    5.9122900423532635e-11, 5.8980215505469407e-11, 5.8874263246475509e-11, 
    5.8799089998887931e-11, 5.874655022069497e-11, 5.8706935485779565e-11, 
    5.8669722575117442e-11, 5.862435515339152e-11, 5.8561006989233439e-11, 
    5.8471259343829618e-11, 5.8348648475500619e-11, 5.8189049763022366e-11, 
    5.7990890921973238e-11, 5.7755168503737036e-11, 5.748530291086039e-11, 
    5.7186841340264658e-11, 5.6867043565932359e-11, 5.653435294213963e-11, 
    5.6197843352129894e-11, 5.5866631629055537e-11, 5.5549311874399301e-11, 
    5.5253443071437547e-11, 5.4985129268994335e-11, 5.4748687595074104e-11, 
    5.4546461833388869e-11, 5.4378758981521604e-11, 5.4243907513158597e-11, 
    5.4138440134240432e-11, 5.4057352570977433e-11, 5.3994429366648191e-11, 
    5.3942588170818126e-11, 5.3894202911347044e-11, 5.3841399590039206e-11, 
    5.3776277814518814e-11, 5.3691083859659836e-11, 5.3578299250153581e-11, 
    5.3430715762668179e-11, 5.3241477156785081e-11, 5.3004166852888183e-11, 
    5.2712926487692519e-11, 5.2362672727429473e-11, 5.1949386189983618e-11, 
    5.1470504382877618e-11, 5.0925335944841562e-11, 5.0315527488680544e-11, 
    4.964544822648582e-11, 4.892250620257481e-11, 4.8157272715867752e-11, 
    4.7363422269815578e-11, 4.6557404974111179e-11, 4.5757898855719326e-11, 
    4.4985012548126768e-11, 4.4259338881902717e-11, 4.3600860080378835e-11, 
    4.3027867023607071e-11, 4.2555906834100503e-11, 4.2196911889806677e-11, 
    4.1958518694323606e-11, 4.1843689623150134e-11, 4.1850603239148735e-11, 
    4.197287502837489e-11, 4.2200002797703729e-11, 4.2518062068655149e-11, 
    4.291052478246968e-11, 4.3359164750607206e-11, 4.3844940784160489e-11, 
    4.4348839800039695e-11, 4.485256639578295e-11, 4.53391254221398e-11, 
    4.5793194613159293e-11, 4.6201385025896728e-11, 4.6552324025192361e-11, 
    4.6836678514766442e-11, 4.7047063509321101e-11, 4.7177966615783544e-11, 
    4.7225636704209528e-11, 4.7188033290376457e-11, 4.7064776967646603e-11, 
    4.685718244751166e-11, 4.6568279093659207e-11, 4.6202888876889876e-11, 
    4.5767649970514476e-11, 4.5271047762467164e-11, 4.4723330980445559e-11, 
    4.4136392589050204e-11, 4.3523508314787516e-11, 4.289901357487996e-11, 
    4.2277828117556041e-11, 4.1674967465276998e-11, 4.1104940279619889e-11, 
    4.0581190477347325e-11, 4.0115517106502751e-11, 3.9717614543369928e-11, 
    3.9394674127125972e-11, 3.9151173184561863e-11, 3.8988779527120088e-11, 
    3.8906471130283819e-11, 3.8900749647302461e-11, 3.8966057866924897e-11, 
    3.909522660586474e-11, 3.9280041185252058e-11, 3.951177055481908e-11, 
    3.9781708402822044e-11, 4.0081595887019513e-11, 4.0403999447294238e-11, 
    4.0742502928619338e-11, 4.10918358718499e-11, 4.1447804139566161e-11, 
    4.1807173969037815e-11, 4.2167408420481934e-11, 4.2526390445069089e-11, 
    4.2882069162130499e-11, 4.3232171261189596e-11, 4.3573902524566274e-11, 
    4.3903775546708127e-11, 4.4217490953396492e-11, 4.4509975497290872e-11, 
    4.4775491909659419e-11, 4.5007907828939814e-11, 4.5200993448720836e-11, 
    4.5348827929283721e-11, 4.544618389460978e-11, 4.5488925378322636e-11, 
    4.5474298302199966e-11, 4.5401184551656449e-11, 4.5270166400006348e-11, 
    4.5083536253379839e-11, 4.4845118026486567e-11, 4.4560044555334475e-11, 
    4.4234397952106906e-11, 4.3874875030530005e-11, 4.3488403278971565e-11, 
    4.308184130424263e-11, 4.2661714421128208e-11, 4.2234087403093882e-11, 
    4.1804478107153513e-11, 4.1377915574535473e-11, 4.0959026300330326e-11, 
    4.0552192231492611e-11, 4.0161674240493719e-11, 3.9791749237846047e-11, 
    3.9446735411235186e-11, 3.913097700429445e-11, 3.8848698462943286e-11, 
    3.8603814137286099e-11, 3.8399607121098644e-11, 3.82384334532308e-11, 
    3.8121366745313953e-11, 3.8047926393638825e-11, 3.8015852545888596e-11, 
    3.8021035738732294e-11, 3.805753495088634e-11, 3.8117799291187586e-11, 
    3.8192993518873262e-11, 3.8273487343686989e-11, 3.8349386866300132e-11, 
    3.8411165369028562e-11, 3.8450234905720862e-11, 3.8459510809598795e-11, 
    3.8433817292806126e-11, 3.8370202924390451e-11, 3.8268038082956695e-11, 
    3.8128986504720269e-11, 3.7956758882049835e-11, 3.7756769646600516e-11, 
    3.7535651202835889e-11, 3.730073824738624e-11, 3.7059498551973998e-11, 
    3.6819037795012452e-11, 3.6585641354857475e-11, 3.6364456391340509e-11, 
    3.6159256405198182e-11, 3.5972383180539231e-11, 3.5804770712714631e-11, 
    3.5656115586697032e-11, 3.5525109113101575e-11, 3.5409768363613416e-11, 
    3.5307745274676098e-11, 3.5216698016185038e-11, 3.5134590062642865e-11, 
    3.5059986615131723e-11, 3.4992232768914252e-11, 3.4931599331623165e-11, 
    3.4879294439781494e-11, 3.4837407457644972e-11, 3.480872927355523e-11, 
    3.4796513284151955e-11, 3.4804133558491457e-11, 3.4834728601738818e-11, 
    3.4890792774088477e-11, 3.497381679230997e-11, 3.5083945038671656e-11, 
    3.5219758588158792e-11, 3.5378131553827734e-11, 3.5554262924860879e-11, 
    3.5741814368109626e-11, 3.5933211820892571e-11, 3.6120044206081568e-11, 
    3.6293569757806419e-11, 3.644522656200515e-11, 3.6567185572000615e-11, 
    3.6652811394078665e-11, 3.6697073860366889e-11, 3.6696795975840069e-11, 
    3.665078419381122e-11, 3.6559808375553446e-11, 3.642645083146417e-11, 
    3.6254792468053349e-11, 3.6050059502402966e-11, 3.5818174915783125e-11, 
    3.5565316717883646e-11, 3.5297457522604636e-11, 3.5019992929907779e-11, 
    3.4737414256199776e-11, 3.4453105917563184e-11, 3.4169246773628921e-11, 
    3.3886854001269469e-11, 3.360592613425398e-11, 3.3325739374105304e-11, 
    3.3045210680671894e-11, 3.2763362765089994e-11, 3.2479796305048014e-11, 
    3.2195178455200688e-11, 3.191164772793588e-11, 3.1633125921836608e-11, 
    3.1365455427958211e-11, 3.111636635588399e-11, 3.0895207723005806e-11, 
    3.0712486477340273e-11, 3.0579201199794094e-11, 3.0506052581188746e-11, 
    3.0502548454110881e-11, 3.057614467424389e-11, 3.0731427380464175e-11, 
    3.0969488493588804e-11, 3.1287530126758752e-11, 3.1678748857707224e-11, 
    3.2132518715681987e-11, 3.2634898757295468e-11, 3.3169387029173602e-11, 
    3.3717908909672035e-11, 3.426191581319494e-11, 3.478355302584028e-11, 
    3.5266738102743996e-11, 3.5698128436786404e-11, 3.6067834691975015e-11, 
    3.6369877628883667e-11, 3.6602296212772854e-11, 3.676696094676324e-11, 
    3.6869061941394931e-11, 3.6916360594616967e-11, 3.6918240383575372e-11, 
    3.6884673326001194e-11, 3.6825182523480625e-11, 3.6747901658389729e-11, 
    3.6658804453544474e-11, 3.6561195979196407e-11, 3.6455490653982799e-11, 
    3.6339295691443435e-11, 3.6207798360945371e-11, 3.6054405479605475e-11, 
    3.5871541940694652e-11, 3.5651563950083333e-11, 3.5387668857892896e-11, 
    3.5074711584913881e-11, 3.4709842467712315e-11, 3.4292930803933112e-11, 
    3.3826712547012855e-11, 3.3316689104448771e-11, 3.2770782463131154e-11, 
    3.2198811480275211e-11, 3.1611843725344034e-11, 3.1021514659045072e-11, 
    3.0439357612922885e-11, 2.9876238559661501e-11, 2.9341917681438918e-11, 
    2.8844778020067786e-11, 2.8391692064177121e-11, 2.7988056424176771e-11, 
    2.7637929903774882e-11, 2.7344237229184738e-11, 2.7109009945448322e-11, 
    2.6933613593802e-11, 2.6818913454588476e-11, 2.6765379073875804e-11, 
    2.6773114310426191e-11, 2.6841803670506115e-11, 2.6970566138764138e-11, 
    2.715779570376616e-11, 2.7400964004391193e-11, 2.76964450782178e-11, 
    2.8039362887736561e-11, 2.8423525081787215e-11, 2.8841436573833243e-11, 
    2.9284419138621098e-11, 2.9742818121430021e-11, 3.0206315448326183e-11, 
    3.0664312599296873e-11, 3.1106360825500998e-11, 3.152259339359871e-11, 
    3.1904152533903649e-11, 3.2243535235105075e-11, 3.2534863810155451e-11, 
    3.2774035035330108e-11, 3.2958751738320449e-11, 3.3088415038819711e-11, 
    3.316392803945091e-11, 3.3187392050470177e-11, 3.3161762022942573e-11, 
    3.3090477450519284e-11, 3.297712012523825e-11, 3.2825120636877824e-11, 
    3.2637557853601855e-11, 3.2417034687091123e-11, 3.216568143369144e-11, 
    3.1885242003780337e-11, 3.1577253913888877e-11, 3.1243255458685588e-11, 
    3.0885039650594549e-11, 3.0504879373721619e-11, 3.010571819483691e-11, 
    2.9691269203813179e-11, 2.9266043304403347e-11, 2.8835259218816751e-11, 
    2.8404670866192965e-11, 2.7980291519341774e-11, 2.7568069723547304e-11, 
    2.717351625566697e-11, 2.6801339916450983e-11, 2.6455088646604002e-11, 
    2.6136868407315115e-11, 2.5847125618757036e-11, 2.5584542206152284e-11, 
    2.5346032613137191e-11, 2.5126869282165233e-11, 2.4920908117337703e-11, 
    2.4720932797423515e-11, 2.4519078016598669e-11, 2.4307328399778652e-11, 
    2.4078036089013361e-11, 2.3824462032152632e-11, 2.3541276916254045e-11, 
    2.3225011612300246e-11, 2.2874389672407431e-11, 2.2490565189892681e-11, 
    2.2077199498179526e-11, 2.1640398204699093e-11, 2.1188481263213532e-11, 
    2.0731638986048912e-11, 2.0281416035453181e-11, 1.9850135651923137e-11, 
    1.9450241918358571e-11, 1.9093616859148774e-11, 1.8790897399626316e-11, 
    1.855086184476326e-11, 1.8379877150494199e-11, 1.8281492619584214e-11, 
    1.8256165834955396e-11, 1.8301177037760011e-11, 1.8410697923727944e-11, 
    1.8576081178937159e-11, 1.8786295294312989e-11, 1.9028525801248293e-11, 
    1.9288883489004557e-11, 1.9553207062860702e-11, 1.9807856763495642e-11, 
    2.0040517615531083e-11, 2.0240894918460554e-11, 2.0401297617485343e-11, 
    2.051705991189654e-11, 2.0586783044508351e-11, 2.0612361838362391e-11, 
    2.0598844040061113e-11, 2.0554086350692206e-11, 2.048827576262127e-11, 
    2.0413308923862368e-11, 2.0342095588318477e-11, 2.0287804009043977e-11, 
    2.0263109545105546e-11, 2.0279440010436822e-11, 2.0346316094434676e-11, 
    2.04707536074077e-11, 2.0656813594647995e-11, 2.0905273125525822e-11, 
    2.1213478825912921e-11, 2.1575368130693664e-11, 2.1981682738078681e-11, 
    2.2420329067572931e-11, 2.287693202456442e-11, 2.3335486934347947e-11, 
    2.3779133358905901e-11, 2.4190961214433945e-11, 2.455483720200167e-11, 
    2.4856171190091099e-11, 2.5082614341845677e-11, 2.5224598495187686e-11, 
    2.5275734874269247e-11, 2.5233025955123108e-11, 2.5096888822215211e-11, 
    2.4870998239207393e-11, 2.456198019130026e-11, 2.4178957544639926e-11, 
    2.3733023480640231e-11, 2.3236651035335338e-11, 2.2703107207868494e-11, 
    2.2145876153961479e-11, 2.1578164985832724e-11, 2.101247419672442e-11, 
    2.0460266884394012e-11, 1.993174529731815e-11, 1.9435701614378409e-11, 
    1.8979452069417868e-11, 1.8568839996215034e-11, 1.820825911003745e-11, 
    1.7900725673907818e-11, 1.7647942191925693e-11, 1.7450380573691435e-11, 
    1.7307344303118824e-11, 1.7217051619844532e-11, 1.7176705267129746e-11, 
    1.7182575694607128e-11, 1.7230109098094079e-11, 1.7314052678085862e-11, 
    1.742859696053149e-11, 1.756756022933854e-11, 1.7724591271276656e-11, 
    1.7893401756975365e-11, 1.8068002357076683e-11, 1.8242957028613522e-11, 
    1.8413629486273764e-11, 1.857641023168043e-11, 1.8728914351178491e-11, 
    1.8870120320267457e-11, 1.9000461516979472e-11, 1.9121828414325711e-11, 
    1.9237482632250325e-11, 1.9351886550685498e-11, 1.9470445200532472e-11, 
    1.959917072067152e-11, 1.9744293054698334e-11, 1.9911845366828204e-11, 
    2.0107251032131196e-11, 2.0334957271110473e-11, 2.0598114660052662e-11, 
    2.0898361159678546e-11, 2.1235702553730858e-11, 2.1608475955810971e-11, 
    2.201343152470213e-11, 2.2445861662170791e-11, 2.2899783396580701e-11, 
    2.3368148201154062e-11, 2.3843060160467572e-11, 2.4315983643131741e-11, 
    2.4777940034131201e-11, 2.5219712329040919e-11, 2.5632047200833622e-11, 
    2.6005889087836989e-11, 2.6332651328861928e-11, 2.6604519199201498e-11, 
    2.6814812137893985e-11, 2.6958346133282822e-11, 2.7031807963360399e-11, 
    2.703407841105316e-11, 2.6966481081469276e-11, 2.6832918200313483e-11, 
    2.6639843170085777e-11, 2.6396072099555372e-11, 2.6112428977098245e-11, 
    2.5801230085333303e-11, 2.5475624012426766e-11, 2.5148864462555652e-11, 
    2.4833561539899368e-11, 2.4540937820102649e-11, 2.4280200619905615e-11, 
    2.4058048592760729e-11, 2.3878343333611185e-11, 2.3742001664009897e-11, 
    2.3647087359583887e-11, 2.3589088029774721e-11, 2.3561367938372342e-11, 
    2.3555728950180486e-11, 2.3563035314951443e-11, 2.3573851140813094e-11, 
    2.3579050515850301e-11, 2.3570331666321364e-11, 2.3540613741906681e-11, 
    2.3484309538936066e-11, 2.3397466496849071e-11, 2.3277767458992773e-11, 
    2.3124444823925272e-11, 2.2938095079055295e-11, 2.2720471660178101e-11, 
    2.2474233270400817e-11, 2.220270751674728e-11, 2.1909665105277334e-11, 
    2.1599127055182684e-11, 2.1275190595366883e-11, 2.0941887821249296e-11, 
    2.0603054517801632e-11, 2.0262229177024038e-11, 1.9922558264986063e-11, 
    1.9586731745452079e-11, 1.9256947133918688e-11, 1.8934916330176952e-11, 
    1.8621924334905689e-11, 1.8318941871961761e-11, 1.80267812557771e-11, 
    1.7746299503800953e-11, 1.7478591788694576e-11, 1.7225169918372294e-11, 
    1.6988075624148502e-11, 1.6769885160930294e-11, 1.6573602773478547e-11, 
    1.6402414714248668e-11, 1.6259306042435213e-11, 1.6146604094494559e-11, 
    1.6065460509243187e-11, 1.6015336869613788e-11, 1.5993589413562323e-11, 
    1.5995192635838327e-11, 1.6012663904862437e-11, 1.603621727828198e-11, 
    1.6054168293439628e-11, 1.6053554654228028e-11, 1.6020939670952506e-11, 
    1.5943339457302013e-11, 1.5809187901003135e-11, 1.5609243280092617e-11, 
    1.5337391517570679e-11, 1.499123386975521e-11, 1.4572436510187914e-11, 
    1.4086803803341444e-11, 1.3544053438156972e-11, 1.2957329600965723e-11, 
    1.2342480403096032e-11, 1.1717141048535149e-11, 1.1099720288913776e-11, 
    1.0508333347823148e-11, 9.9597826531302107e-12, 9.4686366994960568e-12, 
    9.0464922338114306e-12, 8.7014642864775567e-12, 8.4379176086572467e-12, 
    8.2564828180265415e-12, 8.1543147838227045e-12, 8.1255867128375915e-12, 
    8.1621429641530379e-12, 8.2542817830249118e-12, 8.3915743976531227e-12, 
    8.5636431806997198e-12, 8.7608750856680717e-12, 8.9749770727933945e-12, 
    9.1993767488834565e-12, 9.4294254781137958e-12, 9.6624274472068609e-12, 
    9.8975015262954124e-12, 1.0135313040256945e-11, 1.0377692657119527e-11, 
    1.0627196901736665e-11, 1.0886641967231427e-11, 1.1158636205269193e-11, 
    1.1445126891497433e-11, 1.1747011168722802e-11, 1.206380821773987e-11, 
    1.2393423458716421e-11, 1.2732011221982672e-11, 1.3073959850735998e-11, 
    1.3412012364533414e-11, 1.3737523772635781e-11, 1.4040850779382724e-11, 
    1.4311875962594691e-11, 1.4540614242082683e-11, 1.4717891068184446e-11, 
    1.4836020360713949e-11, 1.4889435891364574e-11, 1.4875218177863985e-11, 
    1.4793464693514469e-11, 1.4647447054704581e-11, 1.4443565318714448e-11, 
    1.4191050468004005e-11, 1.3901472560658588e-11, 1.3588067864612172e-11, 
    1.326494102445496e-11, 1.294622088884716e-11, 1.2645226803425031e-11, 
    1.2373701098620443e-11, 1.2141200612999169e-11, 1.1954639088721307e-11, 
    1.1818052864333287e-11, 1.1732572355404997e-11, 1.1696596651347505e-11, 
    1.1706138608337596e-11, 1.1755319172045346e-11, 1.1836938063644507e-11, 
    1.1943103599415057e-11, 1.2065835069163363e-11, 1.2197630968587934e-11, 
    1.2331916303753439e-11, 1.2463377952858872e-11, 1.2588158323005263e-11, 
    1.2703881042005834e-11, 1.2809551715675507e-11, 1.2905324583921525e-11, 
    1.2992176962161641e-11, 1.307153309921584e-11, 1.31448734517944e-11, 
    1.3213386907120569e-11, 1.3277674593835828e-11, 1.33375725110884e-11, 
    1.3392096342489318e-11, 1.343952188643289e-11, 1.3477567178843321e-11, 
    1.3503708249386137e-11, 1.3515541686606064e-11, 1.3511190663772994e-11, 
    1.3489676949708476e-11, 1.3451231787265226e-11, 1.3397482068516595e-11, 
    1.3331492326205298e-11, 1.3257627158451364e-11, 1.3181246448851221e-11, 
    1.3108220315882154e-11, 1.3044347807822124e-11, 1.2994681062888625e-11, 
    1.296286621365297e-11, 1.2950552783231022e-11, 1.2956962476093076e-11, 
    1.2978645617960752e-11, 1.3009525666002465e-11, 1.3041189185271659e-11, 
    1.306346596331208e-11, 1.3065205423137233e-11, 1.3035238736215377e-11, 
    1.2963381085326254e-11, 1.2841423706083949e-11, 1.2664004924497201e-11, 
    1.2429274612419376e-11, 1.2139261980241313e-11, 1.1799975025592517e-11, 
    1.1421155951704576e-11, 1.1015764308870092e-11, 1.0599206847761687e-11, 
    1.0188412778382105e-11, 9.800803696319996e-12, 9.453268790859451e-12, 
    9.1612064191227443e-12, 8.9377143001641589e-12, 8.792941577676584e-12, 
    8.7336941366418006e-12, 8.7632341318380848e-12, 8.8813219654732307e-12, 
    9.0844549774473348e-12, 9.3662860396275209e-12, 9.7181422696297877e-12, 
    1.0129661593007466e-11, 1.0589451378628261e-11, 1.1085751591200799e-11, 
    1.1607037065750682e-11, 1.2142555797706057e-11, 1.2682743699873734e-11, 
    1.3219522548987597e-11, 1.3746450749047717e-11, 1.4258755385202118e-11, 
    1.475322434982772e-11, 1.5228029272963044e-11, 1.5682437596949222e-11, 
    1.6116518103417511e-11, 1.6530822824958834e-11, 1.6926088739978932e-11, 
    1.7302973074561803e-11, 1.7661861731916941e-11, 1.8002726176389473e-11, 
    1.8325059498900507e-11, 1.8627871778635189e-11, 1.8909762533318041e-11, 
    1.916900575294928e-11, 1.9403711879624502e-11, 1.9611989326872622e-11, 
    1.9792130213356836e-11, 1.9942771253611826e-11, 2.0063060778761911e-11, 
    2.015276154480716e-11, 2.0212331654225362e-11, 2.0242937041439001e-11, 
    2.0246421556761612e-11, 2.0225207462768669e-11, 2.0182172056548492e-11, 
    2.0120485371224012e-11, 2.0043448871614257e-11, 1.9954325882892857e-11, 
    1.9856205397246691e-11, 1.9751884437012134e-11, 1.9643786173752122e-11, 
    1.9533901350886454e-11, 1.9423753473380489e-11, 1.9314367762637024e-11, 
    1.9206260349612959e-11, 1.9099411051759302e-11, 1.8993258614326634e-11, 
    1.8886695598729613e-11, 1.8778095879043458e-11, 1.8665367534328816e-11, 
    1.8546057172886482e-11, 1.8417483166944807e-11, 1.8276926889270996e-11, 
    1.8121822316067721e-11, 1.7949975003325859e-11, 1.7759741531977708e-11, 
    1.7550188840835234e-11, 1.732117281035032e-11, 1.7073361207862459e-11, 
    1.6808190290216522e-11, 1.6527756383472457e-11, 1.623466182045515e-11, 
    1.5931854880423208e-11, 1.5622450841930534e-11, 1.5309603452642822e-11, 
    1.4996392337768025e-11, 1.4685773124329068e-11, 1.4380567220433753e-11, 
    1.4083493527355777e-11, 1.3797215676994629e-11, 1.3524414325437e-11, 
    1.3267823515177272e-11, 1.3030251621449947e-11, 1.2814569645422945e-11, 
    1.2623638868369005e-11, 1.2460193310435633e-11, 1.232668156837118e-11, 
    1.2225084589358845e-11, 1.2156730080338037e-11, 1.2122089451695042e-11, 
    1.2120639084932942e-11, 1.2150760404675174e-11, 1.2209714033710905e-11, 
    1.2293687252146706e-11, 1.2397928539470553e-11, 1.2516942675977539e-11, 
    1.2644752461042454e-11, 1.2775175376619913e-11, 1.2902105016489455e-11, 
    1.3019782642383678e-11, 1.3123013549995376e-11, 1.3207314000987133e-11, 
    1.3269007384006465e-11, 1.3305265576549033e-11, 1.3314100260668718e-11, 
    1.3294331200243336e-11, 1.3245555833045644e-11, 1.3168143444683285e-11, 
    1.3063249335336302e-11, 1.2932852041775404e-11, 1.2779820564535478e-11, 
    1.2607957470759678e-11, 1.2422015824565516e-11, 1.2227648521699821e-11, 
    1.2031264630880682e-11, 1.1839770487474687e-11, 1.1660209127421441e-11, 
    1.149930441570631e-11, 1.1362948457442502e-11, 1.125567589822078e-11, 
    1.1180191192302486e-11, 1.1137006359745463e-11, 1.1124234306186856e-11, 
    1.1137589989278622e-11, 1.1170610123386773e-11, 1.1215078126403264e-11, 
    1.126163700155531e-11, 1.1300538377200315e-11, 1.1322435930566934e-11, 
    1.1319181270000337e-11, 1.1284516891488572e-11, 1.1214614925810046e-11, 
    1.1108417781746905e-11, 1.0967746884856297e-11, 1.0797181129791166e-11, 
    1.060372788494827e-11, 1.0396329736985754e-11, 1.0185251728803416e-11, 
    9.9814200832122594e-12, 9.7957564956509871e-12, 9.6385619980275091e-12, 
    9.5189980407549301e-12, 9.4446691030884524e-12, 9.4213245977085178e-12, 
    9.4526907252829622e-12, 9.5404001434857977e-12, 9.6840262452255492e-12, 
    9.8811953974059399e-12, 1.0127764158154629e-11, 1.041806008374305e-11, 
    1.0745159045050517e-11, 1.1101199323293206e-11, 1.1477720739360606e-11, 
    1.1866022526916135e-11, 1.2257503262249654e-11, 1.2643989512193625e-11, 
    1.3018025455741394e-11, 1.3373096104326585e-11, 1.3703787704200703e-11, 
    1.4005871149381353e-11, 1.4276300161365734e-11, 1.4513142902325614e-11, 
    1.4715438782192216e-11, 1.4883023841678977e-11, 1.5016323576583445e-11, 
    1.5116120989860619e-11, 1.5183353144448705e-11, 1.5218920293142208e-11, 
    1.5223528600424365e-11, 1.51975725766011e-11, 1.5141067923887094e-11, 
    1.505363049921279e-11, 1.4934505572413792e-11, 1.4782642584301085e-11, 
    1.4596818857148389e-11, 1.437579229825596e-11, 1.4118491509195792e-11, 
    1.3824218516582509e-11, 1.3492860770732819e-11, 1.3125091661686276e-11, 
    1.2722545283429207e-11, 1.2287949112120943e-11, 1.1825199490367427e-11, 
    1.1339372821199175e-11, 1.0836653742470584e-11, 1.0324190690703275e-11, 
    9.8098736571578727e-12, 9.3020360654885599e-12, 8.8091182517736333e-12, 
    8.3392861339156607e-12, 7.9000465415104411e-12, 7.4978903838282833e-12, 
    7.1379708967185558e-12, 6.8238675111644045e-12, 6.5574329612184868e-12, 
    6.3387571730706666e-12, 6.1662313880984879e-12, 6.0367218426419566e-12, 
    5.9458347758798688e-12, 5.8882253658821036e-12, 5.8579638636138932e-12, 
    5.8488870550748468e-12, 5.854935795087929e-12, 5.8704376712191396e-12, 
    5.8903357279474296e-12, 5.9103545603089879e-12, 5.9271020437688792e-12, 
    5.9381335439581406e-12, 5.9419746194582035e-12,
  // Sqw-Na(6, 0-1999)
    0.027516676840134143, 0.027513822430412459, 0.027505200402471862, 
    0.027490638019522274, 0.027469859183997653, 0.027442500792331927, 
    0.02740813316809761, 0.027366282577290391, 0.027316453828049057, 
    0.027258151231005709, 0.027190896677390997, 0.027114244178465866, 
    0.02702779078854161, 0.02693118430289132, 0.026824128410827767, 
    0.026706386066766199, 0.026577781738629635, 0.026438202962928658, 
    0.02628760136155681, 0.026125993041179556, 0.025953458168101406, 
    0.025770139521955428, 0.025576239972151867, 0.025372019046041021, 
    0.025157788996251464, 0.024933910948806374, 0.024700791758318151, 
    0.024458882076279574, 0.024208675856895168, 0.023950711125705713, 
    0.023685571394797426, 0.023413886716438768, 0.023136333113956215, 
    0.02285362908341881, 0.022566528056420974, 0.02227580614518785, 
    0.021982245107066638, 0.021686611183059229, 0.021389631180486791, 
    0.02109196777455814, 0.020794196400540577, 0.020496786226166099, 
    0.020200087497629065, 0.019904327048135297, 0.019609612992852649, 
    0.019315948691832997, 0.019023255053143326, 0.01873139929556621, 
    0.018440227515527503, 0.018149597910407829, 0.017859411372055489, 
    0.017569636408814909, 0.017280325961142401, 0.016991624575619767, 
    0.016703765484457171, 0.016417058264993799, 0.016131868780796643, 
    0.015848593900289847, 0.015567633950845173, 0.015289365944309295, 
    0.015014120308194949, 0.014742163233859825, 0.014473685911939491, 
    0.014208800996100633, 0.013947545754361457, 0.013689890652110872, 
    0.013435751647568148, 0.013185004308105722, 0.012937497965452736, 
    0.012693068467295763, 0.012451548570018442, 0.012212775556715317, 
    0.01197659616472516, 0.011742869295352306, 0.011511467211573635, 
    0.011282275995995574, 0.011055195959123479, 0.010830142496747252, 
    0.010607047645675778, 0.010385862330331978, 0.010166559071558116, 
    0.0099491347721719758, 0.0097336131145054211, 0.0095200461025724877, 
    0.0093085143448290632, 0.0090991257865656941, 0.0088920127464593886, 
    0.0086873272737897911, 0.0084852350076880297, 0.0082859078756223684, 
    0.0080895161036464002, 0.0078962201136213526, 0.0077061629398768091, 
    0.0075194637974733804, 0.0073362133674846662, 0.0071564712290610169, 
    0.0069802656701978627, 0.0068075958664944054, 0.0066384361570890095, 
    0.0064727419036561115, 0.0063104562278798798, 0.0061515168167453546, 
    0.0059958619841833346, 0.0058434352875555854, 0.0056941882060904279, 
    0.0055480806671265922, 0.0054050795140878488, 0.0052651553011551864, 
    0.0051282780296242553, 0.0049944125758450662, 0.004863514581993386, 
    0.004735527488787839, 0.0046103812016763364, 0.0044879926312625324, 
    0.0043682680753101425, 0.0042511071550769448, 0.0041364078187079295, 
    0.0040240718035726014, 0.0039140099183246832, 0.0038061465603681345, 
    0.0037004230094519683, 0.003596799209192167, 0.0034952539378254239, 
    0.0033957834509472378, 0.0032983988306989676, 0.0032031223833241121, 
    0.0031099834836568578, 0.0030190142718151173, 0.0029302455709343334, 
    0.0028437033258845753, 0.0027594057740311872, 0.0026773614626775179, 
    0.0025975681349092801, 0.0025200124249570117, 0.0024446702420727055, 
    0.002371507681770892, 0.0023004822860608542, 0.0022315444786901381, 
    0.0021646390241794738, 0.0020997063957613493, 0.002036683981350265, 
    0.0019755071019670373, 0.0019161098573559042, 0.0018584258435105688, 
    0.001802388802707718, 0.0017479332668731433, 0.0016949952406114966, 
    0.0016435129443991164, 0.0015934276066148704, 0.0015446842617271922, 
    0.0014972324875113668, 0.0014510270018962673, 0.001406028042963582, 
    0.0013622014739132313, 0.0013195185856478872, 0.0012779556076968684, 
    0.0012374929766462927, 0.0011981144430180926, 0.0011598061167613838, 
    0.0011225555546387992, 0.0010863509792803658, 0.0010511806921323595, 
    0.0010170327061094131, 0.00098389458517264029, 0.00095175344422092779, 
    0.0009205960394189878, 0.00089040887005374268, 0.00086117821913266632, 
    0.00083289007935342647, 0.00080552993965126297, 0.00077908243973984757, 
    0.00075353093007225758, 0.00072885699736879167, 0.0007050400277753405, 
    0.00068205687936312106, 0.00065988172372519432, 0.00063848609536145762, 
    0.00061783916113448837, 0.00059790819462096287, 0.0005786592157909767, 
    0.00056005773841339107, 0.00054206955796567416, 0.00052466151223887713, 
    0.00050780215451513659, 0.00049146229327126341, 0.00047561537023242309, 
    0.00046023766742257723, 0.00044530835101869425, 0.00043080937329504178, 
    0.00041672526257288526, 0.00040304283461335081, 0.00038975085788839489, 
    0.00037683970082246822, 0.00036430098291400411, 0.00035212724510024699, 
    0.00034031164901615933, 0.00032884771063456357, 0.00031772907134793076, 
    0.00030694930856752807, 0.00029650178776139237, 0.00028637955779729004, 
    0.00027657529086940385, 0.00026708126679471546, 0.0002578893990500066, 
    0.00024899129690840032, 0.00024037835501291592, 0.00023204185938024093, 
    0.00022397309777856449, 0.00021616346304570674, 0.00020860454024445284, 
    0.00020128817224666324, 0.00019420650273528574, 0.00018735199985883054, 
    0.00018071746700635665, 0.00017429604870919507, 0.00016808123918035775, 
    0.00016206689856114364, 0.0001562472780789118, 0.00015061705088021866, 
    0.00014517134130500949, 0.00013990574276535837, 0.00013481631388166814, 
    0.00012989954437658894, 0.00012515228620879008, 0.00012057165085710432, 
    0.00011615487953034284, 0.00011189919824376356, 0.00010780167314912027, 
    0.00010385908252593076, 0.00010006782019682067, 9.6423841080229628e-05, 
    9.2922653851284235e-05, 8.9559359252994663e-05, 8.6328726593176445e-05, 
    8.3225296366482723e-05, 8.0243494452854268e-05, 7.7377743248573338e-05, 
    7.4622557237737322e-05, 7.1972614381043431e-05, 6.9422799505880107e-05, 
    6.6968220748527761e-05, 6.460420422221525e-05, 6.2326274860148923e-05, 
    6.0130132500835447e-05, 5.8011631742491108e-05, 5.5966772174468619e-05, 
    5.3991702770559403e-05, 5.2082741072979357e-05, 5.0236404859004277e-05, 
    4.8449451715587119e-05, 4.6718920629990538e-05, 4.5042169429884138e-05, 
    4.3416902583674873e-05, 4.1841185276135452e-05, 4.0313441494986605e-05, 
    3.883243577733722e-05, 3.7397239980750063e-05, 3.6007187757441433e-05, 
    3.4661820213121752e-05, 3.3360826521795713e-05, 3.2103983120855145e-05, 
    3.0891094660842552e-05, 2.9721939279104208e-05, 2.8596220142955245e-05, 
    2.7513524659623715e-05, 2.6473292323576446e-05, 2.5474791858992691e-05, 
    2.4517108074735555e-05, 2.3599138618191587e-05, 2.2719600537653284e-05, 
    2.1877046204438974e-05, 2.1069887707246823e-05, 2.0296428345251769e-05, 
    1.9554899377829972e-05, 1.8843499809937679e-05, 1.8160436775277417e-05, 
    1.7503964069447959e-05, 1.6872416599671119e-05, 1.6264238932166416e-05, 
    1.5678006681657097e-05, 1.5112440123292753e-05, 1.4566410037511336e-05, 
    1.4038936349941712e-05, 1.3529180552191484e-05, 1.3036433159643313e-05, 
    1.2560097582593905e-05, 1.2099671778495767e-05, 1.165472895185626e-05, 
    1.1224898409603555e-05, 1.0809847495598433e-05, 1.0409265337078946e-05, 
    1.0022848948902155e-05, 9.6502920572353592e-06, 9.2912768224725185e-06, 
    8.9454684587887248e-06, 8.6125125717583309e-06, 8.2920348754511034e-06, 
    7.9836428240031489e-06, 7.6869286149759936e-06, 7.4014730065795822e-06, 
    7.1268494395686534e-06, 6.8626280613281264e-06, 6.6083793934024959e-06, 
    6.363677540426703e-06, 6.1281029770333637e-06, 5.9012450475370688e-06, 
    5.6827043531309503e-06, 5.4720951817148017e-06, 5.2690480644833074e-06, 
    5.0732124423549e-06, 4.8842593186317841e-06, 4.7018836889296796e-06, 
    4.5258064937676385e-06, 4.3557758451073659e-06, 4.191567333112252e-06, 
    4.0329833138000236e-06, 3.8798511918843096e-06, 3.7320208264819376e-06, 
    3.5893612788159907e-06, 3.4517571784500837e-06, 3.3191049993358e-06, 
    3.1913095125845121e-06, 3.0682806257071635e-06, 2.9499307424052301e-06, 
    2.8361726949946029e-06, 2.7269182272141831e-06, 2.6220769461562194e-06, 
    2.5215556248660095e-06, 2.4252577214304398e-06, 2.3330829855354182e-06, 
    2.2449270442312694e-06, 2.1606808919408873e-06, 2.080230249534177e-06, 
    2.0034548011239974e-06, 1.9302273596366139e-06, 1.8604130510210365e-06, 
    1.7938686367430773e-06, 1.7304421124321991e-06, 1.6699727221258996e-06, 
    1.6122915115632071e-06, 1.5572225082203935e-06, 1.504584564094591e-06, 
    1.4541938328533627e-06, 1.4058667847615165e-06, 1.3594235984305036e-06, 
    1.314691717919104e-06, 1.2715093335580002e-06, 1.22972854091696e-06, 
    1.1892179540661561e-06, 1.1498645954327775e-06, 1.1115749469027125e-06, 
    1.0742751186831706e-06, 1.0379101627799535e-06, 1.0024426201243033e-06, 
    9.6785043684851109e-07, 9.3412441420713706e-07, 9.012653669971455e-07, 
    8.6928116103571709e-07, 8.3818378441663943e-07, 8.0798658617606435e-07, 
    7.7870179250313164e-07, 7.5033838902543954e-07, 7.2290043754515103e-07, 
    6.9638587753952804e-07, 6.7078584378622201e-07, 6.4608451079808606e-07, 
    6.2225944992429456e-07, 5.99282457220987e-07, 5.7712078009411705e-07, 
    5.5573864272289955e-07, 5.3509894727402549e-07, 5.1516501513882743e-07, 
    4.959022316297199e-07, 4.7727947115694868e-07, 4.5927020516729982e-07, 
    4.4185323025371069e-07, 4.2501299218730833e-07, 4.0873951905827565e-07, 
    3.9302800675729435e-07, 3.778781204402187e-07, 3.6329308375430548e-07, 
    3.4927862584082166e-07, 3.358418463499309e-07, 3.2299004636938823e-07, 
    3.1072956152132853e-07, 2.9906462728576608e-07, 2.8799630619017222e-07, 
    2.7752151279829059e-07, 2.6763218162568031e-07, 2.583146325664949e-07, 
    2.4954919257169228e-07, 2.4131012874328324e-07, 2.3356593323708215e-07, 
    2.2627997587897932e-07, 2.1941150733279402e-07, 2.1291695968187326e-07, 
    2.067514569330815e-07, 2.0087042208437662e-07, 1.952311536698032e-07, 
    1.8979424690745795e-07, 1.8452475199171199e-07, 1.7939299315469e-07, 
    1.743750112394422e-07, 1.6945263469108264e-07, 1.6461322163955895e-07, 
    1.5984914475155151e-07, 1.5515710610197094e-07, 1.5053737113501551e-07, 
    1.459929991495717e-07, 1.4152912715983579e-07, 1.3715233783961986e-07, 
    1.3287011739950695e-07, 1.2869038870165443e-07, 1.246210933411389e-07, 
    1.2066979417759261e-07, 1.1684327706801667e-07, 1.1314714418287709e-07, 
    1.0958540860932801e-07, 1.0616011602237429e-07, 1.0287103150344879e-07, 
    9.9715434211575267e-08, 9.6688059728919617e-08, 9.3781218430683479e-08, 
    9.0985101176246274e-08, 8.8288262649909349e-08, 8.5678251938019776e-08, 
    8.3142341763506483e-08, 8.0668295712643086e-08, 7.8245107300891806e-08, 
    7.5863647637210154e-08, 7.3517167803877961e-08, 7.120161756998523e-08, 
    6.8915760400044896e-08, 6.666108457179023e-08, 6.4441528135639539e-08, 
    6.2263050771811474e-08, 6.0133095709842131e-08, 5.8059990505702342e-08, 
    5.6052335357388415e-08, 5.4118423619280294e-08, 5.226573105191458e-08, 
    5.0500500591088002e-08, 4.8827437961962998e-08, 4.7249523002908506e-08, 
    4.5767931672050669e-08, 4.4382056606719633e-08, 4.308960893771311e-08, 
    4.1886782252254538e-08, 4.0768459743362827e-08, 3.9728448269943081e-08, 
    3.8759726537662981e-08, 3.7854698888092406e-08, 3.700544948457444e-08, 
    3.6203994236518012e-08, 3.5442528111974358e-08, 3.4713664650710491e-08, 
    3.4010661746038787e-08, 3.3327624919651118e-08, 3.2659676229923003e-08, 
    3.2003075676653315e-08, 3.1355282142449186e-08, 3.0714943958375467e-08, 
    3.0081814161902014e-08, 2.9456592631787912e-08, 2.8840704768922823e-08, 
    2.8236034091473745e-08, 2.7644631540768401e-08, 2.7068427934751575e-08, 
    2.6508975778013749e-08, 2.5967243844573278e-08, 2.5443481700977861e-08, 
    2.4937163668052655e-08, 2.4447012680815309e-08, 2.3971096259212901e-08, 
    2.3506979537696829e-08, 2.3051915785947247e-08, 2.2603052528678526e-08, 
    2.2157632302880024e-08, 2.1713169817408961e-08, 2.126759232321532e-08, 
    2.0819335292569005e-08, 2.0367391470737537e-08, 1.9911316050354531e-08, 
    1.9451194757648186e-08, 1.898758361259947e-08, 1.8521430175375352e-08, 
    1.8053985255313372e-08, 1.7586712802994994e-08, 1.7121203428785045e-08, 
    1.6659095165996469e-08, 1.620200298014966e-08, 1.5751457546954234e-08, 
    1.5308852862334291e-08, 1.487540250280554e-08, 1.4452104517716888e-08, 
    1.4039715849299927e-08, 1.3638737570285133e-08, 1.324941295001953e-08, 
    1.287174004513123e-08, 1.2505500232320634e-08, 1.2150302834268538e-08, 
    1.1805644737959187e-08, 1.1470981965633777e-08, 1.1145808757419495e-08, 
    1.0829737980546981e-08, 1.0522576106683393e-08, 1.0224385441213493e-08, 
    9.9355270584923898e-09, 9.6566789535297611e-09, 9.388826085424586e-09, 
    9.1332211193344873e-09, 8.8913175153416778e-09, 8.6646788716735659e-09, 
    8.4548708477516549e-09, 8.2633433212186017e-09, 8.0913115113640516e-09, 
    7.9396445995780596e-09, 7.8087699125481133e-09, 7.6985990973862528e-09, 
    7.6084811562691404e-09, 7.5371849193552084e-09, 7.4829117761512529e-09, 
    7.4433374143393282e-09, 7.4156800836231521e-09, 7.3967916275108093e-09, 
    7.3832670390991961e-09, 7.3715676914342727e-09, 7.3581533929572574e-09, 
    7.3396180466732745e-09, 7.3128237245362324e-09, 7.2750275496659525e-09, 
    7.2239957291255531e-09, 7.1580987820611478e-09, 7.0763823448838063e-09, 
    6.9786082190654072e-09, 6.8652616653771747e-09, 6.737522294618116e-09, 
    6.5971983574015987e-09, 6.4466265148121626e-09, 6.2885421731091852e-09, 
    6.1259277666666445e-09, 5.9618487427568009e-09, 5.7992880957782608e-09, 
    5.6409909693454627e-09, 5.4893299085226558e-09, 5.3461998594729042e-09, 
    5.2129492030838712e-09, 5.0903502291001068e-09, 4.9786087590947305e-09, 
    4.8774096592840596e-09, 4.7859919747820678e-09, 4.7032456950707866e-09, 
    4.6278208919859451e-09, 4.55824006449209e-09, 4.4930052199332761e-09, 
    4.4306928542252789e-09, 4.3700317896897973e-09, 4.3099611144819616e-09, 
    4.2496673045154861e-09, 4.1886014728823567e-09, 4.1264787665999569e-09, 
    4.063262921180527e-09, 3.9991390895453036e-09, 3.9344782203631246e-09, 
    3.8697957965360624e-09, 3.8057075845429736e-09, 3.7428844684888321e-09, 
    3.6820083044789614e-09, 3.6237303924200713e-09, 3.5686342084342425e-09, 
    3.5172037576912574e-09, 3.4697990210779085e-09, 3.4266395470549818e-09, 
    3.3877971345484652e-09, 3.3531978845968222e-09, 3.3226334864572001e-09, 
    3.2957807805286542e-09, 3.2722281335680458e-09, 3.2515063785194613e-09, 
    3.2331218656252419e-09, 3.2165887321465828e-09, 3.2014577539486587e-09, 
    3.1873392913589753e-09, 3.1739185928920871e-09, 3.1609622862945831e-09, 
    3.1483159797701985e-09, 3.1358935679693274e-09, 3.1236598725573132e-09, 
    3.1116086789405116e-09, 3.0997388653719605e-09, 3.0880312422880853e-09, 
    3.0764287877149459e-09, 3.0648223458725413e-09, 3.0530434268098777e-09, 
    3.0408647719900838e-09, 3.0280087097443139e-09, 3.0141623241281965e-09, 
    2.9989979673887115e-09, 2.9821969099831247e-09, 2.9634739162107596e-09, 
    2.9426002236501635e-09, 2.9194228996355413e-09, 2.8938787502836592e-09, 
    2.866001722564817e-09, 2.8359232284425529e-09, 2.8038656367942125e-09, 
    2.7701296033475905e-09, 2.7350765375962035e-09, 2.6991076223891329e-09, 
    2.6626411755600201e-09, 2.6260898982551183e-09, 2.5898396313115764e-09, 
    2.5542308253335118e-09, 2.5195438212810797e-09, 2.4859885433649522e-09, 
    2.4536990612846895e-09, 2.4227329755649537e-09, 2.3930754896976139e-09, 
    2.3646475788738152e-09, 2.3373176052474795e-09, 2.3109154088020623e-09, 
    2.2852479117005875e-09, 2.2601150764164214e-09, 2.2353252459424737e-09, 
    2.2107088165814716e-09, 2.1861295377684539e-09, 2.1614927663061244e-09, 
    2.1367504746594152e-09, 2.1119028362340083e-09, 2.0869967024791452e-09, 
    2.0621212155688919e-09, 2.0374012162857027e-09, 2.012988929090364e-09, 
    1.9890546585870063e-09, 1.9657770226745133e-09, 1.9433333665272998e-09, 
    1.9218907340846075e-09, 1.9015979487672944e-09, 1.8825789578636537e-09, 
    1.864927809926149e-09, 1.848705280244497e-09, 1.8339372343829402e-09, 
    1.8206145886834609e-09, 1.8086947366050441e-09, 1.798104104456567e-09, 
    1.7887416052316802e-09, 1.7804825502385852e-09, 1.7731828330722481e-09, 
    1.7666830108841844e-09, 1.7608122589579377e-09, 1.7553920280191277e-09, 
    1.7502395354616376e-09, 1.7451710638757494e-09, 1.740005296654827e-09, 
    1.7345666648560365e-09, 1.7286888615098822e-09, 1.7222183535031568e-09, 
    1.7150179243045617e-09, 1.7069699513148192e-09, 1.6979793432678867e-09, 
    1.6879757917845905e-09, 1.6769153267613275e-09, 1.664780927058831e-09, 
    1.6515822643226382e-09, 1.637354534253127e-09, 1.622156581097941e-09, 
    1.6060683627482465e-09, 1.5891880739121758e-09, 1.5716289893779616e-09, 
    1.5535163149047304e-09, 1.5349840678068546e-09, 1.5161721909668025e-09, 
    1.497223841558579e-09, 1.4782829497771527e-09, 1.4594919080284443e-09, 
    1.4409894418070476e-09, 1.4229084596560062e-09, 1.4053739430710071e-09, 
    1.3885006872873351e-09, 1.3723910033079219e-09, 1.357132293994969e-09, 
    1.3427946872076005e-09, 1.3294287415022109e-09, 1.3170635162795219e-09, 
    1.30570510429483e-09, 1.2953359117673412e-09, 1.2859147878200813e-09, 
    1.2773782271543206e-09, 1.2696425817075387e-09, 1.2626073747186966e-09, 
    1.2561594625917196e-09, 1.2501779250533803e-09, 1.2445392936980828e-09, 
    1.2391228855921973e-09, 1.2338158081964095e-09, 1.228517416219379e-09, 
    1.223142864519473e-09, 1.217625697133397e-09, 1.2119192583018399e-09, 
    1.2059970394790131e-09, 1.1998519069887186e-09, 1.19349444977447e-09, 
    1.1869504822892356e-09, 1.1802579957422489e-09, 1.1734636223943276e-09, 
    1.1666189147863755e-09, 1.1597764960838218e-09, 1.1529863818824598e-09, 
    1.1462925374093354e-09, 1.1397299346811862e-09, 1.1333221866315572e-09, 
    1.1270799834906612e-09, 1.1210003316271637e-09, 1.1150667746386244e-09, 
    1.1092504842404818e-09, 1.1035122571402799e-09, 1.0978052295929527e-09, 
    1.0920781834275916e-09, 1.0862791635934017e-09, 1.0803592240876665e-09, 
    1.0742759609466207e-09, 1.0679966621825461e-09, 1.0615007385187434e-09, 
    1.054781377012384e-09, 1.0478461713895736e-09, 1.0407167911208455e-09, 
    1.0334275961352396e-09, 1.0260234288000907e-09, 1.0185566286913956e-09, 
    1.0110836162273932e-09, 1.0036612196802861e-09, 9.9634311853923826e-10, 
    9.8917657932322208e-10, 9.8219982158144422e-10, 9.7544009072918337e-10, 
    9.6891263992099835e-10, 9.6262054748567544e-10, 9.5655542402076275e-10, 
    9.5069880987368984e-10, 9.4502418605740859e-10, 9.3949934251706104e-10, 
    9.3408899788308446e-10, 9.2875740130086177e-10, 9.2347085154636895e-10, 
    9.1819987978602345e-10, 9.1292109819938024e-10, 9.0761852746314313e-10, 
    9.0228441479723832e-10, 8.9691943860515876e-10, 8.9153236602466627e-10, 
    8.8613910172161672e-10, 8.8076129242313826e-10, 8.7542447838554255e-10, 
    8.7015603116071278e-10, 8.6498294686073093e-10, 8.5992975059210092e-10, 
    8.5501659507412028e-10, 8.502578001501599e-10, 8.4566083043447572e-10, 
    8.4122588671653498e-10, 8.3694599909981176e-10, 8.3280769084404216e-10, 
    8.2879201157151014e-10, 8.2487592580274983e-10, 8.2103383008400547e-10, 
    8.1723916466899775e-10, 8.1346591508208546e-10, 8.0968999910225325e-10, 
    8.0589040758300096e-10, 8.0205012927181357e-10, 7.9815674756307935e-10, 
    7.9420282550082548e-10, 7.901859751907829e-10, 7.861087140511817e-10, 
    7.8197806922934602e-10, 7.7780500321215995e-10, 7.7360365033790847e-10, 
    7.6939047144473855e-10, 7.651832771557749e-10, 7.6100027945738685e-10, 
    7.5685912674182435e-10, 7.527760419469317e-10, 7.4876503493951872e-10, 
    7.4483727641376245e-10, 7.4100059203922289e-10, 7.3725912769044798e-10, 
    7.33613135951954e-10, 7.3005893445807911e-10, 7.265889399595092e-10, 
    7.2319189238007304e-10, 7.1985316365263185e-10, 7.165552401134183e-10, 
    7.1327832206007791e-10, 7.1000110738193098e-10, 7.0670169138562496e-10, 
    7.033586232627129e-10, 6.9995201061993848e-10, 6.9646469303759467e-10, 
    6.9288332971379317e-10, 6.8919939268460189e-10, 6.8540989449540572e-10, 
    6.8151785424826746e-10, 6.7753234987376692e-10, 6.734681949376379e-10, 
    6.6934516158598246e-10, 6.6518685406783446e-10, 6.610192230916715e-10, 
    6.5686892051927336e-10, 6.5276152712768317e-10, 6.4871989748555982e-10, 
    6.4476269059075941e-10, 6.409032851599611e-10, 6.3714912152827225e-10, 
    6.3350158900982229e-10, 6.2995640487589228e-10, 6.2650451726310578e-10, 
    6.2313334979296727e-10, 6.1982835680015143e-10, 6.1657464201516269e-10, 
    6.1335857388564813e-10, 6.1016915219100334e-10, 6.0699910063175857e-10, 
    6.0384551104818786e-10, 6.0071007718050394e-10, 5.9759883902973047e-10, 
    5.9452156211127558e-10, 5.9149075231719028e-10, 5.8852046307914533e-10, 
    5.8562495738629492e-10, 5.8281738239267531e-10, 5.8010850892424247e-10, 
    5.7750569213253959e-10, 5.7501205267858608e-10, 5.7262601457007406e-10, 
    5.7034113781101853e-10, 5.6814633888258237e-10, 5.6602638638047302e-10, 
    5.6396270335940041e-10, 5.6193434731083271e-10, 5.5991913969373158e-10, 
    5.578947837537294e-10, 5.5583997539329678e-10, 5.5373532906646523e-10, 
    5.5156415151389343e-10, 5.4931293978133419e-10, 5.4697167373359666e-10, 
    5.4453385510347263e-10, 5.4199638808566143e-10, 5.3935929175394367e-10, 
    5.3662537622306296e-10, 5.3379986388875344e-10, 5.308900664266294e-10, 
    5.2790506900391671e-10, 5.2485551444369143e-10, 5.2175337807131264e-10, 
    5.1861180526181901e-10, 5.1544489467037971e-10, 5.1226746688040891e-10, 
    5.090947339712044e-10, 5.0594191891061501e-10, 5.0282378160184964e-10, 
    4.9975412071149124e-10, 4.9674524047951459e-10, 4.9380747559338793e-10, 
    4.9094877619583978e-10, 4.881744394537473e-10, 4.8548695961847664e-10, 
    4.8288608744549487e-10, 4.8036901187679402e-10, 4.7793073653541244e-10, 
    4.7556452823974174e-10, 4.732624746058644e-10, 4.7101603229832163e-10, 
    4.6881659175612651e-10, 4.6665592770748008e-10, 4.6452659292991995e-10, 
    4.6242216245490166e-10, 4.6033738099157898e-10, 4.5826814730025489e-10, 
    4.5621144204971331e-10, 4.5416512072925542e-10, 4.5212770299645392e-10, 
    4.5009808288755031e-10, 4.4807527616757599e-10, 4.4605815776969621e-10, 
    4.4404526656439554e-10, 4.4203461586599995e-10, 4.4002361197233969e-10, 
    4.3800900217238304e-10, 4.3598692398653791e-10, 4.3395299690029261e-10, 
    4.3190251416329075e-10, 4.2983066792891427e-10, 4.2773284869102676e-10, 
    4.256049493487885e-10, 4.2344370544122713e-10, 4.2124696718002302e-10, 
    4.1901396021313187e-10, 4.1674544046841407e-10, 4.1444377724400377e-10, 
    4.1211289510973467e-10, 4.0975815661566721e-10, 4.0738611304391285e-10, 
    4.0500422693117468e-10, 4.026205150697726e-10, 4.0024322018297709e-10, 
    3.9788046948797189e-10, 3.9554000323434776e-10, 3.9322892623678945e-10, 
    3.9095355666617708e-10, 3.8871931599863678e-10, 3.8653070113820091e-10, 
    3.8439129509779434e-10, 3.8230384666960035e-10, 3.8027036493315444e-10, 
    3.7829226603048651e-10, 3.7637051574435846e-10, 3.7450579231101958e-10, 
    3.7269860449684088e-10, 3.7094940533914755e-10, 3.6925860469075001e-10, 
    3.6762655202919521e-10, 3.6605339237178422e-10, 3.64538884378175e-10, 
    3.6308209646773638e-10, 3.6168112392750676e-10, 3.6033275884330747e-10, 
    3.5903224537029854e-10, 3.5777309117611136e-10, 3.5654705834863256e-10, 
    3.5534426393618681e-10, 3.5415348564130623e-10, 3.529625903300052e-10, 
    3.5175910738935005e-10, 3.5053082540497882e-10, 3.4926643721704036e-10, 
    3.4795609282400382e-10, 3.4659186924916066e-10, 3.4516806433588876e-10, 
    3.4368135181648486e-10, 3.4213074147564893e-10, 3.4051742964396968e-10, 
    3.388445119400015e-10, 3.3711667106546159e-10, 3.3533983690192216e-10, 
    3.3352090534192705e-10, 3.3166749587633707e-10, 3.2978781750707359e-10, 
    3.27890585135474e-10, 3.2598501524378073e-10, 3.2408080094144168e-10, 
    3.2218812489730348e-10, 3.2031755019141655e-10, 3.1847989388020039e-10, 
    3.1668595565894086e-10, 3.1494620316902122e-10, 3.1327035450700245e-10, 
    3.1166696575900965e-10, 3.1014301573682459e-10, 3.0870357845255073e-10, 
    3.0735157364290972e-10, 3.0608767337851415e-10, 3.0491031959869525e-10, 
    3.0381588623890114e-10, 3.0279890083145573e-10, 3.0185234575309584e-10, 
    3.0096793827710388e-10, 3.0013640105234217e-10, 2.9934763981843813e-10, 
    2.985908954876786e-10, 2.9785480794016263e-10, 2.9712749893755574e-10, 
    2.9639663764046839e-10, 2.9564960930695042e-10, 2.948737731551761e-10, 
    2.9405686799362796e-10, 2.9318750314087192e-10, 2.9225580714799424e-10, 
    2.9125405691704341e-10, 2.9017733979985033e-10, 2.8902406894411779e-10, 
    2.8779636341218935e-10, 2.8650014692883559e-10, 2.8514501092826254e-10, 
    2.8374376339871111e-10, 2.8231173287239438e-10, 2.8086584504730608e-10, 
    2.7942357851061145e-10, 2.7800183372756825e-10, 2.7661587044488227e-10, 
    2.7527833988785665e-10, 2.7399853751665159e-10, 2.7278186728468195e-10, 
    2.7162962856522543e-10, 2.7053905869900219e-10, 2.6950368633010769e-10, 
    2.6851390494573143e-10, 2.6755778475758362e-10, 2.6662199547485006e-10, 
    2.6569285063194021e-10, 2.6475732549249977e-10, 2.638040568761047e-10, 
    2.6282418498084907e-10, 2.6181205187159672e-10, 2.6076564090373466e-10, 
    2.5968680133472775e-10, 2.5858115280933294e-10, 2.5745778526962259e-10, 
    2.5632866363631483e-10, 2.5520786934620711e-10, 2.5411068057052787e-10, 
    2.530525752617791e-10, 2.5204819812634494e-10, 2.5111040867116318e-10, 
    2.5024939819373456e-10, 2.4947201242069136e-10, 2.4878123534119904e-10, 
    2.4817594101557216e-10, 2.4765085764269725e-10, 2.4719680208212641e-10, 
    2.4680112248332947e-10, 2.4644836021460751e-10, 2.4612105861680377e-10, 
    2.4580070332685703e-10, 2.4546870105569632e-10, 2.4510738441524967e-10, 
    2.4470090900624161e-10, 2.4423607449560374e-10, 2.43702933784308e-10, 
    2.4309522109597546e-10, 2.4241051064686903e-10, 2.4165017252028865e-10, 
    2.4081906025201164e-10, 2.3992504296118138e-10, 2.3897834322753068e-10, 
    2.3799082421438653e-10, 2.3697519900146066e-10, 2.3594430565951659e-10, 
    2.3491042420636833e-10, 2.3388474188923404e-10, 2.328769313714851e-10, 
    2.3189491268742589e-10, 2.3094472337242078e-10, 2.3003054437873921e-10, 
    2.2915478759749229e-10, 2.283182756134704e-10, 2.2752041570005825e-10, 
    2.2675940437804539e-10, 2.2603238000555966e-10, 2.2533557366049373e-10, 
    2.2466438957466013e-10, 2.2401349282535129e-10, 2.2337682981084561e-10, 
    2.2274768123189153e-10, 2.2211868316862671e-10, 2.214818992247478e-10, 
    2.2082889126354046e-10, 2.2015087189512148e-10, 2.1943888646877174e-10, 
    2.1868408874135542e-10, 2.1787805899907971e-10, 2.1701322806305038e-10, 
    2.1608331945905254e-10, 2.1508386129471106e-10, 2.1401267334912438e-10, 
    2.1287033551345937e-10, 2.1166053235431857e-10, 2.1039028243719461e-10, 
    2.0906994378565129e-10, 2.0771301577373788e-10, 2.0633566995550945e-10, 
    2.049560576723346e-10, 2.0359340152284405e-10, 2.0226695140600226e-10, 
    2.0099484669690586e-10, 1.9979304244729665e-10, 1.9867430949206927e-10, 
    1.9764749392270491e-10, 1.9671702005187904e-10, 1.9588274928804709e-10, 
    1.9514015663620554e-10, 1.9448084761614255e-10, 1.9389331210281497e-10, 
    1.9336388512841571e-10, 1.9287777510765259e-10, 1.9242009188018425e-10, 
    1.9197675042995785e-10, 1.9153522543286663e-10, 1.910850219105477e-10, 
    1.9061795449723533e-10, 1.901281480473431e-10, 1.8961186671673247e-10, 
    1.8906716898695641e-10, 1.8849350674476153e-10, 1.8789127478797766e-10, 
    1.8726141645030327e-10, 1.8660507658806585e-10, 1.8592336944668597e-10, 
    1.8521722138242209e-10, 1.8448733911724189e-10, 1.8373423347463086e-10, 
    1.8295833408444577e-10, 1.821601360027217e-10, 1.8134039540390192e-10, 
    1.8050033350312927e-10, 1.7964185635985215e-10, 1.7876774012874392e-10, 
    1.7788180054209952e-10, 1.7698898276243496e-10, 1.7609537374622579e-10, 
    1.7520808337075506e-10, 1.7433501984294863e-10, 1.7348450068608052e-10, 
    1.72664776235673e-10, 1.7188345079908852e-10, 1.7114690371176736e-10, 
    1.7045970837419261e-10, 1.6982420179228246e-10, 1.6924019171212273e-10, 
    1.6870489906714149e-10, 1.6821310657051673e-10, 1.6775754643884531e-10, 
    1.6732943951737934e-10, 1.6691915948100022e-10, 1.6651689871991898e-10, 
    1.6611330371514495e-10, 1.6569996620611986e-10, 1.6526976969958343e-10, 
    1.6481704491162992e-10, 1.6433758250999721e-10, 1.6382852593249178e-10, 
    1.6328822683966839e-10, 1.6271610089013552e-10, 1.6211255666463409e-10, 
    1.6147901487821831e-10, 1.6081801950600095e-10, 1.6013339844369281e-10, 
    1.5943044759530942e-10, 1.5871601887766945e-10, 1.579985026096058e-10, 
    1.5728760136291411e-10, 1.5659390871240104e-10, 1.5592826103222494e-10, 
    1.5530096217449499e-10, 1.5472088570650775e-10, 1.5419463068134638e-10, 
    1.5372577651816386e-10, 1.5331437203107188e-10, 1.5295670519408703e-10, 
    1.5264542343112226e-10, 1.5236997752985839e-10, 1.5211738197056154e-10, 
    1.518731739927548e-10, 1.5162252804352242e-10, 1.5135135810187016e-10, 
    1.5104735120965457e-10, 1.5070079448515623e-10, 1.50305168012415e-10, 
    1.4985742273012853e-10, 1.4935798557198095e-10, 1.4881047453519124e-10, 
    1.4822121104313081e-10, 1.4759854813607442e-10, 1.46952138019897e-10, 
    1.462921499675411e-10, 1.4562855308070073e-10, 1.4497044457718033e-10, 
    1.4432553022589837e-10, 1.4369970591459836e-10, 1.4309680347717539e-10, 
    1.4251846461404528e-10, 1.4196416671442647e-10, 1.4143134992121633e-10, 
    1.4091569097657899e-10, 1.4041144950840217e-10, 1.3991189533403352e-10, 
    1.3940977824722588e-10, 1.3889781032185688e-10, 1.3836911239651214e-10, 
    1.3781761564445509e-10, 1.3723834182941134e-10, 1.3662759531094181e-10, 
    1.3598300676265297e-10, 1.3530347837971919e-10, 1.3458900834459579e-10, 
    1.3384047273765774e-10, 1.3305936596611022e-10, 1.32247582139472e-10, 
    1.3140724257188973e-10, 1.3054062545217967e-10, 1.2965020057040581e-10, 
    1.2873877081762519e-10, 1.2780968617949518e-10, 1.2686713519400558e-10, 
    1.2591639928284527e-10, 1.2496411029243035e-10, 1.2401837234989212e-10, 
    1.2308878974894934e-10, 1.2218629896285978e-10, 1.2132286322717774e-10, 
    1.2051097765915712e-10, 1.1976306466203338e-10, 1.1909074217296378e-10, 
    1.1850408925403413e-10, 1.1801091021467098e-10, 1.1761611653243177e-10, 
    1.1732123979146493e-10, 1.1712418441846358e-10, 1.1701918872937348e-10, 
    1.1699708276439853e-10, 1.1704574592823816e-10, 1.1715081345296607e-10, 
    1.1729649977716604e-10, 1.1746652732647865e-10, 1.1764501700519109e-10, 
    1.1781733055994087e-10, 1.1797072516903542e-10, 1.1809484034551224e-10, 
    1.1818192920872786e-10, 1.1822689740814131e-10, 1.1822711144906972e-10, 
    1.1818209375546867e-10, 1.1809308678425445e-10, 1.1796261393540432e-10, 
    1.1779403139358476e-10, 1.1759117046608693e-10, 1.1735801675886254e-10, 
    1.1709851984115244e-10, 1.1681642823018826e-10, 1.1651521833604576e-10, 
    1.1619799851214123e-10, 1.1586745308514883e-10, 1.1552572478570129e-10, 
    1.1517430795723318e-10, 1.1481390178482166e-10, 1.1444429554093177e-10, 
    1.1406425459907042e-10, 1.1367152302430597e-10, 1.1326287721833678e-10, 
    1.1283433505023834e-10, 1.1238145310408678e-10, 1.1189976085490552e-10, 
    1.1138524058143035e-10, 1.1083487318264203e-10, 1.1024713456915855e-10, 
    1.0962245018363396e-10, 1.0896347688428501e-10, 1.0827527424515384e-10, 
    1.0756522455245006e-10, 1.0684280072589075e-10, 1.0611911668277434e-10, 
    1.054063601164975e-10, 1.0471708202253706e-10, 1.0406349327442565e-10, 
    1.0345672000245266e-10, 1.0290620096595897e-10, 1.0241914725289585e-10, 
    1.0200021266396621e-10, 1.0165130614879756e-10, 1.0137162806925915e-10, 
    1.0115782495674722e-10, 1.0100434470389282e-10, 1.0090383656803222e-10, 
    1.0084767089097336e-10, 1.0082642715358402e-10, 1.0083040606411033e-10, 
    1.0085003062841162e-10, 1.0087622387374092e-10, 1.0090061920664291e-10, 
    1.0091572633432724e-10, 1.0091495707130806e-10, 1.0089260728120427e-10, 
    1.0084374326266662e-10, 1.0076411967826333e-10, 1.0065003249914352e-10, 
    1.0049827606876297e-10, 1.0030609760764855e-10, 1.000712615135935e-10, 
    9.9792136403605465e-11, 9.9467877512573028e-11, 9.9098611800849313e-11, 
    9.8685661594340818e-11, 9.8231713234407948e-11, 9.7740984291280113e-11, 
    9.7219257192070775e-11, 9.6673884743199311e-11, 9.6113640852760629e-11, 
    9.554852119867639e-11, 9.4989406822809137e-11, 9.4447697063836296e-11, 
    9.3934839166428714e-11, 9.34618659545328e-11, 9.303887969089656e-11, 
    9.2674594411527839e-11, 9.2375848373227927e-11, 9.2147237134026835e-11, 
    9.1990771843486471e-11, 9.1905682834339458e-11, 9.1888310217858421e-11, 
    9.1932179132707814e-11, 9.202817851767421e-11, 9.2164958212352606e-11, 
    9.2329422599519888e-11, 9.2507411653857436e-11, 9.268442451634973e-11, 
    9.284644188768368e-11, 9.2980704669649433e-11, 9.3076461250361563e-11, 
    9.3125552943578273e-11, 9.3122866971859734e-11, 9.3066536398703303e-11, 
    9.2957961672162714e-11, 9.2801558622059996e-11, 9.2604352725456319e-11, 
    9.2375379650165044e-11, 9.2125015660940025e-11, 9.1864214332978579e-11, 
    9.1603801388954673e-11, 9.1353788594368357e-11, 9.1122822802083996e-11, 
    9.0917722666962266e-11, 9.0743199470017769e-11, 9.0601667314350452e-11, 
    9.0493238896474512e-11, 9.041580079396983e-11, 9.0365241181295456e-11, 
    9.0335719865858091e-11, 9.0320063739063746e-11, 9.0310188009898949e-11, 
    9.0297597876207494e-11, 9.0273860131007348e-11, 9.0231123155245196e-11, 
    9.0162555454162931e-11, 9.0062756262071121e-11, 8.9928019954893571e-11, 
    8.9756516707091592e-11, 8.9548284937836526e-11, 8.930510257668542e-11, 
    8.903017927944385e-11, 8.8727756125161743e-11, 8.8402592148195517e-11, 
    8.8059442571579004e-11, 8.7702526355991306e-11, 8.7335102826796447e-11, 
    8.6959140558728538e-11, 8.6575182843317598e-11, 8.6182366632007892e-11, 
    8.5778660159828266e-11, 8.5361227385497722e-11, 8.4926955335083749e-11, 
    8.4473017356787462e-11, 8.3997488058912881e-11, 8.3499833666310149e-11, 
    8.2981330435693916e-11, 8.2445271149054083e-11, 8.1896995902113702e-11, 
    8.134364415031531e-11, 8.0793758378718954e-11, 8.0256671589692109e-11, 
    7.9741825126622392e-11, 7.9257994874229158e-11, 7.8812610993637377e-11, 
    7.8411152637561008e-11, 7.8056757484473631e-11, 7.7750037403872593e-11, 
    7.748918052381485e-11, 7.7270266746241087e-11, 7.708784533692813e-11, 
    7.6935640061674714e-11, 7.6807383427406923e-11, 7.6697624003515171e-11, 
    7.6602488821479129e-11, 7.6520259838319012e-11, 7.6451761127607415e-11, 
    7.6400450902997109e-11, 7.6372269206640705e-11, 7.6375178470695166e-11, 
    7.6418500697603021e-11, 7.6512031958149507e-11, 7.6665078818778042e-11, 
    7.6885426204033225e-11, 7.7178393554913954e-11, 7.7545978455406856e-11, 
    7.7986242595944052e-11, 7.8492936033549742e-11, 7.9055442164869932e-11, 
    7.9659015467396989e-11, 8.02853552734701e-11, 8.0913432005705529e-11, 
    8.1520564738898349e-11, 8.2083623163084894e-11, 8.258032967541974e-11, 
    8.2990498058954021e-11, 8.3297201651297192e-11, 8.3487702025043984e-11, 
    8.3554155081426405e-11, 8.3493961778111502e-11, 8.3309826343686317e-11, 
    8.3009440633631238e-11, 8.2604898673004461e-11, 8.2111813399806137e-11, 
    8.1548279521641369e-11, 8.0933700676440713e-11, 8.0287618871160497e-11, 
    7.9628574331767802e-11, 7.897315066357293e-11, 7.833519121024051e-11, 
    7.7725294118388232e-11, 7.7150571647905513e-11, 7.6614706770886458e-11, 
    7.6118221197680028e-11, 7.5658987969155932e-11, 7.5232862557757127e-11, 
    7.4834407813986635e-11, 7.4457588982602897e-11, 7.4096441743765692e-11, 
    7.3745593657410877e-11, 7.3400666411235979e-11, 7.3058489348755545e-11, 
    7.2717191046584456e-11, 7.2376129963794759e-11, 7.2035772521706515e-11, 
    7.1697485211803923e-11, 7.1363344405406573e-11, 7.1035958191618625e-11, 
    7.0718348329737927e-11, 7.041385460581132e-11, 7.0126111327403248e-11, 
    6.9859031837237689e-11, 6.9616798097777441e-11, 6.9403807209061377e-11, 
    6.922458528784656e-11, 6.9083599585031668e-11, 6.898501815098651e-11, 
    6.8932397522490542e-11, 6.8928339763991412e-11, 6.8974109539251264e-11, 
    6.9069318062875272e-11, 6.9211652780054256e-11, 6.9396743771818087e-11, 
    6.9618134805878602e-11, 6.9867432304313638e-11, 7.0134602530939901e-11, 
    7.0408412949377258e-11, 7.0676964975931973e-11, 7.0928326198664573e-11, 
    7.1151158132861056e-11, 7.1335352234555568e-11, 7.1472556131496943e-11, 
    7.1556635574694405e-11, 7.1583962177404999e-11, 7.1553575411667722e-11, 
    7.146716458052836e-11, 7.1328919514486376e-11, 7.1145199553484845e-11, 
    7.092412192769971e-11, 7.0675005985930428e-11, 7.0407780281359724e-11, 
    7.0132318033584904e-11, 6.9857778487130089e-11, 6.9591971180268023e-11, 
    6.9340797115206217e-11, 6.9107774321700287e-11, 6.8893742434632976e-11, 
    6.8696717771841032e-11, 6.8511986379197752e-11, 6.8332367360902508e-11, 
    6.8148724433805998e-11, 6.7950627376557187e-11, 6.7727173206729856e-11, 
    6.7467853398034718e-11, 6.7163448258966821e-11, 6.6806822566368731e-11, 
    6.6393598121135171e-11, 6.5922579785407306e-11, 6.5395961965426885e-11, 
    6.4819225690594121e-11, 6.420079537992745e-11, 6.3551424587153424e-11, 
    6.2883422460598494e-11, 6.2209749154742087e-11, 6.1543095759375117e-11, 
    6.08950027874514e-11, 6.027512604596794e-11, 5.9690679311292829e-11, 
    5.9146130528644628e-11, 5.8643132198262943e-11, 5.8180734016364893e-11, 
    5.7755766186026937e-11, 5.736342869794089e-11, 5.6997968955863899e-11, 
    5.6653407906795094e-11, 5.6324206151378928e-11, 5.600587264546936e-11, 
    5.5695401776068638e-11, 5.5391559139154059e-11, 5.5094957918002148e-11, 
    5.480798504399381e-11, 5.4534517859561846e-11, 5.427954919947634e-11, 
    5.4048692364567549e-11, 5.384765553076794e-11, 5.3681681531520144e-11, 
    5.3555051541129194e-11, 5.3470624182224169e-11, 5.3429490901266805e-11, 
    5.3430727541326938e-11, 5.3471288333497953e-11, 5.3546007786248375e-11, 
    5.3647762895464292e-11, 5.3767732617961369e-11, 5.389579844596781e-11, 
    5.4021025576011525e-11, 5.4132240624847096e-11, 5.4218638258318033e-11, 
    5.4270439531099188e-11, 5.4279503531889771e-11, 5.4239906596504408e-11, 
    5.4148414090759482e-11, 5.4004833040628513e-11, 5.3812173952783995e-11, 
    5.3576652233501174e-11, 5.3307461553464618e-11, 5.3016364634856916e-11, 
    5.2717075622363376e-11, 5.2424502041881039e-11, 5.215385159651606e-11, 
    5.1919696291285681e-11, 5.1735012339168618e-11, 5.1610301958367803e-11, 
    5.1552829086326375e-11, 5.1566058728220836e-11, 5.1649319814364481e-11, 
    5.179775040711295e-11, 5.2002537151914749e-11, 5.2251445687868076e-11, 
    5.2529591200693237e-11, 5.2820441076908805e-11, 5.3106934083945305e-11, 
    5.3372666451412313e-11, 5.3603009555979955e-11, 5.3786097384063252e-11, 
    5.3913572778592183e-11, 5.3981045345021072e-11, 5.3988190507386249e-11, 
    5.3938514185096201e-11, 5.3838789339052483e-11, 5.3698228052425587e-11, 
    5.3527467620560369e-11, 5.3337499490514663e-11, 5.3138604029353912e-11, 
    5.2939450681615636e-11, 5.2746408539158501e-11, 5.2563157824840871e-11, 
    5.2390601256532849e-11, 5.2227103246999942e-11, 5.2068984097340995e-11, 
    5.191121579487821e-11, 5.1748238474920275e-11, 5.1574784856756337e-11, 
    5.1386623176384438e-11, 5.1181159125819123e-11, 5.0957806267163781e-11, 
    5.0718125588303173e-11, 5.046571692717132e-11, 5.0205901766840908e-11, 
    4.9945223326723496e-11, 4.9690862099451775e-11, 4.9450000415371305e-11, 
    4.922922259755754e-11, 4.9034009705320169e-11, 4.886836321799609e-11, 
    4.8734567200516473e-11, 4.8633133293733681e-11, 4.8562881408311473e-11, 
    4.8521170404127471e-11, 4.8504206832127268e-11, 4.8507447349025307e-11, 
    4.8526030882097807e-11, 4.8555214476444525e-11, 4.8590790075870848e-11, 
    4.8629442661530947e-11, 4.8669041761694185e-11, 4.8708834717335853e-11, 
    4.8749515445912961e-11, 4.8793178420322393e-11, 4.8843139389266226e-11, 
    4.8903633466031874e-11, 4.8979405462846586e-11, 4.9075225894817022e-11, 
    4.9195372386868255e-11, 4.9343122852572402e-11, 4.9520299891143981e-11, 
    4.9726929869383339e-11, 4.9961040336243782e-11, 5.0218611867988335e-11, 
    5.0493712938468357e-11, 5.0778781363916222e-11, 5.106502080425249e-11, 
    5.1342899723901452e-11, 5.1602678313775769e-11, 5.1834929398908812e-11, 
    5.203101195558178e-11, 5.2183470398912323e-11, 5.2286337354260298e-11, 
    5.2335345042805277e-11, 5.2328046479011554e-11, 5.2263867386445165e-11, 
    5.2144102372164064e-11, 5.197187225718636e-11, 5.1752057688499266e-11, 
    5.1491200380406498e-11, 5.1197385327463742e-11, 5.0880084158230713e-11, 
    5.0549939151493373e-11, 5.0218485825511433e-11, 4.9897815483130801e-11, 
    4.9600148609336824e-11, 4.9337343794787469e-11, 4.9120351575290374e-11, 
    4.8958662206459733e-11, 4.8859735747414302e-11, 4.8828502642840494e-11, 
    4.8866944466276498e-11, 4.8973790994482664e-11, 4.9144382393817963e-11, 
    4.9370714267383055e-11, 4.9641653612109647e-11, 4.9943365479755716e-11, 
    5.0259893995678408e-11, 5.0573897210734356e-11, 5.0867473208753086e-11, 
    5.1123065646377651e-11, 5.1324349695301437e-11, 5.145706379962521e-11, 
    5.150973502727537e-11, 5.147424637832832e-11, 5.1346196255611705e-11, 
    5.1125051855218954e-11, 5.0814055515169519e-11, 5.0419940666340367e-11, 
    4.9952442448742762e-11, 4.9423667103561907e-11, 4.8847362873611728e-11, 
    4.823816347970868e-11, 4.7610828105740376e-11, 4.6979553724093348e-11, 
    4.6357375031174413e-11, 4.5755701239593303e-11, 4.518397518921478e-11, 
    4.4649475486238235e-11, 4.415724240450859e-11, 4.3710116722478875e-11, 
    4.3308871379015899e-11, 4.295241851636133e-11, 4.2638059739152703e-11, 
    4.2361795158179356e-11, 4.2118626876997152e-11, 4.1902888709599524e-11, 
    4.1708560316201169e-11, 4.1529554507355667e-11, 4.1359974745783576e-11, 
    4.1194325965413716e-11, 4.1027645717587508e-11, 4.0855600929830439e-11, 
    4.0674491655784745e-11, 4.0481198302216039e-11, 4.027308158791994e-11, 
    4.0047854114423922e-11, 3.9803438380826983e-11, 3.9537837559488977e-11, 
    3.9249050462009447e-11, 3.8935034805319598e-11, 3.8593730301584662e-11, 
    3.8223170311694534e-11, 3.782163222890656e-11, 3.7387841314137199e-11, 
    3.6921210974290898e-11, 3.64220679558982e-11, 3.5891868369794961e-11, 
    3.5333370213568388e-11, 3.4750738988769766e-11, 3.4149586492684735e-11, 
    3.3536931942220847e-11, 3.29210857827566e-11, 3.2311464838345672e-11, 
    3.171834632876516e-11, 3.1152571726325655e-11, 3.0625212114385188e-11, 
    3.0147208323164206e-11, 2.9729003762323116e-11, 2.938016753330612e-11, 
    2.9109039121243512e-11, 2.8922389938045715e-11, 2.8825138645627057e-11, 
    2.8820108352872233e-11, 2.8907872823705814e-11, 2.908667921703789e-11, 
    2.9352464160001793e-11, 2.9698992496337866e-11, 3.0118075939135917e-11, 
    3.059990938820263e-11, 3.1133466674974873e-11, 3.1706964952517408e-11, 
    3.2308343152907486e-11, 3.2925738505492791e-11, 3.3547902535111669e-11, 
    3.4164537696746021e-11, 3.4766541186364716e-11, 3.5346107019025123e-11, 
    3.5896704482675485e-11, 3.6412943183603684e-11, 3.6890345691855293e-11, 
    3.732506490597709e-11, 3.771359039736635e-11, 3.8052491549353474e-11, 
    3.8338243799994838e-11, 3.8567172655793745e-11, 3.8735526247436129e-11, 
    3.8839692177587588e-11, 3.8876525747128163e-11, 3.8843766184788602e-11, 
    3.8740482958004772e-11, 3.8567493650226875e-11, 3.8327705827854285e-11, 
    3.8026321444551017e-11, 3.7670868890822333e-11, 3.7271053618495285e-11, 
    3.6838414620165308e-11, 3.6385833570000914e-11, 3.5926910769685607e-11, 
    3.5475279098945308e-11, 3.5043909464785759e-11, 3.4644463098888771e-11, 
    3.4286726072019187e-11, 3.3978197320726366e-11, 3.3723801147760053e-11, 
    3.3525779282683345e-11, 3.3383726360826353e-11, 3.3294767519628807e-11, 
    3.3253830897324206e-11, 3.3254028463440172e-11, 3.3287065966916086e-11, 
    3.3343706204524024e-11, 3.3414221675958449e-11, 3.3488848739806894e-11, 
    3.3558199050855574e-11, 3.3613637660329068e-11, 3.3647602538324018e-11, 
    3.3653857671708545e-11, 3.3627674126005624e-11, 3.3565936583949885e-11, 
    3.3467164219944533e-11, 3.3331469046034434e-11, 3.3160442724235861e-11, 
    3.2957006921399663e-11, 3.2725208974640142e-11, 3.2470019322807115e-11, 
    3.2197135748167554e-11, 3.191279557766732e-11, 3.162360533426429e-11, 
    3.1336417942287342e-11, 3.1058211050838038e-11, 3.0795998365264175e-11, 
    3.0556725501926286e-11, 3.0347163639736608e-11, 3.0173760977093363e-11, 
    3.0042475530930776e-11, 2.9958543201592864e-11, 2.9926238498136624e-11, 
    2.9948574247228247e-11, 3.0027026365435574e-11, 3.0161249824306599e-11, 
    3.0348853583073443e-11, 3.0585244636126392e-11, 3.0863586170387082e-11, 
    3.1174856284846849e-11, 3.1508085284310968e-11, 3.185071603184788e-11, 
    3.2189131905764519e-11, 3.2509286059683331e-11, 3.2797451385322425e-11, 
    3.3040988282794432e-11, 3.3229126488465646e-11, 3.3353665326771525e-11, 
    3.3409564243984746e-11, 3.3395317940028683e-11, 3.3313141345215411e-11, 
    3.316888951265666e-11, 3.2971737480143066e-11, 3.27336173500802e-11, 
    3.2468481678466768e-11, 3.2191418952449728e-11, 3.1917722198469814e-11, 
    3.1661966176669178e-11, 3.1437177025687534e-11, 3.1254138464532159e-11, 
    3.1120915876069413e-11, 3.1042582730492299e-11, 3.102118857339879e-11, 
    3.1055938464057889e-11, 3.1143570052344262e-11, 3.1278839068553934e-11, 
    3.1455138864517495e-11, 3.1665133880483156e-11, 3.1901406971714235e-11, 
    3.2157035566676606e-11, 3.2426107098733008e-11, 3.2704100905499045e-11, 
    3.2988152673982162e-11, 3.3277162458032676e-11, 3.3571771381746342e-11, 
    3.3874163105605917e-11, 3.4187769784066226e-11, 3.4516822136950654e-11, 
    3.4865841461798122e-11, 3.5239069861224799e-11, 3.5639896083595962e-11, 
    3.6070320437413459e-11, 3.653051854127252e-11, 3.7018534362630473e-11, 
    3.7530156227416531e-11, 3.8058986024571625e-11, 3.8596732413661982e-11, 
    3.9133664674061074e-11, 3.9659259124266394e-11, 4.0162935218030128e-11, 
    4.0634840219054812e-11, 4.1066585640426255e-11, 4.1451892845622297e-11, 
    4.1787042994686345e-11, 4.2071112653124814e-11, 4.2305949291897784e-11, 
    4.2495888583965841e-11, 4.2647230985075827e-11, 4.2767545379413035e-11, 
    4.2864843561261961e-11, 4.2946734617074016e-11, 4.3019604331896574e-11, 
    4.3087941858449039e-11, 4.315383614600309e-11, 4.3216710660414243e-11, 
    4.327330219517584e-11, 4.3317881229557125e-11, 4.3342691878487665e-11, 
    4.3338560631329955e-11, 4.3295611331718239e-11, 4.3204045312485977e-11, 
    4.3054898149854521e-11, 4.2840746160792074e-11, 4.2556286646490712e-11, 
    4.2198780113171789e-11, 4.1768320269883916e-11, 4.1267928878005015e-11, 
    4.0703455606306067e-11, 4.0083325791609577e-11, 3.9418122421916286e-11, 
    3.8720059700352788e-11, 3.8002345873662089e-11, 3.7278504020782353e-11, 
    3.6561690064600771e-11, 3.5864032675026853e-11, 3.5196058726829792e-11, 
    3.4566249373983958e-11, 3.3980737312776364e-11, 3.3443204385373176e-11, 
    3.2954962005573984e-11, 3.2515224880630837e-11, 3.2121549991792828e-11, 
    3.1770402445576311e-11, 3.1457796080405117e-11, 3.1179948465715634e-11, 
    3.0933877772684201e-11, 3.0717890449384992e-11, 3.0531911261026576e-11, 
    3.0377614517714492e-11, 3.0258343826394792e-11, 3.017883435945187e-11, 
    3.0144774394702233e-11, 3.0162233733440698e-11, 3.0237013458937367e-11, 
    3.037399455233793e-11, 3.0576526029193398e-11, 3.0845897589191353e-11, 
    3.1180940384926038e-11, 3.1577766709971161e-11, 3.2029668714819843e-11, 
    3.2527170545762056e-11, 3.3058216297497205e-11, 3.360848897716168e-11, 
    3.4161856666469275e-11, 3.4700911333160604e-11, 3.5207590556883862e-11, 
    3.5663876324209342e-11, 3.605255731107107e-11, 3.6358008789417896e-11, 
    3.6566977391396336e-11, 3.6669327899328249e-11, 3.6658715709713793e-11, 
    3.6533118476130898e-11, 3.6295185244573338e-11, 3.5952366051637685e-11, 
    3.5516766470453472e-11, 3.5004721852830126e-11, 3.4436093428043284e-11, 
    3.3833295342307872e-11, 3.3220109476643623e-11, 3.2620357076907931e-11, 
    3.2056519344382499e-11, 3.1548397081615464e-11, 3.1111919074544437e-11, 
    3.0758191595503306e-11, 3.0492875727249299e-11, 3.0315932063098296e-11, 
    3.0221779868270822e-11, 3.0199839151334122e-11, 3.0235429183704692e-11, 
    3.0310932410194554e-11, 3.0407156571462322e-11, 3.0504746846761804e-11, 
    3.0585565779043477e-11, 3.0633920892844132e-11, 3.0637545571037216e-11, 
    3.0588291271893243e-11, 3.0482471784807432e-11, 3.0320868478013054e-11, 
    3.0108427083481384e-11, 2.9853669621475868e-11, 2.9567918732590798e-11, 
    2.9264377118535988e-11, 2.8957165837520206e-11, 2.8660358174683573e-11, 
    2.8387115120014214e-11, 2.8148920503595093e-11, 2.7954987166244447e-11, 
    2.7811835304936412e-11, 2.7723058143278326e-11, 2.7689272934213086e-11, 
    2.7708249521852556e-11, 2.7775197886996934e-11, 2.78832040767608e-11, 
    2.8023779089718356e-11, 2.8187494073070708e-11, 2.8364654363176622e-11, 
    2.854600269862689e-11, 2.872334472402689e-11, 2.8890109598144335e-11, 
    2.9041760202012655e-11, 2.9176030605257675e-11, 2.9292966963478713e-11, 
    2.9394772288807826e-11, 2.9485452813030697e-11, 2.957031727994584e-11, 
    2.9655361255116694e-11, 2.9746618665614118e-11, 2.9849516070087631e-11, 
    2.9968299999150714e-11, 3.0105582174342029e-11, 3.0262038989272413e-11, 
    3.0436255911961517e-11, 3.0624731074684106e-11, 3.0822004920919469e-11, 
    3.1020904724109945e-11, 3.1212852459786573e-11, 3.1388239169977091e-11, 
    3.1536825460749893e-11, 3.1648171380715066e-11, 3.171208703483482e-11, 
    3.171911878045675e-11, 3.1661030754847879e-11, 3.1531330284932054e-11, 
    3.1325755358043689e-11, 3.1042734164607053e-11, 3.0683755333034321e-11, 
    3.0253604425717703e-11, 2.9760421125514163e-11, 2.9215542725042149e-11, 
    2.863310291127853e-11, 2.8029415301301666e-11, 2.7422137246073508e-11, 
    2.6829301446507225e-11, 2.6268269374596081e-11, 2.575470836041204e-11, 
    2.5301670889418112e-11, 2.4918873653456158e-11, 2.4612215608893354e-11, 
    2.4383603245821615e-11, 2.4231046212234889e-11, 2.4149051331916784e-11, 
    2.4129207411578253e-11, 2.416093825929333e-11, 2.4232310406787107e-11, 
    2.4330846986118762e-11, 2.4444263227303804e-11, 2.4561080561533934e-11, 
    2.4671101987245576e-11, 2.4765740733419033e-11, 2.4838214824457991e-11, 
    2.4883651641189265e-11, 2.4899122296090412e-11,
  // Sqw-Na(7, 0-1999)
    0.023501517064793455, 0.023502513929617781, 0.023505371511282978, 
    0.023509696919003415, 0.023514855531213255, 0.023520000261875919, 
    0.023524110503033782, 0.023526038781915695, 0.023524562724274799, 
    0.023518439575631225, 0.023506460335024612, 0.0234875005337974, 
    0.023460564865840722, 0.023424823249868675, 0.023379636462525027, 
    0.023324570186747169, 0.023259397118545896, 0.023184087601336098, 
    0.023098790040424613, 0.023003803025631795, 0.0228995416030662, 
    0.022786500449944472, 0.022665216800297101, 0.022536235844704537, 
    0.022400081001278938, 0.022257230959112299, 0.022108104770621837, 
    0.021953055563437688, 0.021792372707188545, 0.021626291558628122, 
    0.02145500927231456, 0.021278704653135853, 0.021097559685539086, 
    0.020911780237528734, 0.020721613527233552, 0.020527360260324728, 
    0.020329379880774857, 0.020128088085344543, 0.019923946571676687, 
    0.019717445841106213, 0.019509082670105274, 0.019299334508364751, 
    0.0190886334777088, 0.018877342777480322, 0.018665738122933932, 
    0.018453996364238244, 0.018242192702566114, 0.018030307016657886, 
    0.017818238841717526, 0.017605829616747587, 0.017392890046592207, 
    0.017179229902566859, 0.016964687371062444, 0.016749155173765296, 
    0.016532601104309066, 0.016315081292647131, 0.016096745327523785, 
    0.015877833228910659, 0.015658665054670114, 0.015439624552856298, 
    0.015221138666390317, 0.01500365483268885, 0.0147876179112924, 
    0.014573448269170116, 0.014361522134328635, 0.014152154883080102, 
    0.013945587538520729, 0.013741976489884114, 0.013541386324660344, 
    0.013343785691352372, 0.0131490462406145, 0.012956944862807516, 
    0.01276716957808023, 0.012579329475348608, 0.012392968994871583, 
    0.012207586592780375, 0.012022657436848124, 0.011837659313901424, 
    0.011652100454514196, 0.011465547581059702, 0.01127765223395117, 
    0.011088173379940286, 0.01089699447747472, 0.0107041335557854, 
    0.010509745414286087, 0.010314115701715428, 0.010117647312720541, 
    0.0099208401654913552, 0.0097242659302720445, 0.009528539616366934, 
    0.0093342900689741722, 0.0091421313751783757, 0.0089526369507855336, 
    0.0087663177136942331, 0.008583605293889341, 0.0084048407388634516, 
    0.0082302686994580685, 0.00806003667169225, 0.0078941985612759284, 
    0.0077327216511624153, 0.0075754959944441423, 0.0074223453144051819, 
    0.0072730386450590165, 0.0071273021524214967, 0.0069848307969482002, 
    0.0068452996899852807, 0.0067083751285693495, 0.0065737253438086897, 
    0.0064410309656235997, 0.0063099951053745195, 0.0061803528168442468, 
    0.0060518795529317564, 0.0059243981293495675, 0.0057977836702571917, 
    0.005671966063770616, 0.0055469296002820167, 0.0054227096883082719, 
    0.0052993868108084999, 0.0051770781595298961, 0.0050559276234622636, 
    0.0049360949724765249, 0.0048177451428200709, 0.0047010384872401261, 
    0.0045861227061617747, 0.0044731269501070868, 0.0043621583112775364, 
    0.0042533006432222279, 0.0041466154000309747, 0.0040421440017937398, 
    0.0039399111310437661, 0.0038399283517667731, 0.0037421975109799967, 
    0.0036467135142484179, 0.0035534662348396906, 0.0034624414929225081, 
    0.0033736211997734151, 0.0032869828818050538, 0.0032024988682317597, 
    0.0031201354414327645, 0.0030398522160852803, 0.0029616019438093648, 
    0.0028853308498758123, 0.0028109795136185677, 0.0027384842188454498, 
    0.0026677786353908051, 0.0025987956541426382, 0.0025314691870359268, 
    0.0024657357584292197, 0.0024015357499539971, 0.0023388142106699266, 
    0.0022775212008583636, 0.0022176116939312922, 0.0021590451103863598, 
    0.0021017845953737657, 0.002045796173609895, 0.0019910479201571164, 
    0.0019375092729431874, 0.0018851505847147228, 0.001833942972125183, 
    0.0017838584730652377, 0.001734870476275092, 0.0016869543460105124, 
    0.0016400881346080583, 0.0015942532612140308, 0.0015494350375383303, 
    0.0015056229406465011, 0.0014628105655193433, 0.0014209952315175011, 
    0.0013801772609988224, 0.0013403589889898126, 0.001301543594597567, 
    0.0012637338638855158, 0.0012269309983582964, 0.0011911335733209942, 
    0.001156336728489036, 0.0011225316431441406, 0.0010897053145198727, 
    0.0010578406257380996, 0.0010269166626832365, 0.00099690922072013318, 
    0.00096779143363232337, 0.00093953445846051088, 0.00091210815945001289, 
    0.00088548174936071999, 0.00085962436364992627, 0.00083450555922042651, 
    0.00081009574181165327, 0.00078636653299759825, 0.00076329108868096191, 
    0.00074084437673220592, 0.00071900341381323537, 0.0006977474528453249, 
    0.00067705810549600833, 0.00065691938051208848, 0.00063731761992276642, 
    0.00061824132125233426, 0.00059968084405160693, 0.00058162801160503252, 
    0.0005640756314562531, 0.00054701696925525233, 0.0005304452175647975, 
    0.00051435300354419201, 0.0004987319765330534, 0.00048357250896608497, 
    0.00046886353288172342, 0.00045459252107111548, 0.00044074560830770497, 
    0.00042730783565376052, 0.00041426349080787866, 0.00040159651068799861, 
    0.00038929090934276958, 0.00037733119484617051, 0.00036570274268949408, 
    0.0003543920997009075, 0.00034338720085350826, 0.00033267749051883256, 
    0.00032225394880308725, 0.00031210903165618774, 0.00030223653970624367, 
    0.00029263143472522523, 0.00028328962405337678, 0.00027420773231615113, 
    0.00026538287678411546, 0.00025681245843491517, 0.00024849397599290658, 
    0.00024042486577177891, 0.00023260236671300379, 0.00022502340803837845, 
    0.00021768451653516381, 0.00021058174146436985, 0.00020371059694796118, 
    0.00019706602381106716, 0.00019064237455783446, 0.00018443342588417982, 
    0.00017843242253242633, 0.00017263215431917084, 0.00016702506505834102, 
    0.00016160338835117261, 0.00015635930147060961, 0.00015128508551838233, 
    0.00014637327827479022, 0.00014161680610079718, 0.00013700908302545525, 
    0.00013254406860884873, 0.000128216280887105, 0.00012402076605775447, 
    0.0001199530318116072, 0.00011600895562623104, 0.00011218468227378174, 
    0.00010847652583291696, 0.00010488089045786401, 0.00010139422116613048, 
    9.8012991346671781e-05, 9.4733728176268526e-05, 9.1553071411399373e-05, 
    8.8467855885886963e-05, 8.5475204203647282e-05, 8.2572614114988512e-05, 
    7.9758025192985574e-05, 7.7029851682798949e-05, 7.4386972481898302e-05, 
    7.1828674575117408e-05, 6.935455217023018e-05, 6.6964369467647291e-05, 
    6.4657899703023252e-05, 6.2434756229669603e-05, 6.029423258928939e-05, 
    5.8235167661996442e-05, 5.6255849265790386e-05, 5.4353965404921559e-05, 
    5.2526607316295281e-05, 5.077032318075448e-05, 4.9081216474919607e-05, 
    4.7455078966582668e-05, 4.5887545667679223e-05, 4.4374257836296597e-05, 
    4.2911020354021253e-05, 4.1493941330683985e-05, 4.0119544313687534e-05, 
    3.878484664661878e-05, 3.7487400950858949e-05, 3.6225300041525858e-05, 
    3.4997148535476166e-05, 3.3802006746004138e-05, 3.2639314050102198e-05, 
    3.1508799713468899e-05, 3.0410389191731067e-05, 2.9344113287247786e-05, 
    2.831002636558152e-05, 2.7308138293260365e-05, 2.6338363025496705e-05, 
    2.5400485023804273e-05, 2.4494143070616467e-05, 2.3618829695207032e-05, 
    2.2773903414476989e-05, 2.195861036806879e-05, 2.1172111690157506e-05, 
    2.041351307892966e-05, 1.9681893437207666e-05, 1.8976330087077218e-05, 
    1.8295918819174648e-05, 1.7639787839311975e-05, 1.7007105441223506e-05, 
    1.6397081901704293e-05, 1.5808966613567208e-05, 1.5242041815406642e-05, 
    1.4695614432941415e-05, 1.4169007524150024e-05, 1.3661552641092099e-05, 
    1.3172584123377814e-05, 1.270143596497719e-05, 1.224744149868382e-05, 
    1.180993576681304e-05, 1.1388260136054191e-05, 1.0981768496349613e-05, 
    1.0589834275128156e-05, 1.0211857496170451e-05, 9.8472712023738457e-06, 
    9.4955467145124353e-06, 9.1561973819699097e-06, 8.8287806612259512e-06, 
    8.5128985087507892e-06, 8.208196178535617e-06, 7.914359569686074e-06, 
    7.6311112829518073e-06, 7.3582055361665393e-06, 7.0954220762781977e-06, 
    6.8425592303907965e-06, 6.5994262695198006e-06, 6.3658353197114458e-06, 
    6.1415931347374638e-06, 5.9264931274534312e-06, 5.7203081203685982e-06, 
    5.5227843022980962e-06, 5.3336368521046114e-06, 5.1525476098985144e-06, 
    4.9791650449650555e-06, 4.8131066040358722e-06, 4.6539633417821025e-06, 
    4.5013065604111334e-06, 4.3546960344847949e-06, 4.2136892861348683e-06, 
    4.0778513108164637e-06, 3.9467641379745214e-06, 3.8200356397510532e-06, 
    3.6973070700746937e-06, 3.5782589169489964e-06, 3.4626147766981541e-06, 
    3.3501431005287624e-06, 3.2406568142868045e-06, 3.1340109602818785e-06, 
    3.030098646477015e-06, 2.9288456996707862e-06, 2.830204496288401e-06, 
    2.7341474763163991e-06, 2.6406608299131571e-06, 2.5497387815928476e-06, 
    2.4613787927426785e-06, 2.3755778710130376e-06, 2.2923300338329036e-06, 
    2.2116248399609929e-06, 2.1334467964480729e-06, 2.0577753800021363e-06, 
    1.9845853895194445e-06, 1.9138473682771103e-06, 1.8455278939986819e-06, 
    1.7795896182442402e-06, 1.7159910293542873e-06, 1.654685998174585e-06, 
    1.5956232313006585e-06, 1.5387457921218966e-06, 1.4839908537243401e-06, 
    1.4312898200696618e-06, 1.3805689009824094e-06, 1.3317501604492944e-06, 
    1.2847529890717905e-06, 1.2394958891899499e-06, 1.1958984153700733e-06, 
    1.1538830878360368e-06, 1.1133770960858785e-06, 1.0743136319156136e-06, 
    1.0366327334435306e-06, 1.0002815770810144e-06, 9.6521421706406311e-07, 
    9.3139083308777705e-07, 8.9877659962377995e-07, 8.6734032799355377e-07, 
    8.3705305089780965e-07, 8.0788671516744868e-07, 7.7981312373982017e-07, 
    7.5280322412862244e-07, 7.2682678515121607e-07, 7.0185244274195414e-07, 
    6.7784803971881098e-07, 6.5478114039833963e-07, 6.3261957754116126e-07, 
    6.1133188893208355e-07, 5.908875258818786e-07, 5.7125676113773052e-07, 
    5.5241028326219908e-07, 5.3431852759405119e-07, 5.1695085075356783e-07, 
    5.0027469552257825e-07, 4.8425490945088197e-07, 4.6885336943078795e-07, 
    4.5402902796579466e-07, 4.3973843956725102e-07, 4.2593675767155991e-07, 
    4.1257912356803618e-07, 3.9962231095431172e-07, 3.8702645061677613e-07, 
    3.7475664624474372e-07, 3.6278430456630052e-07, 3.5108803930011853e-07, 
    3.3965406136481409e-07, 3.2847602984106076e-07, 3.1755439894276297e-07, 
    3.0689534841173344e-07, 2.9650942075758453e-07, 2.8641000647243411e-07, 
    2.766118163270469e-07, 2.6712946194558368e-07, 2.5797623567323723e-07, 
    2.4916314531449594e-07, 2.4069822345266467e-07, 2.3258610080845497e-07, 
    2.2482781092336484e-07, 2.174207819109275e-07, 2.1035896869863415e-07, 
    2.0363308535221033e-07, 1.9723090761032388e-07, 1.9113762853301089e-07, 
    1.8533626087347348e-07, 1.7980808715425962e-07, 1.7453316000305601e-07, 
    1.6949085210126132e-07, 1.6466044686326376e-07, 1.6002175095954131e-07, 
    1.5555569903909117e-07, 1.512449132412785e-07, 1.4707417620406155e-07, 
    1.43030778574598e-07, 1.3910470982113034e-07, 1.3528867452153113e-07, 
    1.3157793266159648e-07, 1.2796998049090756e-07, 1.244641044764851e-07, 
    1.2106085381734873e-07, 1.1776148386320337e-07, 1.1456742390609512e-07, 
    1.114798172025158e-07, 1.0849917053985934e-07, 1.0562513590612985e-07, 
    1.0285643065832343e-07, 1.0019088606436381e-07, 9.7625600169470258e-08, 
    9.5157159987687629e-08, 9.2781892207288783e-08, 9.0496100466595892e-08, 
    8.8296251704544267e-08, 8.6179082842967043e-08, 8.414161181175767e-08, 
    8.218105159248823e-08, 8.0294641361689501e-08, 7.8479422280404228e-08, 
    7.6731995813669269e-08, 7.5048307082150351e-08, 7.342349470207832e-08, 
    7.1851840513497329e-08, 7.0326839581889748e-08, 6.8841393525855296e-08, 
    6.7388112307464215e-08, 6.5959692817803016e-08, 6.4549330934758916e-08, 
    6.3151117911179237e-08, 6.1760374272601102e-08, 6.0373883226923085e-08, 
    5.8990000497848062e-08, 5.7608634673807304e-08, 5.6231109832119887e-08, 
    5.4859936155969678e-08, 5.3498523515414498e-08, 5.2150875302973982e-08, 
    5.0821296372922359e-08, 4.9514140112137627e-08, 4.8233608530718989e-08, 
    4.6983607358630815e-08, 4.576764868151816e-08, 4.4588787323462538e-08, 
    4.3449575656162135e-08, 4.2352023542742434e-08, 4.129755560359279e-08, 
    4.0286964322314106e-08, 3.9320364046159088e-08, 3.8397155187398558e-08, 
    3.7516010034185852e-08, 3.6674890327475584e-08, 3.5871103548126826e-08, 
    3.5101399568057289e-08, 3.4362103996323884e-08, 3.364927943978372e-08, 
    3.2958902580944673e-08, 3.2287043123856109e-08, 3.1630031181945476e-08, 
    3.0984601289239071e-08, 3.0348004521918775e-08, 2.9718083416478975e-08, 
    2.9093308126346439e-08, 2.8472775036945248e-08, 2.7856171799377288e-08, 
    2.7243714185627936e-08, 2.6636061554767098e-08, 2.6034218046234523e-08, 
    2.5439426941326952e-08, 2.4853065091646773e-08, 2.4276543809627777e-08, 
    2.3711221226312398e-08, 2.3158329946956862e-08, 2.2618921751190554e-08, 
    2.2093829646725538e-08, 2.1583645650541509e-08, 2.1088711755246834e-08, 
    2.0609120749575693e-08, 2.0144723932386449e-08, 1.9695143362936923e-08, 
    1.925978786184495e-08, 1.8837873137501524e-08, 1.8428447928250498e-08, 
    1.8030428393583061e-08, 1.7642643057480844e-08, 1.7263889265765636e-08, 
    1.6893000413539389e-08, 1.6528920665596438e-08, 1.6170781761870246e-08, 
    1.581797438282218e-08, 1.5470205927570681e-08, 1.5127536626454145e-08, 
    1.4790387808319836e-08, 1.4459518687906263e-08, 1.4135971861783165e-08, 
    1.3820991194973644e-08, 1.3515919457308046e-08, 1.3222085294864826e-08, 
    1.2940690660685941e-08, 1.2672709339014093e-08, 1.2418805977899643e-08, 
    1.2179282162992388e-08, 1.1954053181828047e-08, 1.1742655544449727e-08, 
    1.1544282564828115e-08, 1.1357842780026296e-08, 1.1182034796740238e-08, 
    1.1015431358055686e-08, 1.0856565872270894e-08, 1.0704015278610912e-08, 
    1.0556474449763891e-08, 1.0412818333927434e-08, 1.0272149460262648e-08, 
    1.0133829152547765e-08, 9.9974918791786891e-09, 9.863042549123248e-09, 
    9.7306374997932345e-09, 9.6006502228935209e-09, 9.4736238314812353e-09, 
    9.3502127289262357e-09, 9.231116947816326e-09, 9.1170130297962788e-09, 
    9.0084860024673654e-09, 8.9059670569136904e-09, 8.8096815901923348e-09, 
    8.7196115465699524e-09, 8.6354753654996055e-09, 8.5567273765920816e-09, 
    8.4825773519254091e-09, 8.4120290937298242e-09, 8.3439357293703988e-09, 
    8.2770677437204546e-09, 8.2101889890950144e-09, 8.1421349476997267e-09, 
    8.0718875647226494e-09, 7.9986409086509484e-09, 7.9218528996466987e-09, 
    7.8412791729255433e-09, 7.7569868155801275e-09, 7.669347035887099e-09, 
    7.5790077033320195e-09, 7.4868479517889996e-09, 7.3939185344708292e-09, 
    7.3013723105839644e-09, 7.210389986169148e-09, 7.1221060910227882e-09, 
    7.0375401201134323e-09, 6.9575369026524653e-09, 6.88271962698882e-09, 
    6.8134577033998015e-09, 6.749850794297524e-09, 6.6917290794708257e-09, 
    6.6386690832509437e-09, 6.5900233282239697e-09, 6.5449617028815335e-09, 
    6.5025216449532273e-09, 6.46166423728329e-09, 6.4213328710964171e-09, 
    6.3805114087437333e-09, 6.3382786553405574e-09, 6.2938564708026566e-09, 
    6.2466489613520243e-09, 6.1962709351830686e-09, 6.142564074822389e-09, 
    6.085600216847907e-09, 6.0256715258905737e-09, 5.9632683048366248e-09, 
    5.8990456524623646e-09, 5.8337810811629245e-09, 5.7683254997580169e-09, 
    5.7035506768697909e-09, 5.640296261955806e-09, 5.5793198029969548e-09, 
    5.5212527489032972e-09, 5.4665652761252537e-09, 5.4155420053882875e-09, 
    5.3682700847217563e-09, 5.3246400818084454e-09, 5.2843594211129935e-09, 
    5.2469770159273444e-09, 5.2119172094915136e-09, 5.1785202896488551e-09, 
    5.1460867557806232e-09, 5.1139220795484345e-09, 5.0813791048049493e-09, 
    5.0478952694611317e-09, 5.0130226463260555e-09, 4.9764490996426772e-09, 
    4.9380098628683776e-09, 4.8976892311322572e-09, 4.8556129826238301e-09, 
    4.8120324043167743e-09, 4.7673015273100255e-09, 4.7218491777235496e-09, 
    4.6761479304602825e-09, 4.63068182367611e-09, 4.5859149097671641e-09, 
    4.5422623218215237e-09, 4.5000655690596831e-09, 4.4595732276966129e-09, 
    4.4209281091345768e-09, 4.3841613721825545e-09, 4.349193870003092e-09, 
    4.3158443546965979e-09, 4.2838440273604285e-09, 4.2528562867050641e-09, 
    4.2225004236493282e-09, 4.1923775626692951e-09, 4.1620972285645283e-09, 
    4.1313026742692397e-09, 4.099693404746006e-09, 4.0670433462910825e-09, 
    4.0332136995612129e-09, 3.9981596221147986e-09, 3.9619306413354787e-09, 
    3.9246648827792158e-09, 3.8865778859225645e-09, 3.8479468887515683e-09, 
    3.8090919570172394e-09, 3.7703552585723017e-09, 3.7320800283547751e-09, 
    3.6945904723484803e-09, 3.6581739217429987e-09, 3.6230660805661397e-09, 
    3.589440172348686e-09, 3.5574002733700164e-09, 3.5269790888007445e-09, 
    3.498139947579761e-09, 3.4707827778495553e-09, 3.4447534483223106e-09, 
    3.419855905868251e-09, 3.3958662212025646e-09, 3.3725477786519098e-09, 
    3.3496665769903188e-09, 3.3270058428989671e-09, 3.3043789495001813e-09, 
    3.2816399658452926e-09, 3.258691056077262e-09, 3.2354864021194609e-09, 
    3.2120322912866106e-09, 3.1883835039632477e-09, 3.1646361896712968e-09, 
    3.1409178803415925e-09, 3.1173752831743171e-09, 3.0941609027380488e-09, 
    3.0714193960671151e-09, 3.0492748053311216e-09, 3.0278195402751521e-09, 
    3.0071060310145414e-09, 2.9871415834255482e-09, 2.9678868740374898e-09, 
    2.9492580544850841e-09, 2.9311323393211913e-09, 2.9133564711393682e-09, 
    2.8957574404038462e-09, 2.8781544701163416e-09, 2.8603714144459709e-09, 
    2.8422484981085929e-09, 2.8236526490757703e-09, 2.8044855914576661e-09, 
    2.7846893257739131e-09, 2.7642486134211173e-09, 2.7431905721646326e-09, 
    2.7215814850048761e-09, 2.6995213161209232e-09, 2.6771363854467276e-09, 
    2.6545708976021487e-09, 2.6319778713151883e-09, 2.6095101773078303e-09, 
    2.5873121197984895e-09, 2.5655121232700233e-09, 2.544216779436524e-09, 
    2.5235065578293979e-09, 2.5034332547403741e-09, 2.4840192667726015e-09, 
    2.4652585642705114e-09, 2.4471192899253259e-09, 2.4295476757125448e-09, 
    2.4124731075556346e-09, 2.3958139096785933e-09, 2.3794835984472348e-09, 
    2.3633971254907549e-09, 2.3474768580837157e-09, 2.3316578510192721e-09, 
    2.3158921751261755e-09, 2.3001519935359371e-09, 2.2844312498844302e-09, 
    2.2687457945408494e-09, 2.2531320170467393e-09, 2.2376439694875102e-09, 
    2.2223492501574233e-09, 2.2073238228026859e-09, 2.1926462157951994e-09, 
    2.1783914223101786e-09, 2.1646250245830524e-09, 2.1513979100086319e-09, 
    2.1387420590479053e-09, 2.1266676581855983e-09, 2.1151618305927833e-09, 
    2.1041890057350165e-09, 2.0936929430305556e-09, 2.0836001586609927e-09, 
    2.0738245153608506e-09, 2.0642725075792379e-09, 2.0548488933296365e-09, 
    2.045462142546864e-09, 2.0360293935295594e-09, 2.0264805164527568e-09, 
    2.0167611354217456e-09, 2.0068344331764425e-09, 1.996681808514725e-09, 
    1.986302399739173e-09, 1.975711708254483e-09, 1.9649394587802843e-09, 
    1.9540269628441355e-09, 1.9430241274472927e-09, 1.9319863544288364e-09, 
    1.920971387203503e-09, 1.910036298914286e-09, 1.8992346231038875e-09, 
    1.8886137714489406e-09, 1.8782127295174748e-09, 1.8680601693466022e-09, 
    1.8581730134557087e-09, 1.8485555689937931e-09, 1.8391992677529726e-09, 
    1.8300831467909869e-09, 1.8211750280422478e-09, 1.8124334474098363e-09, 
    1.8038102087307597e-09, 1.7952534792701525e-09, 1.7867112047728815e-09, 
    1.7781346512278278e-09, 1.7694817681764987e-09, 1.7607201828711717e-09, 
    1.7518295134738811e-09, 1.7428028794225293e-09, 1.7336474068761877e-09, 
    1.7243837407243547e-09, 1.715044537829596e-09, 1.7056720897089929e-09, 
    1.6963152296088613e-09, 1.6870258077381526e-09, 1.6778549421022932e-09, 
    1.6688494220876597e-09, 1.6600484707030883e-09, 1.6514811583059165e-09, 
    1.6431646030806435e-09, 1.6351031264244946e-09, 1.627288337710108e-09, 
    1.619700163262365e-09, 1.6123086282955086e-09, 1.6050762972063003e-09, 
    1.5979610747503909e-09, 1.5909191963060325e-09, 1.5839081154793825e-09, 
    1.5768891325637594e-09, 1.5698295292426511e-09, 1.5627041414184634e-09, 
    1.5554962599581334e-09, 1.5481978817374186e-09, 1.5408093310816779e-09, 
    1.5333383634946682e-09, 1.5257988442803927e-09, 1.5182091744961079e-09, 
    1.5105905709954851e-09, 1.5029653719431468e-09, 1.4953554433760496e-09, 
    1.4877808209331734e-09, 1.4802586055119426e-09, 1.472802194957386e-09, 
    1.465420805603223e-09, 1.4581193358461786e-09, 1.4508984858515305e-09, 
    1.4437551513749821e-09, 1.4366830029203715e-09, 1.4296732426735659e-09, 
    1.422715467355287e-09, 1.4157986082587608e-09, 1.4089118692125285e-09, 
    1.4020456491513402e-09, 1.3951923606835858e-09, 1.3883471214154103e-09, 
    1.3815082506297156e-09, 1.3746775566838149e-09, 1.3678603645329614e-09, 
    1.3610653013199686e-09, 1.3543038140912297e-09, 1.3475894823381954e-09, 
    1.3409371277230238e-09, 1.3343618060911809e-09, 1.3278777157443811e-09, 
    1.3214971175941502e-09, 1.3152293095798827e-09, 1.3090797503030282e-09, 
    1.3030493524419482e-09, 1.297134043185837e-09, 1.2913245876571619e-09, 
    1.2856067336018242e-09, 1.2799616538817304e-09, 1.2743667069456474e-09, 
    1.2687964602842438e-09, 1.2632239512938851e-09, 1.2576220860992334e-09, 
    1.2519651360457305e-09, 1.2462302026858794e-09, 1.2403985854917574e-09, 
    1.2344569249736114e-09, 1.2283980847764241e-09, 1.2222216464525783e-09, 
    1.2159340420277702e-09, 1.2095482433012568e-09, 1.2030830793382075e-09, 
    1.1965621718667241e-09, 1.1900126047050121e-09, 1.1834633803182515e-09, 
    1.1769438060306556e-09, 1.1704818783474914e-09, 1.1641028160168971e-09, 
    1.1578278086208534e-09, 1.1516730894142773e-09, 1.1456493375136711e-09, 
    1.139761492727308e-09, 1.1340089059068669e-09, 1.1283858509231118e-09, 
    1.1228822704124946e-09, 1.1174847306231959e-09, 1.1121774467678265e-09, 
    1.1069433413881789e-09, 1.1017649910139065e-09, 1.0966254791462798e-09, 
    1.0915090558418328e-09, 1.0864016333029184e-09, 1.0812910915483291e-09, 
    1.0761674561581874e-09, 1.0710229442901387e-09, 1.0658519600395463e-09, 
    1.0606510149012989e-09, 1.0554186538044725e-09, 1.0501553490723804e-09, 
    1.0448633995505914e-09, 1.0395467721854805e-09, 1.0342109384146516e-09, 
    1.0288626225542063e-09, 1.0235095116658652e-09, 1.0181598683010806e-09, 
    1.0128221181452015e-09, 1.0075043669209076e-09, 1.0022139320213357e-09, 
    9.9695687266418389e-10, 9.9173761029466328e-10, 9.8655859318341728e-10, 
    9.8142013418342962e-10, 9.7632036514120952e-10, 9.7125537683086915e-10, 
    9.6621951102964536e-10, 9.6120583271957636e-10, 9.562067328277629e-10, 
    9.5121465041221812e-10, 9.4622282996795529e-10, 9.4122610282859897e-10, 
    9.3622157245913337e-10, 9.3120918954300292e-10, 9.2619210585224962e-10, 
    9.2117680638014088e-10, 9.1617295811232939e-10, 9.111930075472273e-10, 
    9.0625152049650172e-10, 9.0136435586772408e-10, 8.965476968109053e-10, 
    8.9181707923057474e-10, 8.871864439182957e-10, 8.8266734970842834e-10, 
    8.7826835310732455e-10, 8.7399464687117582e-10, 8.6984791771150815e-10, 
    8.6582646331649903e-10, 8.6192548754634853e-10, 8.5813758795571267e-10, 
    8.5445328933892496e-10, 8.5086168231963068e-10, 8.4735100976450295e-10, 
    8.4390925455086391e-10, 8.4052460992409312e-10, 8.3718590495796696e-10, 
    8.3388288392503138e-10, 8.3060642001575786e-10, 8.2734859336682999e-10, 
    8.2410269452170358e-10, 8.208630988860748e-10, 8.1762508764394916e-10, 
    8.1438456856776574e-10, 8.1113778007005092e-10, 8.0788094154326048e-10, 
    8.0460996535460057e-10, 8.013201995046723e-10, 7.9800631487385914e-10, 
    7.9466229396435138e-10, 7.9128162811041911e-10, 7.8785765546793856e-10, 
    7.8438408304867187e-10, 7.8085559772059378e-10, 7.7726856342994643e-10, 
    7.7362168147809617e-10, 7.6991659077743074e-10, 7.6615825330360265e-10, 
    7.6235517366029389e-10, 7.585192845449542e-10, 7.5466560266253628e-10, 
    7.5081157464527776e-10, 7.4697623447812112e-10, 7.431791687857051e-10, 
    7.3943945206417898e-10, 7.3577456365586087e-10, 7.321994565770046e-10, 
    7.2872578604743044e-10, 7.2536140962401461e-10, 7.2211014209255778e-10, 
    7.1897180892851836e-10, 7.1594251454216199e-10, 7.1301513829105659e-10, 
    7.1017992271943699e-10, 7.0742516203917573e-10, 7.0473784310212663e-10, 
    7.0210426823567347e-10, 6.995105665273029e-10, 6.9694315048937747e-10, 
    6.9438904768301616e-10, 6.9183621516692945e-10, 6.8927380394230528e-10, 
    6.8669242770040678e-10, 6.8408441273251834e-10, 6.8144407717262879e-10, 
    6.7876794285536683e-10, 6.7605493190530052e-10, 6.7330642891187652e-10, 
    6.7052624122393145e-10, 6.6772037473605883e-10, 6.6489668118144764e-10, 
    6.620643359611159e-10, 6.5923323697653902e-10, 6.564133251893696e-10, 
    6.5361394609061207e-10, 6.5084324425249537e-10, 6.4810771223467886e-10, 
    6.4541187127090987e-10, 6.427581526358988e-10, 6.4014692387767241e-10, 
    6.3757669454815315e-10, 6.350444365439559e-10, 6.325460008864748e-10, 
    6.300765636570437e-10, 6.2763110993428362e-10, 6.2520486677469339e-10, 
    6.2279371327689395e-10, 6.2039449600153894e-10, 6.1800528914692504e-10, 
    6.1562553294333518e-10, 6.1325610560389037e-10, 6.1089926490699374e-10, 
    6.0855853393189011e-10, 6.0623844909618533e-10, 6.0394428187699619e-10, 
    6.0168165720256149e-10, 5.9945615990359693e-10, 5.972729120090151e-10, 
    5.9513617548735134e-10, 5.9304897228058234e-10, 5.9101280324266037e-10, 
    5.8902742378861766e-10, 5.8709076572042301e-10, 5.8519894041442063e-10, 
    5.8334639867215028e-10, 5.8152618602631341e-10, 5.7973031385721315e-10, 
    5.7795020891743798e-10, 5.7617721931967537e-10, 5.7440314219943668e-10, 
    5.7262073860774607e-10, 5.7082419287333392e-10, 5.6900950382848928e-10, 
    5.6717473012049591e-10, 5.6532013154850943e-10, 5.6344812768345381e-10, 
    5.615631271132061e-10, 5.5967118661031024e-10, 5.5777957392615194e-10, 
    5.5589621292180095e-10, 5.5402910741162734e-10, 5.5218574261776171e-10, 
    5.503725485689482e-10, 5.485944369176625e-10, 5.468544746736665e-10, 
    5.4515368168300275e-10, 5.4349099670694731e-10, 5.4186336403876859e-10, 
    5.4026595303646163e-10, 5.3869245224352598e-10, 5.3713542375209936e-10, 
    5.35586664295155e-10, 5.340375579707802e-10, 5.3247937479436819e-10, 
    5.3090354577991403e-10, 5.2930185630783078e-10, 5.2766663658709397e-10, 
    5.2599089496654697e-10, 5.2426847555545273e-10, 5.2249419473406577e-10, 
    5.206640120207823e-10, 5.1877518950157738e-10, 5.1682646807908122e-10, 
    5.1481818143993993e-10, 5.1275234870478802e-10, 5.1063266015711963e-10, 
    5.0846438073797672e-10, 5.062541291930034e-10, 5.0400957325078346e-10, 
    5.0173902668276626e-10, 4.9945102241593542e-10, 4.9715386480102867e-10, 
    4.9485525730077541e-10, 4.9256198707158674e-10, 4.9027976929262036e-10, 
    4.8801320170923167e-10, 4.8576588263735425e-10, 4.8354062183387786e-10, 
    4.8133974658464491e-10, 4.7916541720778906e-10, 4.7701993644818076e-10, 
    4.7490595869245178e-10, 4.7282660662224396e-10, 4.7078543854299832e-10, 
    4.6878628794843906e-10, 4.6683297906929253e-10, 4.6492896340909367e-10, 
    4.6307691167149411e-10, 4.6127832455911311e-10, 4.595331878158996e-10, 
    4.5783973868898084e-10, 4.5619434297397026e-10, 4.5459151593297697e-10, 
    4.530240651314598e-10, 4.5148336951682421e-10, 4.4995972370985403e-10, 
    4.4844278370189239e-10, 4.4692202537512239e-10, 4.4538723305142442e-10, 
    4.4382896330870893e-10, 4.4223898317818562e-10, 4.4061064690487517e-10, 
    4.3893920843463264e-10, 4.3722203682882792e-10, 4.3545874357775673e-10, 
    4.3365116903132703e-10, 4.3180327601946925e-10, 4.2992089429914094e-10, 
    4.2801138567450951e-10, 4.2608319710735274e-10, 4.2414538020926173e-10, 
    4.2220709127935775e-10, 4.2027714043853523e-10, 4.1836359760740805e-10, 
    4.1647352768297365e-10, 4.1461284751904438e-10, 4.1278631333511502e-10, 
    4.1099762263128766e-10, 4.0924960566555496e-10, 4.0754443636144704e-10, 
    4.0588386306874312e-10, 4.0426936716688865e-10, 4.0270226910177191e-10, 
    4.0118371537607266e-10, 3.9971459585419365e-10, 3.98295385403755e-10, 
    3.9692595015441998e-10, 3.956053502067188e-10, 3.9433169408201168e-10, 
    3.9310205870439982e-10, 3.9191251051027677e-10, 3.9075821997548044e-10, 
    3.8963368045010855e-10, 3.8853298292832637e-10, 3.8745013986555538e-10, 
    3.8637940437509855e-10, 3.8531555832196723e-10, 3.8425413000104637e-10, 
    3.831915262804375e-10, 3.8212505967490822e-10, 3.8105288217920169e-10, 
    3.7997382177700237e-10, 3.7888716667712814e-10, 3.777923893817834e-10, 
    3.7668889091576673e-10, 3.7557573895793865e-10, 3.7445148265812842e-10, 
    3.7331402915069969e-10, 3.7216061529433122e-10, 3.7098786558245409e-10, 
    3.6979195734650139e-10, 3.6856883768715364e-10, 3.6731452598766414e-10, 
    3.660254319104705e-10, 3.6469869146378382e-10, 3.6333247172646218e-10, 
    3.6192623721603489e-10, 3.6048093645706299e-10, 3.5899911912941175e-10, 
    3.5748493098498215e-10, 3.5594403749666632e-10, 3.5438342265676522e-10, 
    3.528111213792295e-10, 3.512358591054133e-10, 3.4966665813698536e-10, 
    3.4811239531972156e-10, 3.465813751167192e-10, 3.4508091175310222e-10, 
    3.4361698205353469e-10, 3.4219393022102929e-10, 3.408142860571422e-10, 
    3.3947867260259731e-10, 3.3818584225843884e-10, 3.3693279180487663e-10, 
    3.3571500393013373e-10, 3.3452674917166183e-10, 3.3336146392777348e-10, 
    3.3221215067090101e-10, 3.3107181484735126e-10, 3.299338550344446e-10, 
    3.2879245171484613e-10, 3.2764286775975645e-10, 3.2648168844022876e-10, 
    3.2530694999118075e-10, 3.2411817032599119e-10, 3.2291625584636942e-10, 
    3.2170331590402054e-10, 3.2048235350425217e-10, 3.192569117670671e-10, 
    3.1803066022825747e-10, 3.1680699098421537e-10, 3.1558864893173427e-10, 
    3.1437745474247886e-10, 3.1317413835638639e-10, 3.1197832559277378e-10, 
    3.1078866202604775e-10, 3.0960308715754464e-10, 3.0841920889654789e-10, 
    3.072347532099591e-10, 3.060480082491018e-10, 3.0485823651952051e-10, 
    3.0366596432043723e-10, 3.0247314814478326e-10, 3.012831447154608e-10, 
    3.0010053308565935e-10, 2.9893074718036618e-10, 2.9777961552645845e-10, 
    2.9665280565224033e-10, 2.9555528284080088e-10, 2.9449078158201595e-10, 
    2.9346141622685038e-10, 2.9246740229357484e-10, 2.9150697336450323e-10, 
    2.9057645389012883e-10, 2.8967051826893414e-10, 2.8878257122034073e-10, 
    2.8790526821298668e-10, 2.8703105830804554e-10, 2.8615277450121164e-10, 
    2.8526417274672862e-10, 2.8436040207657014e-10, 2.8343835162658336e-10, 
    2.8249687254406105e-10, 2.8153682841497102e-10, 2.8056101286553326e-10, 
    2.795739035978275e-10, 2.7858132112045157e-10, 2.7758998356128471e-10, 
    2.7660704780568446e-10, 2.7563962484143426e-10, 2.746943661204922e-10, 
    2.7377710090379751e-10, 2.7289259566947796e-10, 2.7204438318227894e-10, 
    2.7123471593339858e-10, 2.7046455923879941e-10, 2.6973365442969284e-10, 
    2.6904056582277145e-10, 2.683827324896489e-10, 2.6775646167190977e-10, 
    2.6715690308541453e-10, 2.6657797464545317e-10, 2.6601231100803972e-10, 
    2.6545120673380173e-10, 2.6488466925727085e-10, 2.6430154192074491e-10, 
    2.6368978305841666e-10, 2.6303686152720953e-10, 2.623302992163657e-10, 
    2.6155829411337021e-10, 2.6071041574379089e-10, 2.5977828870076369e-10, 
    2.5875623795529002e-10, 2.5764179954731673e-10, 2.5643611286678894e-10, 
    2.5514409279614177e-10, 2.5377443308469824e-10, 2.5233939014524956e-10, 
    2.5085440211449117e-10, 2.4933751979951143e-10, 2.4780874685947429e-10, 
    2.4628924955883615e-10, 2.4480055933564357e-10, 2.4336372699337264e-10, 
    2.4199854662708502e-10, 2.4072281565311441e-10, 2.3955173184935956e-10, 
    2.3849738261777364e-10, 2.3756841462163007e-10, 2.3676982232192434e-10, 
    2.3610291372840166e-10, 2.3556538104041934e-10, 2.3515150763141057e-10, 
    2.3485242271218709e-10, 2.3465645091185671e-10, 2.3454945180375057e-10, 
    2.3451521688509811e-10, 2.3453584684395774e-10, 2.3459217548089358e-10, 
    2.3466419721536149e-10, 2.3473157295152595e-10, 2.347741511820707e-10, 
    2.3477258827837143e-10, 2.347089899193165e-10, 2.3456761424359319e-10, 
    2.3433553260675597e-10, 2.3400327809803973e-10, 2.3356536328209381e-10, 
    2.3302067269476292e-10, 2.323726343331564e-10, 2.3162919753182425e-10, 
    2.3080253068365777e-10, 2.2990851936888136e-10, 2.2896601067318103e-10, 
    2.2799591223403538e-10, 2.2702012524983418e-10, 2.2606044757716581e-10, 
    2.2513743822389346e-10, 2.2426937680125325e-10, 2.2347132650874178e-10, 
    2.2275440604518968e-10, 2.2212524437834386e-10, 2.2158574181617404e-10, 
    2.2113305399515413e-10, 2.2075987989619688e-10, 2.2045497322898499e-10, 
    2.2020390017205484e-10, 2.1998993685533745e-10, 2.1979512103845374e-10, 
    2.1960132741063284e-10, 2.1939136651070713e-10, 2.191499704142806e-10, 
    2.1886468514897204e-10, 2.1852653831020113e-10, 2.1813051059309473e-10, 
    2.1767571233877735e-10, 2.1716532823142304e-10, 2.1660625779863528e-10, 
    2.1600855211893343e-10, 2.1538461034551034e-10, 2.1474826102103663e-10, 
    2.1411374176691852e-10, 2.1349470285504018e-10, 2.1290324165590598e-10, 
    2.1234911936534397e-10, 2.1183914165908382e-10, 2.1137679815594807e-10, 
    2.1096213761034496e-10, 2.105919155341984e-10, 2.1025993554605341e-10, 
    2.0995760701867219e-10, 2.0967460666812991e-10, 2.0939963305059498e-10, 
    2.0912114277696651e-10, 2.0882806698971837e-10, 2.0851042128226017e-10, 
    2.0815981978734105e-10, 2.0776980651772681e-10, 2.0733608364658728e-10, 
    2.0685655542729543e-10, 2.0633127006313117e-10, 2.057622096231197e-10, 
    2.0515301399024488e-10, 2.04508605024211e-10, 2.0383478821265147e-10, 
    2.0313780335862562e-10, 2.0242390726248615e-10, 2.0169895182975568e-10, 
    2.0096804148541546e-10, 2.0023522728407736e-10, 1.9950331619763445e-10, 
    1.9877375469673768e-10, 1.9804664430880522e-10, 1.9732084999740863e-10, 
    1.9659425017609944e-10, 1.9586405366828611e-10, 1.9512724067256175e-10, 
    1.9438103543282336e-10, 1.9362343295475235e-10, 1.9285367229967509e-10, 
    1.9207267563351074e-10, 1.9128335901076308e-10, 1.9049081090214509e-10, 
    1.8970224375144557e-10, 1.8892679015752247e-10, 1.8817507234039812e-10, 
    1.8745863004862833e-10, 1.8678919411090664e-10, 1.8617794639064187e-10, 
    1.8563476227950671e-10, 1.851675801628961e-10, 1.8478190492798309e-10, 
    1.844805508847069e-10, 1.8426357971548558e-10, 1.8412849905980261e-10, 
    1.8407062121533006e-10, 1.8408357933796059e-10, 1.8415987733916699e-10, 
    1.8429144708535931e-10, 1.8447008857344312e-10, 1.8468780172353483e-10, 
    1.8493690571564115e-10, 1.8521002528138162e-10, 1.854998916490879e-10, 
    1.8579907225774821e-10, 1.8609962747383592e-10, 1.8639281966417898e-10, 
    1.8666888924003824e-10, 1.8691698910187737e-10, 1.8712525102810838e-10, 
    1.8728106758908608e-10, 1.8737150707176355e-10, 1.8738389007296125e-10, 
    1.8730642122841168e-10, 1.8712889826334665e-10, 1.8684336209528703e-10, 
    1.8644471392228279e-10, 1.8593118354919655e-10, 1.8530468644272624e-10, 
    1.845709629155321e-10, 1.8373957444226701e-10, 1.8282367575664982e-10, 
    1.8183964074721643e-10, 1.8080648320921692e-10, 1.7974517142709494e-10, 
    1.7867779609496862e-10, 1.7762668444386166e-10, 1.7661343893817567e-10, 
    1.756580053863399e-10, 1.7477776671523457e-10, 1.7398675682023434e-10, 
    1.7329498697117099e-10, 1.7270799522690529e-10, 1.7222659530189031e-10, 
    1.7184688555757343e-10, 1.7156051170780218e-10, 1.713551928341673e-10, 
    1.7121542455335421e-10, 1.711234065940415e-10, 1.7106003963073959e-10, 
    1.7100600105516604e-10, 1.7094274818351838e-10, 1.7085346439417205e-10, 
    1.7072380396340533e-10, 1.7054246976770264e-10, 1.7030153260154487e-10, 
    1.6999655474632409e-10, 1.6962646981504738e-10, 1.6919333205155072e-10, 
    1.6870190117996775e-10, 1.6815919063822162e-10, 1.6757397911391862e-10, 
    1.669563680057881e-10, 1.6631735764027566e-10, 1.6566853479506941e-10, 
    1.6502178573917439e-10, 1.6438907490334209e-10, 1.6378221192401667e-10, 
    1.6321262762808881e-10, 1.6269105001846459e-10, 1.6222714651747267e-10, 
    1.6182905888643002e-10, 1.6150290164201334e-10, 1.6125218644647675e-10, 
    1.6107732275294019e-10, 1.6097516968159578e-10, 1.6093878799841221e-10, 
    1.6095737364540269e-10, 1.6101651140740298e-10, 1.6109870629939974e-10, 
    1.611842391622619e-10, 1.6125224836337992e-10, 1.6128204516097384e-10, 
    1.6125449211040276e-10, 1.6115338322148182e-10, 1.6096665169678195e-10, 
    1.6068734677890911e-10, 1.6031421794042162e-10, 1.5985190130414775e-10, 
    1.5931062631126489e-10, 1.5870551570887964e-10, 1.5805546397555106e-10, 
    1.5738177452415339e-10, 1.5670658619408185e-10, 1.5605129919263842e-10, 
    1.5543507027671667e-10, 1.5487353416733255e-10, 1.5437781345384465e-10, 
    1.5395391412804802e-10, 1.5360246498084047e-10, 1.5331887154158487e-10, 
    1.5309376806061167e-10, 1.5291377120320028e-10, 1.5276238342874152e-10, 
    1.5262104546945812e-10, 1.5247019688922459e-10, 1.5229032605668601e-10, 
    1.5206290216800312e-10, 1.5177121990713002e-10, 1.5140106364340501e-10, 
    1.5094125020057474e-10, 1.50383982202836e-10, 1.4972509360866794e-10, 
    1.4896412668881673e-10, 1.4810432742627864e-10, 1.4715248839513856e-10, 
    1.4611874013917164e-10, 1.4501620799651699e-10, 1.4386062010997767e-10, 
    1.4266979292765668e-10, 1.4146307274744724e-10, 1.4026067051702792e-10, 
    1.3908297018036544e-10, 1.3794976388425563e-10, 1.368795162919183e-10, 
    1.3588860555958714e-10, 1.3499066216912604e-10, 1.3419599698076975e-10, 
    1.3351118672940289e-10, 1.3293881055434055e-10, 1.3247742252900102e-10, 
    1.321217026251381e-10, 1.3186283908235647e-10, 1.3168906463040604e-10, 
    1.3158637401997708e-10, 1.3153929201078897e-10, 1.3153172863107959e-10, 
    1.315477953294093e-10, 1.3157257062805923e-10, 1.3159273012489729e-10, 
    1.3159705127262759e-10, 1.3157671809491575e-10, 1.3152546636152367e-10, 
    1.3143951879592203e-10, 1.313173934884919e-10, 1.3115953357591623e-10, 
    1.3096787812468721e-10, 1.3074535067492911e-10, 1.304953617792999e-10, 
    1.3022133409510636e-10, 1.2992633310682066e-10, 1.2961278247056431e-10, 
    1.292823565480114e-10, 1.2893598871955873e-10, 1.2857404263591872e-10, 
    1.2819658566640022e-10, 1.2780375295004481e-10, 1.2739611639207981e-10, 
    1.2697504782406835e-10, 1.2654297754567527e-10, 1.2610354011282745e-10, 
    1.2566152662739183e-10, 1.2522268576790968e-10, 1.2479332727735092e-10, 
    1.2437980593511398e-10, 1.2398789482498632e-10, 1.2362216449397403e-10, 
    1.2328538537323039e-10, 1.2297808815308371e-10, 1.2269828396488108e-10, 
    1.224414368329649e-10, 1.2220068394437979e-10, 1.2196731327619236e-10, 
    1.2173142212174921e-10, 1.2148276612374574e-10, 1.2121165439824737e-10, 
    1.2090985983074455e-10, 1.2057140826228048e-10, 1.2019322205497234e-10, 
    1.1977550751126211e-10, 1.1932189575283465e-10, 1.1883928176942874e-10, 
    1.183374154577583e-10, 1.1782826512652585e-10, 1.1732521363052816e-10, 
    1.1684216500391012e-10, 1.163926465778668e-10, 1.1598894111602885e-10, 
    1.156413763809268e-10, 1.1535775745222895e-10, 1.1514302353544096e-10, 
    1.1499908997523832e-10, 1.1492492450364065e-10, 1.1491677844645405e-10, 
    1.1496858208313627e-10, 1.1507243545775052e-10, 1.152191666663086e-10, 
    1.1539888921383645e-10, 1.1560156149116012e-10, 1.1581745378715782e-10, 
    1.1603756536974969e-10, 1.1625391645074611e-10, 1.1645975710128272e-10, 
    1.1664964211047994e-10, 1.1681943854009989e-10, 1.1696622930960747e-10, 
    1.1708816330083213e-10, 1.1718427411456785e-10, 1.1725428424234337e-10, 
    1.172984076960634e-10, 1.1731720555669374e-10, 1.1731147179063589e-10, 
    1.1728219312144922e-10, 1.1723053967401127e-10, 1.171579255397354e-10, 
    1.1706609440559139e-10, 1.1695721715818531e-10, 1.1683397851141308e-10, 
    1.1669963187589883e-10, 1.1655800355628897e-10, 1.164134332547841e-10, 
    1.1627063551613977e-10, 1.1613450420762863e-10, 1.1600985594801796e-10, 
    1.1590114678842006e-10, 1.1581216366664378e-10, 1.1574574873065955e-10, 
    1.1570354898226734e-10, 1.1568584501850106e-10, 1.1569143248868904e-10, 
    1.1571761343482489e-10, 1.1576025636834428e-10, 1.158139358149241e-10, 
    1.1587214821401017e-10, 1.1592757016770725e-10, 1.1597235424283646e-10, 
    1.1599845176748036e-10, 1.1599794032069822e-10, 1.1596336275759453e-10, 
    1.1588804611292765e-10, 1.1576642998860606e-10, 1.1559435869354604e-10, 
    1.1536936683874137e-10, 1.1509091498515184e-10, 1.147605744567929e-10, 
    1.1438214386965135e-10, 1.139616617005692e-10, 1.1350730557876901e-10, 
    1.1302916025648384e-10, 1.1253884515592458e-10, 1.1204902009262198e-10, 
    1.1157276338592849e-10, 1.1112288993556748e-10, 1.1071123435108169e-10, 
    1.1034796152516144e-10, 1.1004094858192653e-10, 1.0979530303956889e-10, 
    1.0961306752589538e-10, 1.0949310441086972e-10, 1.0943120708167656e-10, 
    1.0942040570033518e-10, 1.0945142742082693e-10, 1.0951330082691214e-10, 
    1.0959401788614418e-10, 1.096812095435399e-10, 1.0976277980214006e-10, 
    1.0982745671030462e-10, 1.0986520233100229e-10, 1.0986749582830973e-10, 
    1.0982747308048548e-10, 1.097399373983926e-10, 1.0960125084540888e-10, 
    1.0940917775837794e-10, 1.0916267845147936e-10, 1.0886171138877154e-10, 
    1.0850705592303006e-10, 1.0810018538603153e-10, 1.0764318938458008e-10, 
    1.0713874662981093e-10, 1.0659012551435674e-10, 1.0600120239531403e-10, 
    1.0537646875802121e-10, 1.0472100702604781e-10, 1.0404041482811854e-10, 
    1.0334066719625162e-10, 1.0262792703289006e-10, 1.0190830248467809e-10, 
    1.0118756512353764e-10, 1.0047087690847284e-10, 9.9762533008930444e-11, 
    9.9065765367008875e-11, 9.8382633021682344e-11, 9.7714014826082228e-11, 
    9.7059729632222715e-11, 9.6418769958538156e-11, 9.5789635339051771e-11, 
    9.5170753708340783e-11, 9.4560922431548187e-11, 9.3959747591218341e-11, 
    9.3368018870305832e-11, 9.2787958716652811e-11, 9.2223339329433443e-11, 
    9.1679405169191173e-11, 9.1162607606148826e-11, 9.0680174196290723e-11, 
    9.0239530383983616e-11, 8.9847637102301864e-11, 8.9510293497982637e-11, 
    8.9231496509398768e-11, 8.9012901315893735e-11, 8.885345763186327e-11, 
    8.8749271599887565e-11, 8.8693695206313036e-11, 8.8677657918044667e-11, 
    8.8690219448724644e-11, 8.8719286957557492e-11, 8.8752452153669153e-11, 
    8.877787412112764e-11, 8.8785123684535662e-11, 8.8765945835475786e-11, 
    8.8714860742203544e-11, 8.8629561096325461e-11, 8.8511086681044766e-11, 
    8.8363751038762943e-11, 8.8194843047718646e-11, 8.8014104344957805e-11, 
    8.7833043481913771e-11, 8.7664119523401457e-11, 8.7519865452920242e-11, 
    8.7412002037043078e-11, 8.7350615225042512e-11, 8.7343452598333155e-11, 
    8.7395388788493379e-11, 8.7508096084587764e-11, 8.7679942636558889e-11, 
    8.7906116431148937e-11, 8.8178961324033129e-11, 8.8488489541648693e-11, 
    8.882302430973266e-11, 8.9169913100207654e-11, 8.9516252959792153e-11, 
    8.9849579344689872e-11, 9.0158458352969099e-11, 9.0432944366775061e-11, 
    9.0664889713465171e-11, 9.0848095728556405e-11, 9.0978306387063939e-11, 
    9.105305697035992e-11, 9.1071428666141923e-11, 9.1033733156303736e-11, 
    9.0941172200241352e-11, 9.079551985500135e-11, 9.0598870560029848e-11, 
    9.0353481755205653e-11, 9.0061742876219428e-11, 8.9726265041876619e-11, 
    8.935009942341599e-11, 8.8937029555149294e-11, 8.8491920850816697e-11, 
    8.802104572100818e-11, 8.7532332494818637e-11, 8.7035481204047983e-11, 
    8.6541890433881407e-11, 8.6064368359655906e-11, 8.5616642690548028e-11, 
    8.5212667258784467e-11, 8.4865810000807792e-11, 8.4587973821144871e-11, 
    8.4388738853120235e-11, 8.4274630598188747e-11, 8.4248564105900849e-11, 
    8.4309537221749779e-11, 8.4452611086788105e-11, 8.4669149847190625e-11, 
    8.4947328946664199e-11, 8.5272836057002492e-11, 8.5629702312541847e-11, 
    8.6001193104321095e-11, 8.637068130161751e-11, 8.6722427690378546e-11, 
    8.7042245083830026e-11, 8.7317980234451587e-11, 8.7539837840868738e-11, 
    8.7700517951435289e-11, 8.7795211662701762e-11, 8.78214751681693e-11, 
    8.7779008577370376e-11, 8.7669380528465502e-11, 8.7495730280041414e-11, 
    8.7262453414020148e-11, 8.6974917832447672e-11, 8.6639192854118818e-11, 
    8.6261829656564191e-11, 8.5849660029993844e-11, 8.5409642434196648e-11, 
    8.4948748489137257e-11, 8.4473883919670759e-11, 8.3991821785670825e-11, 
    8.3509178812028882e-11, 8.3032393216027537e-11, 8.2567711491203741e-11, 
    8.2121162835425104e-11, 8.1698518904442975e-11, 8.1305222716186891e-11, 
    8.0946286297566325e-11, 8.0626145770842531e-11, 8.0348505687887555e-11, 
    8.011614435301622e-11, 7.993074649260528e-11, 7.9792742086266559e-11, 
    7.9701202240445574e-11, 7.9653806923168309e-11, 7.9646893456174237e-11, 
    7.9675583118952895e-11, 7.9734009663517164e-11, 7.9815602324382919e-11, 
    7.9913428753169635e-11, 8.0020532032096271e-11, 8.0130276658669204e-11, 
    8.0236623226914907e-11, 8.0334338894859385e-11, 8.0419131574594629e-11, 
    8.0487683029467455e-11, 8.0537589642897682e-11, 8.0567260362129392e-11, 
    8.0575756100307954e-11, 8.0562635865828591e-11, 8.0527803799072883e-11, 
    8.0471415974374782e-11, 8.0393827636848046e-11, 8.0295613079068363e-11, 
    8.0177629130455529e-11, 8.0041128448501898e-11, 7.9887866926973766e-11, 
    7.9720216151709544e-11, 7.9541227235999432e-11, 7.9354643320571456e-11, 
    7.9164846745682275e-11, 7.8976753944091077e-11, 7.8795631550354804e-11, 
    7.8626920418147512e-11, 7.847602780663197e-11, 7.8348162696593575e-11, 
    7.824819584352468e-11, 7.8180588880192549e-11, 7.8149363750624268e-11, 
    7.8158126940672554e-11, 7.8210101063101829e-11, 7.8308160903209907e-11, 
    7.8454815584136265e-11, 7.8652156958982458e-11, 7.8901704902405886e-11, 
    7.9204209278794959e-11, 7.9559383180186737e-11, 7.9965626049346149e-11, 
    8.0419758398130437e-11, 8.0916829824307816e-11, 8.1450036205117859e-11, 
    8.2010783422407912e-11, 8.2588911483789617e-11, 8.3173091121974466e-11, 
    8.3751342182933908e-11, 8.4311665265826796e-11, 8.4842718459180682e-11, 
    8.5334473312142855e-11, 8.5778782023843075e-11, 8.6169823493249731e-11, 
    8.6504358965780483e-11, 8.6781791434638773e-11, 8.7004023845824978e-11, 
    8.717512742006496e-11, 8.730084701544539e-11, 8.7388013011526818e-11, 
    8.7443879032224146e-11, 8.7475472972610559e-11, 8.7488973153108774e-11, 
    8.7489190365179261e-11, 8.7479153426326044e-11, 8.7459845736690926e-11, 
    8.743008410603106e-11, 8.7386554472080812e-11, 8.7323991866017943e-11, 
    8.7235500111625853e-11, 8.7112983186298981e-11, 8.6947681199247395e-11, 
    8.673077609023203e-11, 8.6454042846680739e-11, 8.6110507318792399e-11, 
    8.5695075370636335e-11, 8.5205084958870986e-11, 8.4640755577358452e-11, 
    8.4005459828790602e-11, 8.3305822386683775e-11, 8.2551597215673063e-11, 
    8.1755327312861222e-11, 8.0931786270813745e-11, 8.009724721054499e-11, 
    7.9268627244467999e-11, 7.8462567268299038e-11, 7.7694527164689684e-11, 
    7.6977988012335645e-11, 7.6323810596614967e-11, 7.5739842538716548e-11, 
    7.523077081177493e-11, 7.4798258506679848e-11, 7.4441326352873395e-11, 
    7.4156936452772644e-11, 7.3940700775031498e-11, 7.3787648362656942e-11, 
    7.3692937765926843e-11, 7.3652466729551471e-11, 7.3663301803392792e-11, 
    7.3723896371737351e-11, 7.3834086425605594e-11, 7.3994871488717042e-11, 
    7.4208044466176184e-11, 7.4475697745487275e-11, 7.4799661332922174e-11, 
    7.5180969858748012e-11, 7.5619374504553672e-11, 7.611295551619785e-11, 
    7.6657861369379205e-11, 7.7248178165750774e-11, 7.7875932339243776e-11, 
    7.8531214054635256e-11, 7.9202392311806113e-11, 7.9876416146915289e-11, 
    8.0539180150122249e-11, 8.1175935432565646e-11, 8.1771733472441626e-11, 
    8.2311892569015377e-11, 8.278250048416942e-11, 8.3170912824482949e-11, 
    8.3466243582453044e-11, 8.3659838358657121e-11, 8.3745701256691529e-11, 
    8.3720840029137815e-11, 8.358549835652767e-11, 8.3343259017007332e-11, 
    8.3000973428735037e-11, 8.2568524881684984e-11, 8.205840801600465e-11, 
    8.148515157105456e-11, 8.0864600583984664e-11, 8.021312388875405e-11, 
    7.9546783824694531e-11, 7.8880540439272602e-11, 7.8227542291849806e-11, 
    7.7598563455965011e-11, 7.7001623490389934e-11, 7.6441813669903337e-11, 
    7.592133539610501e-11, 7.5439740565785922e-11, 7.4994337422567691e-11, 
    7.458072344205213e-11, 7.4193408819314584e-11, 7.3826454002276647e-11, 
    7.3474088889248834e-11, 7.3131263760968794e-11, 7.2794083029876613e-11, 
    7.246011656995734e-11, 7.2128547641031495e-11, 7.1800171274321786e-11, 
    7.1477244024699607e-11, 7.1163202701780784e-11, 7.0862289926006618e-11, 
    7.0579110699252846e-11, 7.031817702729286e-11, 7.0083468037586613e-11, 
    6.9878062804090332e-11, 6.9703862883495426e-11, 6.9561434941159785e-11, 
    6.9449989038873809e-11, 6.9367477642746813e-11, 6.9310815430789746e-11, 
    6.9276179493181266e-11, 6.9259371949419845e-11, 6.9256200904424902e-11, 
    6.9262852342189737e-11, 6.9276218956448786e-11, 6.9294160454176386e-11, 
    6.9315695966389063e-11, 6.9341095523107916e-11, 6.9371886643785292e-11, 
    6.9410770598219088e-11, 6.9461452746695923e-11, 6.952839198999169e-11, 
    6.961649347256796e-11, 6.9730732694798728e-11, 6.9875740171818446e-11, 
    7.0055364835260526e-11, 7.0272236494271388e-11, 7.052735861394741e-11, 
    7.0819746696313534e-11, 7.1146163142628488e-11, 7.1500969151478544e-11, 
    7.1876107907900978e-11, 7.2261243678589937e-11, 7.2644052942304295e-11, 
    7.3010665929911408e-11, 7.3346233680382847e-11, 7.3635589105755374e-11, 
    7.3863977535587083e-11, 7.4017794423287991e-11, 7.4085308954909854e-11, 
    7.4057328063436852e-11, 7.392774828318809e-11, 7.3693998365933252e-11, 
    7.3357322677843917e-11, 7.2922900442467219e-11, 7.2399798759327804e-11, 
    7.1800748716467495e-11, 7.1141753979193775e-11, 7.0441545982867311e-11, 
    6.9720892323310047e-11, 6.9001794887158027e-11, 6.8306590502639663e-11, 
    6.7657005666585447e-11, 6.7073192730295095e-11, 6.6572803749784636e-11, 
    6.6170147976612073e-11, 6.5875480902285276e-11, 6.5694473672765714e-11, 
    6.5627898711288006e-11, 6.5671559634810978e-11, 6.5816475995446054e-11, 
    6.6049318570808261e-11, 6.6353069903092208e-11, 6.670787092083194e-11, 
    6.7092015012563831e-11, 6.7483014425773362e-11, 6.7858692177274789e-11, 
    6.8198241229005308e-11, 6.8483191311040389e-11, 6.8698253658952444e-11, 
    6.8832004350400832e-11, 6.8877383640830062e-11,
  // Sqw-Na(8, 0-1999)
    0.020925215872861367, 0.020922136582194942, 0.020912976261888948, 
    0.02089796201066935, 0.020877454249665642, 0.020851921129086196, 
    0.020821905620903317, 0.020787987944837723, 0.020750746350248629, 
    0.020710719392985747, 0.020668372681704367, 0.020624072625821877, 
    0.020578069029855164, 0.020530487508854518, 0.020481331735432057, 
    0.020430494575874994, 0.020377776340797994, 0.020322907763955265, 
    0.020265575005350811, 0.020205443988933789, 0.020142181724551411, 
    0.020075472878059154, 0.020005030654493345, 0.019930601933570529, 
    0.019851967422020715, 0.019768938249741987, 0.019681350848102505, 
    0.019589062058471322, 0.019491946221372344, 0.019389895530245636, 
    0.01928282427521787, 0.019170676853795705, 0.01905343869948237, 
    0.018931148682246907, 0.018803911151723713, 0.018671905677856249, 
    0.018535392708736113, 0.018394713786776744, 0.018250285582746953, 
    0.018102587737787605, 0.017952145248122733, 0.017799506787416288, 
    0.017645220852060862, 0.017489811873326547, 0.017333758436939548, 
    0.017177475490083107, 0.017021301936812325, 0.016865494392647461, 
    0.016710227173694504, 0.016555597927663705, 0.016401637759529648, 
    0.0162483243302411, 0.016095596251374165, 0.015943367167191004, 
    0.015791538180644021, 0.015640007686814731, 0.015488678154409298, 
    0.01533745986704285, 0.01518627203299888, 0.015035041945497462, 
    0.01488370300099259, 0.014732192363284357, 0.014580448922463716, 
    0.014428411982445473, 0.014276020868435739, 0.014123215422591477, 
    0.013969937187864387, 0.013816130986144771, 0.013661746579677288, 
    0.013506740151691742, 0.013351075430639849, 0.013194724385945487, 
    0.013037667517712336, 0.012879893831429061, 0.012721400623912929, 
    0.012562193210516675, 0.012402284705047586, 0.012241695935277392, 
    0.012080455549864835, 0.011918600354164834, 0.011756175903754289, 
    0.011593237380483127, 0.01142985076734631, 0.011266094315710977, 
    0.011102060254786451, 0.010937856628304342, 0.010773609064506594, 
    0.010609462207189002, 0.010445580476563859, 0.01028214780813025, 
    0.010119366050018964, 0.0099574517902049908, 0.0097966315293324027, 
    0.0096371352964382123, 0.0094791889988292289, 0.0093230059748795318, 
    0.0091687783519497097, 0.0090166688797862979, 0.0088668039016710828, 
    0.0087192680422230971, 0.0085741010443711255, 0.0084312969994053081, 
    0.0082908060084532081, 0.0081525381164581669, 0.0080163691920550131, 
    0.0078821483033071973, 0.0077497060670331103, 0.0076188634280949007, 
    0.0074894403485927146, 0.0073612639459730914, 0.0072341757028867035, 
    0.0071080374698669554, 0.0069827360855106947, 0.0068581865403967148, 
    0.0067343337043843359, 0.0066111527170695421, 0.0064886482036050647, 
    0.0063668525191906819, 0.0062458232429626632, 0.0061256401354401729, 
    0.0060064017455174167, 0.0058882218087135804, 0.0057712255263083134, 
    0.0056555457652349593, 0.0055413191814705541, 0.005428682253587923, 
    0.0053177672227190586, 0.00520869796979393, 0.0051015859142718939, 
    0.004996526079540666, 0.004893593524694196, 0.0047928403764315591, 
    0.0046942936972576461, 0.0045979543915723349, 0.0045037972813621596, 
    0.0044117723870630366, 0.0043218073414266062, 0.0042338107623889369, 
    0.0041476763317068004, 0.0040632872819197433, 0.0039805209905696762, 
    0.0038992534151757372, 0.0038193631655548278, 0.0037407350870425462, 
    0.0036632633026770067, 0.0035868537200823359, 0.0035114260402459184, 
    0.0034369153080751531, 0.0033632730230464271, 0.0032904677926264216, 
    0.0032184854747797278, 0.0031473287320849591, 0.003077015919020367, 
    0.003007579250838833, 0.002939062255810347, 0.0028715165851832588, 
    0.0028049983352582035, 0.0027395641096234695, 0.0026752671035118105, 
    0.0026121535159804609, 0.002550259583440104, 0.0024896094797832035, 
    0.0024302142492400509, 0.0023720718378610096, 0.0023151681807808957, 
    0.0022594791987083787, 0.0022049734709378536, 0.0021516152934922686, 
    0.0020993678058233755, 0.0020481958794690046, 0.0019980685044697559, 
    0.0019489604776977978, 0.0019008532823374875, 0.001853735138962635, 
    0.0018076002953361877, 0.001762447694861069, 0.0017182792155101727, 
    0.0016750976980544003, 0.0016329049837515688, 0.0015917001597083944, 
    0.0015514781697468379, 0.0015122288963274921, 0.001473936762091844, 
    0.0014365808447365106, 0.0014001354518830985, 0.0013645710672461847, 
    0.0013298555575774812, 0.0012959555214735554, 0.0012628376644759759, 
    0.0012304700972297186, 0.0011988234716382822, 0.0011678718909642432, 
    0.0011375935512483294, 0.0011079710916419342, 0.001078991649455705, 
    0.0010506466317540797, 0.0010229312293677404, 0.00099584371151746794, 
    0.00096938454992107135, 0.00094355543005321613, 0.00091835821357743295, 
    0.00089379391910525592, 0.00086986178758536551, 0.00084655849325570014, 
    0.00082387755110503735, 0.00080180895765929257, 0.00078033908467161923, 
    0.0007594508264721591, 0.00073912398310298721, 0.00071933584472621312, 
    0.00070006192969028936, 0.00068127682015302956, 0.00066295503576540389, 
    0.00064507188747724912, 0.00062760425934505143, 0.00061053127524106701, 
    0.00059383481834284521, 0.00057749988302483, 0.0005615147502743285, 
    0.00054587098830676396, 0.00053056328925533503, 0.00051558916050868414, 
    0.00050094849546379833, 0.00048664305319353241, 0.0004726758797915863, 
    0.00045905070586804741, 0.00044577135466621011, 0.00043284119339725638, 
    0.00042026265655769002, 0.00040803686428897515, 0.00039616335155305879, 
    0.00038463991555313519, 0.000373462580118752, 0.00036262566748556985, 
    0.00035212196079493406, 0.00034194293535670179, 0.00033207903368330581, 
    0.00032251995868461374, 0.00031325496111520186, 0.00030427310106677271, 
    0.00029556346849766952, 0.00028711535388409169, 0.00027891836640943856, 
    0.00027096250304212339, 0.00026323817680624234, 0.00025573621604965024, 
    0.00024844784822520839, 0.00024136468147439605, 0.0002344786951994472, 
    0.00022778224712759879, 0.00022126809962271985, 0.00021492946288193139, 
    0.00020876004795418156, 0.00020275411900782939, 0.00019690653257791859, 
    0.0001912127520047324, 0.00018566882794415155, 0.00018027134032841673, 
    0.00017501730278740926, 0.00016990403639079003, 0.00016492902465482836, 
    0.00016008976520440256, 0.00015538363468753063, 0.0001508077822913499, 
    0.00014635906370642933, 0.00014203402221565645, 0.00013782891758948947, 
    0.00013373979760232028, 0.0001297626021191161, 0.00012589328648989132, 
    0.00012212794975555684, 0.00011846295388449112, 0.00011489502257940887, 
    0.000111421311561227, 0.00010803944600358237, 0.00010474752436136227, 
    0.0001015440907605211, 9.8428080162397852e-05, 9.5398741668118356e-05, 
    9.2455545753902297e-05, 8.9598081191851045e-05, 8.6825947198450679e-05, 
    8.4138646180933333e-05, 8.1535482423967308e-05, 7.9015472141760897e-05, 
    7.6577270370076285e-05, 7.4219119976573654e-05, 7.1938827418661759e-05, 
    6.9733768627874718e-05, 6.7600926517912661e-05, 6.5536959201249262e-05, 
    6.3538295290162182e-05, 6.1601249976358889e-05, 5.9722153296098568e-05, 
    5.789748043418866e-05, 5.6123973360092604e-05, 5.4398743649455345e-05, 
    5.2719348002761883e-05, 5.1083830553905259e-05, 4.9490729267591718e-05, 
    4.793904717413461e-05, 4.6428192479107377e-05, 4.4957894336369959e-05, 
    4.3528102993026177e-05, 4.2138883922973121e-05, 4.0790315418247769e-05, 
    3.9482397988792183e-05, 3.8214982030779419e-05, 3.6987717836004265e-05, 
    3.580002944448992e-05, 3.4651111395181163e-05, 3.3539945370605704e-05, 
    3.2465332249627416e-05, 3.1425934281082063e-05, 3.0420321976706774e-05, 
    2.9447020820349176e-05, 2.8504553858078148e-05, 2.7591477489315638e-05, 
    2.6706409123569537e-05, 2.584804661806688e-05, 2.5015180417066822e-05, 
    2.4206699976424071e-05, 2.3421596334715523e-05, 2.2658962604180423e-05, 
    2.1917993767064923e-05, 2.1197986581307044e-05, 2.0498339744381289e-05, 
    1.981855385822342e-05, 1.9158230282184538e-05, 1.8517067726569699e-05, 
    1.7894855454869768e-05, 1.7291462218606191e-05, 1.6706820496133901e-05, 
    1.6140906173930917e-05, 1.5593714408366565e-05, 1.5065232953433933e-05, 
    1.455541466082582e-05, 1.4064151102136394e-05, 1.3591249300800694e-05, 
    1.3136413394460371e-05, 1.2699232697873286e-05, 1.2279177144960469e-05, 
    1.1875600507281397e-05, 1.1487751175685217e-05, 1.1114789708765751e-05, 
    1.0755811850575971e-05, 1.0409875342229852e-05, 1.0076028628732639e-05, 
    9.7533395060207237e-06, 9.4409218622938895e-06, 9.1379589218492411e-06, 
    8.8437217669420049e-06, 8.5575823494983233e-06, 8.2790206637213696e-06, 
    8.0076261854800125e-06, 7.7430940578647821e-06, 7.4852167862231792e-06, 
    7.2338723893195101e-06, 6.9890100360969767e-06, 6.7506341947592316e-06, 
    6.518788251933421e-06, 6.2935384495141583e-06, 6.0749588556272378e-06, 
    5.8631179511604139e-06, 5.6580672819607203e-06, 5.4598325023908745e-06, 
    5.2684070140443283e-06, 5.0837482808212221e-06, 4.9057767733620888e-06, 
    4.7343773638147314e-06, 4.5694028600819145e-06, 4.410679248047705e-06, 
    4.2580121121683474e-06, 4.1111936431870736e-06, 3.9700096249697048e-06, 
    3.8342458269144988e-06, 3.7036933109967006e-06, 3.5781522868456792e-06, 
    3.4574343001070167e-06, 3.34136270429945e-06, 3.2297715268186411e-06, 
    3.1225029825430351e-06, 3.0194040011192274e-06, 2.9203222105014394e-06, 
    2.8251018549532234e-06, 2.7335801217282439e-06, 2.6455843076148147e-06, 
    2.5609301799725601e-06, 2.4794217804550673e-06, 2.4008527916354095e-06, 
    2.3250094444445827e-06, 2.2516747996866728e-06, 2.1806341010282683e-06, 
    2.1116807845122231e-06, 2.0446226523183902e-06, 1.9792876878842941e-06, 
    1.9155290101180663e-06, 1.8532285374823497e-06, 1.7922990499408417e-06, 
    1.7326844862789669e-06, 1.6743584772163858e-06, 1.6173212723948864e-06, 
    1.5615953520356869e-06, 1.5072201083155266e-06, 1.4542460278189985e-06, 
    1.402728804879288e-06, 1.3527237710931892e-06, 1.3042809513807652e-06, 
    1.2574409649473898e-06, 1.2122318962436095e-06, 1.1686671773843181e-06, 
    1.1267444586377388e-06, 1.0864453989721666e-06, 1.0477362833355031e-06, 
    1.010569360814153e-06, 9.7488479230041196e-07, 9.4061309025645192e-07, 
    9.0767792400462064e-07, 8.759991496462414e-07, 8.4549590815447083e-07, 
    8.1608962201920949e-07, 7.877067173225438e-07, 7.6028090794383816e-07, 
    7.3375490586403128e-07, 7.0808146442276573e-07, 6.8322371697133263e-07, 
    6.5915483397129684e-07, 6.3585707971497783e-07, 6.1332039654572215e-07, 
    5.9154067429837585e-07, 5.705178712196779e-07, 5.5025414130014415e-07, 
    5.3075209415604161e-07, 5.1201327492661191e-07, 4.940369093528518e-07, 
    4.7681892196932318e-07, 4.6035120759509374e-07, 4.4462112250536306e-07, 
    4.2961116064542647e-07, 4.1529879072726505e-07, 4.0165644594315338e-07, 
    3.8865167512645611e-07, 3.7624747596350956e-07, 3.6440283450535724e-07, 
    3.530734881114541e-07, 3.4221291258733738e-07, 3.3177351054681412e-07, 
    3.2170795223999087e-07, 3.1197059587750342e-07, 3.025188974235366e-07, 
    2.9331471192868937e-07, 2.8432539216967618e-07, 2.7552460416832169e-07, 
    2.6689280207109675e-07, 2.5841733263722126e-07, 2.5009216976388191e-07, 
    2.419173076173595e-07, 2.338978654269921e-07, 2.2604297502136984e-07, 
    2.1836453402513865e-07, 2.1087591205920804e-07, 2.0359069594361706e-07, 
    1.9652155234455496e-07, 1.8967927439200023e-07, 1.8307206245983791e-07, 
    1.7670507034352531e-07, 1.7058022682703337e-07, 1.6469632142003134e-07, 
    1.5904932258776232e-07, 1.5363287998928548e-07, 1.4843894966062672e-07, 
    1.4345847522912764e-07, 1.3868205864012839e-07, 1.3410056142699647e-07, 
    1.2970559013166167e-07, 1.2548983622365964e-07, 1.2144725856430814e-07, 
    1.1757311361119455e-07, 1.1386385226811056e-07, 1.1031691200619656e-07, 
    1.0693043719265894e-07, 1.0370296073680959e-07, 1.0063307620828921e-07, 
    9.7719124025229581e-08, 9.4958908590467562e-08, 9.2349457776347815e-08, 
    8.9886831667130798e-08, 8.7565985216457036e-08, 8.5380688181748252e-08, 
    8.3323505694080161e-08, 8.1385842189805956e-08, 7.9558050585429786e-08, 
    7.7829605880588289e-08, 7.6189339032454935e-08, 7.4625722019694581e-08, 
    7.3127190489451627e-08, 7.1682485782609268e-08, 7.0280995461637086e-08, 
    6.8913070161417116e-08, 6.757029586445447e-08, 6.6245703634055927e-08, 
    6.4933903815927326e-08, 6.363113719276305e-08, 6.2335241928027848e-08, 
    6.1045540522771981e-08, 5.9762656195835989e-08, 5.8488271586746027e-08, 
    5.722484554271881e-08, 5.5975305073909393e-08, 5.4742730491377255e-08, 
    5.3530051468876818e-08, 5.2339771420478246e-08, 5.1173736129757997e-08, 
    5.0032960869986993e-08, 4.8917527221086227e-08, 4.7826557203654345e-08, 
    4.6758267275086566e-08, 4.5710099286171165e-08, 4.4678919137995276e-08, 
    4.3661268071230748e-08, 4.265364618881973e-08, 4.1652804444817353e-08, 
    4.0656019721834701e-08, 3.9661329017361511e-08, 3.8667702193057143e-08, 
    3.7675138888340914e-08, 3.6684682354665425e-08, 3.5698351180352263e-08, 
    3.4718997267694271e-08, 3.3750104959528109e-08, 3.2795550320921712e-08, 
    3.1859341829619234e-08, 3.0945363217777488e-08, 3.0057137198880884e-08, 
    2.9197624946055394e-08, 2.8369072093416184e-08, 2.7572907399599686e-08, 
    2.6809696467691329e-08, 2.6079149423491992e-08, 2.5380179171394523e-08, 
    2.4711004695993493e-08, 2.406929258313822e-08, 2.3452328299670442e-08, 
    2.2857207641258281e-08, 2.2281037121369304e-08, 2.1721131152650632e-08, 
    2.1175192907697329e-08, 2.0641466158904399e-08, 2.0118846359299204e-08, 
    1.9606941928572954e-08, 1.9106080146462325e-08, 1.8617256818765859e-08, 
    1.8142033543016165e-08, 1.7682391384817482e-08, 1.7240553442327562e-08, 
    1.6818791631941331e-08, 1.6419233748676703e-08, 1.6043686389882774e-08, 
    1.5693486814107426e-08, 1.536939356776229e-08, 1.5071521364232873e-08, 
    1.479932166256156e-08, 1.4551606197369991e-08, 1.4326607735556559e-08, 
    1.4122069834681284e-08, 1.3935356408434565e-08, 1.376357140578383e-08, 
    1.3603679729890775e-08, 1.3452621574234182e-08, 1.3307414243149484e-08, 
    1.3165237231470833e-08, 1.3023498560387454e-08, 1.2879881992113097e-08, 
    1.2732376641130853e-08, 1.2579291509080699e-08, 1.2419258459003458e-08, 
    1.2251227216433607e-08, 1.2074455871344527e-08, 1.1888499395193075e-08, 
    1.1693197844545583e-08, 1.1488664423546037e-08, 1.1275272743831378e-08, 
    1.1053641524946243e-08, 1.08246149164653e-08, 1.0589236596008459e-08, 
    1.0348716797113871e-08, 1.0104392297059684e-08, 9.857680948936836e-09, 
    9.6100332618498598e-09, 9.362884603308493e-09, 9.1176116398236655e-09, 
    8.8754965528636649e-09, 8.637701423488725e-09, 8.4052541001804327e-09, 
    8.1790451671123985e-09, 7.9598344426971987e-09, 7.7482641680343836e-09, 
    7.5448756370991902e-09, 7.3501258562685815e-09, 7.1644014677460684e-09, 
    6.9880279123834596e-09, 6.8212731071026696e-09, 6.6643458258066872e-09, 
    6.517390085501031e-09, 6.3804772784649862e-09, 6.2535981774390353e-09, 
    6.1366566236485233e-09, 6.029466437581355e-09, 5.9317522343434407e-09, 
    5.8431543691307224e-09, 5.7632373778165467e-09, 5.691501007122975e-09, 
    5.6273925019137799e-09, 5.5703190127687358e-09, 5.5196589616364249e-09, 
    5.4747717666949014e-09, 5.4350055282269574e-09, 5.3997029113860203e-09, 
    5.3682055630956909e-09, 5.339857847089711e-09, 5.3140105169068948e-09, 
    5.2900251024694471e-09, 5.2672793521407184e-09, 5.2451740387125763e-09, 
    5.2231408930285897e-09, 5.2006513507188938e-09, 5.1772253230085255e-09, 
    5.1524392930257613e-09, 5.1259327555732575e-09, 5.0974123195967905e-09, 
    5.0666527868433716e-09, 5.0334950331219207e-09, 4.9978406889514569e-09, 
    4.9596442119796409e-09, 4.9189031215453151e-09, 4.875647622552403e-09, 
    4.8299308166910997e-09, 4.7818208299568672e-09, 4.7313957907685129e-09, 
    4.6787424142614588e-09, 4.62395825728915e-09, 4.5671573644170378e-09, 
    4.5084783416495472e-09, 4.4480936966062298e-09, 4.386218858317032e-09, 
    4.3231195055742635e-09, 4.2591157759569838e-09, 4.1945825208607735e-09, 
    4.1299450204317526e-09, 4.0656702848810514e-09, 4.0022543550711168e-09, 
    3.9402065943929179e-09, 3.8800320134405369e-09, 3.8222129845225742e-09, 
    3.7671914712071405e-09, 3.7153529284407575e-09, 3.667012613923742e-09, 
    3.6224050134472512e-09, 3.5816766049343848e-09, 3.5448821953197014e-09, 
    3.5119846569994203e-09, 3.4828580067426038e-09, 3.4572934605372959e-09, 
    3.4350082137267305e-09, 3.4156565003979399e-09, 3.3988425532396448e-09, 
    3.3841349096376586e-09, 3.3710815875367613e-09, 3.3592254791635115e-09, 
    3.3481194265461698e-09, 3.3373403013439159e-09, 3.3265016348067148e-09, 
    3.3152642535501075e-09, 3.3033446397487264e-09, 3.2905207136388994e-09, 
    3.2766350363777271e-09, 3.2615953589188009e-09, 3.245372754740321e-09, 
    3.2279974353862022e-09, 3.2095526337945404e-09, 3.1901667724591061e-09, 
    3.1700043642475108e-09, 3.1492559093642072e-09, 3.1281273289279081e-09, 
    3.1068292353420939e-09, 3.0855665819315769e-09, 3.0645290498098945e-09, 
    3.0438826590427319e-09, 3.0237628749263028e-09, 3.004269578206496e-09, 
    2.985463959115459e-09, 2.967367475354096e-09, 2.9499626611962457e-09, 
    2.9331956886569753e-09, 2.9169802831854316e-09, 2.9012027028445462e-09, 
    2.8857273414509938e-09, 2.8704026956707811e-09, 2.8550673220610572e-09, 
    2.8395556707682787e-09, 2.823703585715497e-09, 2.8073535046194978e-09, 
    2.7903592563377123e-09, 2.7725905662951785e-09, 2.7539371338370675e-09, 
    2.7343123567943228e-09, 2.713656491324397e-09, 2.691939197867618e-09, 
    2.6691612257841911e-09, 2.6453551303970207e-09, 2.6205848228455725e-09, 
    2.5949439358831067e-09, 2.5685529320147636e-09, 2.5415551204383079e-09, 
    2.5141116735249366e-09, 2.486395969422178e-09, 2.458587485913921e-09, 
    2.4308656315094976e-09, 2.4034037481044897e-09, 2.376363666765394e-09, 
    2.3498909702675388e-09, 2.3241112419551897e-09, 2.2991273376109463e-09, 
    2.275017857982271e-09, 2.2518367507803901e-09, 2.2296140853521544e-09, 
    2.2083578402923193e-09, 2.1880566705010674e-09, 2.1686833757021786e-09, 
    2.150198955129131e-09, 2.132556908950434e-09, 2.1157075905490239e-09, 
    2.0996022180752182e-09, 2.0841963653911118e-09, 2.069452564327373e-09, 
    2.0553419124460447e-09, 2.0418444654656717e-09, 2.0289484746153156e-09, 
    2.0166484665040759e-09, 2.0049424356635793e-09, 1.9938283470358506e-09, 
    1.9833003833403245e-09, 1.9733452452959154e-09, 1.9639389488608559e-09, 
    1.9550443883819696e-09, 1.9466099777096573e-09, 1.9385694693753399e-09, 
    1.9308430399752766e-09, 1.92333950551074e-09, 1.9159595728871255e-09, 
    1.9085997877140979e-09, 1.9011569653165208e-09, 1.8935326870998572e-09, 
    1.8856376328538597e-09, 1.8773953660423908e-09, 1.868745411485904e-09, 
    1.8596453681029884e-09, 1.8500720234752793e-09, 1.8400213679707174e-09, 
    1.829507625988131e-09, 1.8185613487181215e-09, 1.8072268032814029e-09, 
    1.7955587952680961e-09, 1.7836192223499826e-09, 1.7714735147395336e-09, 
    1.7591872411197984e-09, 1.7468229890661028e-09, 1.7344377328935941e-09, 
    1.7220807254287787e-09, 1.7097920313104062e-09, 1.6976016438639698e-09, 
    1.6855292796262171e-09, 1.6735847121076463e-09, 1.6617686864988653e-09, 
    1.650074265530201e-09, 1.6384886049144684e-09, 1.6269949888066649e-09, 
    1.6155750959780082e-09, 1.6042112808409795e-09, 1.5928888450145813e-09, 
    1.5815980610227905e-09, 1.570335900298104e-09, 1.5591072755444163e-09, 
    1.5479257651522249e-09, 1.5368137000052602e-09, 1.5258016470771043e-09, 
    1.5149272650573114e-09, 1.5042336617158673e-09, 1.4937672877917725e-09, 
    1.4835756031995691e-09, 1.4737045924322602e-09, 1.4641963727097685e-09, 
    1.4550869764315999e-09, 1.446404521521566e-09, 1.4381677950524548e-09, 
    1.4303853810162823e-09, 1.4230552747490659e-09, 1.4161650365863881e-09, 
    1.409692362284694e-09, 1.4036060533637714e-09, 1.397867228582511e-09, 
    1.3924307653789791e-09, 1.387246807440575e-09, 1.3822623458381291e-09, 
    1.3774227610671665e-09, 1.3726733538194306e-09, 1.3679607736793221e-09, 
    1.363234415631333e-09, 1.3584476820011726e-09, 1.3535591685579362e-09, 
    1.3485336801832227e-09, 1.3433430910988476e-09, 1.3379669534459794e-09, 
    1.3323928613719604e-09, 1.3266164629958235e-09, 1.3206411728148517e-09, 
    1.3144774919462813e-09, 1.308142037021863e-09, 1.301656256317568e-09, 
    1.295044972350372e-09, 1.2883347822499166e-09, 1.2815524957660766e-09, 
    1.2747236652693466e-09, 1.267871377565404e-09, 1.2610153231361611e-09, 
    1.2541712950417547e-09, 1.2473510546372479e-09, 1.2405626287364215e-09, 
    1.2338109251185658e-09, 1.2270986406867981e-09, 1.2204272977185952e-09, 
    1.2137983513485469e-09, 1.2072141687771121e-09, 1.2006788567707815e-09, 
    1.1941987568147001e-09, 1.1877826395167623e-09, 1.1814414860536837e-09, 
    1.1751879612533151e-09, 1.1690355479545949e-09, 1.1629975048895856e-09, 
    1.1570856707192647e-09, 1.1513093199356287e-09, 1.1456741082943382e-09, 
    1.1401812984548306e-09, 1.1348272689002677e-09, 1.1296034529555469e-09, 
    1.1244966573690811e-09, 1.1194898086893437e-09, 1.1145630093067975e-09, 
    1.1096948996991803e-09, 1.104864138133253e-09, 1.1000509519389763e-09, 
    1.0952385652450576e-09, 1.0904144633608623e-09, 1.0855713227799606e-09, 
    1.08070760818285e-09, 1.075827734535557e-09, 1.0709418364896777e-09, 
    1.0660651080857173e-09, 1.0612168274499154e-09, 1.0564190515234374e-09, 
    1.0516951501398823e-09, 1.047068177077869e-09, 1.0425592697179842e-09, 
    1.0381860925578309e-09, 1.0339614886789603e-09, 1.0298923503750089e-09, 
    1.0259788695573148e-09, 1.0222141188892194e-09, 1.0185841009291268e-09, 
    1.0150681724875836e-09, 1.0116399155377354e-09, 1.0082683272560766e-09, 
    1.0049193369992371e-09, 1.0015574781134595e-09, 9.981476878292733e-10, 
    9.9465705466234567e-10, 9.9105646140736699e-10, 9.8732194287430107e-10, 
    9.8343575928558024e-10, 9.7938701515541825e-10, 9.7517188631247184e-10, 
    9.707933403120573e-10, 9.6626046539229644e-10, 9.6158738497888044e-10, 
    9.567919152924887e-10, 9.5189397135375181e-10, 9.4691396557655065e-10, 
    9.4187121045229242e-10, 9.3678255231075751e-10, 9.316612462522182e-10, 
    9.2651626786725257e-10, 9.213520090365088e-10, 9.1616847354103184e-10, 
    9.1096186873102717e-10, 9.0572561964941352e-10, 9.0045160857811837e-10, 
    8.9513164715717576e-10, 8.8975893997175196e-10, 8.8432950244513734e-10, 
    8.7884331538269575e-10, 8.7330521232923051e-10, 8.6772532600732155e-10, 
    8.6211914412295129e-10, 8.5650707819178204e-10, 8.5091365979002049e-10, 
    8.4536635024429551e-10, 8.3989412970923854e-10, 8.3452588738841504e-10, 
    8.2928881075869338e-10, 8.2420682720258698e-10, 8.1929925203449892e-10, 
    8.1457968022283255e-10, 8.1005526473349036e-10, 8.0572633286992904e-10, 
    8.0158646244243384e-10, 7.976229030782484e-10, 7.9381741595938239e-10, 
    7.9014737766228886e-10, 7.8658718066041957e-10, 7.8310973529089528e-10, 
    7.7968809092367608e-10, 7.7629696873025557e-10, 7.7291421049558387e-10, 
    7.6952193342764079e-10, 7.6610743112975199e-10, 7.6266364715019845e-10, 
    7.5918928466702905e-10, 7.5568845278405122e-10, 7.5216996721071272e-10, 
    7.4864628176757689e-10, 7.4513221648477331e-10, 7.4164352111435342e-10, 
    7.3819546361190724e-10, 7.3480148137713284e-10, 7.3147209374998491e-10, 
    7.2821407136731182e-10, 7.2502999797838602e-10, 7.2191816016051553e-10, 
    7.188728393548028e-10, 7.1588487385513004e-10, 7.1294250160093259e-10, 
    7.1003230769212652e-10, 7.0714027365594378e-10, 7.0425275197814378e-10, 
    7.0135735528797574e-10, 6.9844361857088162e-10, 6.955034640057363e-10, 
    6.9253137918767476e-10, 6.8952437031743949e-10, 6.8648164247209322e-10, 
    6.8340415098007628e-10, 6.8029396542573365e-10, 6.7715364372198909e-10, 
    6.7398559356582835e-10, 6.7079157363821845e-10, 6.6757233958560979e-10, 
    6.6432754522461629e-10, 6.6105585305821764e-10, 6.5775533541577315e-10, 
    6.5442403466590029e-10, 6.5106071663229091e-10, 6.476656442036287e-10, 
    6.4424134970655556e-10, 6.4079322238529481e-10, 6.3732990465429444e-10, 
    6.3386334307889777e-10, 6.3040853392544026e-10, 6.2698288124032057e-10, 
    6.2360529435429228e-10, 6.2029501615568727e-10, 6.170703694924637e-10, 
    6.1394744596996256e-10, 6.109389564478512e-10, 6.0805327760809685e-10, 
    6.0529383389731914e-10, 6.0265880561881073e-10, 6.0014126572357914e-10, 
    5.977296267997333e-10, 5.9540843917576414e-10, 5.9315938524641762e-10, 
    5.9096246336949251e-10, 5.8879717318856194e-10, 5.8664371808923179e-10, 
    5.8448405575861737e-10, 5.8230281299591992e-10, 5.8008795479754124e-10, 
    5.7783125050192104e-10, 5.7552844957995861e-10, 5.7317926150583525e-10, 
    5.7078707281214807e-10, 5.6835850936726326e-10, 5.6590280803137361e-10, 
    5.6343112491951743e-10, 5.6095575606546519e-10, 5.58489394414109e-10, 
    5.5604441401851122e-10, 5.5363228982357576e-10, 5.5126312771011477e-10, 
    5.4894538903637852e-10, 5.4668575268351772e-10, 5.4448917400508432e-10, 
    5.4235903068008825e-10, 5.4029740521154007e-10, 5.3830536376829923e-10, 
    5.363832763490388e-10, 5.3453102302004604e-10, 5.3274816568353485e-10, 
    5.3103395895185229e-10, 5.293872740576583e-10, 5.2780640351206542e-10, 
    5.2628881173784693e-10, 5.2483083371420795e-10, 5.2342743945077357e-10, 
    5.2207204025572105e-10, 5.2075646326753394e-10, 5.1947104396094924e-10, 
    5.1820493957217269e-10, 5.16946563743774e-10, 5.1568419985759271e-10, 
    5.1440666961946521e-10, 5.1310405643345074e-10, 5.1176836092755e-10, 
    5.1039406284691354e-10, 5.0897848867803668e-10, 5.0752198536387414e-10, 
    5.0602781356890893e-10, 5.0450183594172462e-10, 5.0295194645162307e-10, 
    5.0138735740585591e-10, 4.9981774650034901e-10, 4.9825239798169466e-10, 
    4.9669935429465355e-10, 4.9516471861048826e-10, 4.936521054344909e-10, 
    4.9216235104078533e-10, 4.9069342938881575e-10, 4.8924065753434045e-10, 
    4.8779708065436059e-10, 4.8635406866098455e-10, 4.8490199938780308e-10, 
    4.8343101937028037e-10, 4.8193176203276254e-10, 4.8039600591883957e-10, 
    4.7881718001024955e-10, 4.7719071712334292e-10, 4.7551419436828922e-10, 
    4.7378730145976786e-10, 4.720116015701317e-10, 4.7019016281078246e-10, 
    4.6832705061122957e-10, 4.6642677689456984e-10, 4.6449371037652827e-10, 
    4.6253155018140353e-10, 4.6054287062749002e-10, 4.5852882850435108e-10, 
    4.5648901638532285e-10, 4.5442154603256054e-10, 4.5232330842576363e-10, 
    4.5019045258732553e-10, 4.480189919409664e-10, 4.4580556195837771e-10, 
    4.4354816952698256e-10, 4.4124695260423362e-10, 4.3890478614440678e-10, 
    4.3652772126780155e-10, 4.3412513858386435e-10, 4.3170963344843399e-10, 
    4.2929656033693138e-10, 4.2690331221424205e-10, 4.2454834018056256e-10, 
    4.2225002742256667e-10, 4.2002549565278926e-10, 4.1788947950337777e-10, 
    4.1585334741994581e-10, 4.1392440152252436e-10, 4.1210548960332725e-10, 
    4.1039499357566327e-10, 4.0878716573540573e-10, 4.0727278619280306e-10, 
    4.0584004399650244e-10, 4.0447556535001721e-10, 4.0316544463483883e-10, 
    4.0189619025570667e-10, 4.0065547833243544e-10, 3.9943265445235016e-10, 
    3.9821894092001735e-10, 3.9700738151479122e-10, 3.957925204792323e-10, 
    3.9456995310103213e-10, 3.9333577116128277e-10, 3.9208605338545536e-10, 
    3.9081643808501506e-10, 3.8952189320926402e-10, 3.8819667643850238e-10, 
    3.8683453158092895e-10, 3.8542906817962334e-10, 3.8397430532860165e-10, 
    3.8246527062252661e-10, 3.8089863289493615e-10, 3.7927324289993991e-10, 
    3.7759055748422322e-10, 3.7585487572873868e-10, 3.7407337877651379e-10, 
    3.7225595627469937e-10, 3.7041485504141004e-10, 3.6856415612293136e-10, 
    3.6671915410557561e-10, 3.6489566540796142e-10, 3.6310933298735928e-10, 
    3.6137495426964373e-10, 3.5970589372330329e-10, 3.581135714968665e-10, 
    3.5660708799785398e-10, 3.5519294877097241e-10, 3.5387492866479709e-10, 
    3.5265402100930199e-10, 3.5152851756971461e-10, 3.5049415674908788e-10, 
    3.4954437026783792e-10, 3.486705838617981e-10, 3.47862589013377e-10, 
    3.4710895221446034e-10, 3.463974672308878e-10, 3.457156049349627e-10, 
    3.4505098512177283e-10, 3.4439178740693845e-10, 3.4372714352335751e-10, 
    3.4304743934150844e-10, 3.4234454514881451e-10, 3.416119562394026e-10, 
    3.4084484747667895e-10, 3.4004005251826231e-10, 3.3919599320457214e-10, 
    3.3831256715667321e-10, 3.3739102940146007e-10, 3.3643385547679559e-10, 
    3.3544463154442254e-10, 3.3442790928632211e-10, 3.3338907657070864e-10, 
    3.3233416907504627e-10, 3.312696441419503e-10, 3.3020206809883013e-10, 
    3.2913775972997729e-10, 3.2808234276001333e-10, 3.2704029726226501e-10, 
    3.2601451394646725e-10, 3.2500592540576015e-10, 3.2401325456397012e-10, 
    3.2303295097344629e-10, 3.2205932923754408e-10, 3.2108494656989957e-10, 
    3.2010116859331097e-10, 3.1909893167581566e-10, 3.1806958869604407e-10, 
    3.1700579511385418e-10, 3.1590232224201733e-10, 3.1475673031576748e-10, 
    3.135698121058266e-10, 3.1234578414959262e-10, 3.1109217076276424e-10, 
    3.0981941779555175e-10, 3.0854024321377761e-10, 3.0726879754880493e-10, 
    3.0601968892819293e-10, 3.0480697484944467e-10, 3.0364315747923953e-10, 
    3.0253831121035749e-10, 3.0149935562311781e-10, 3.0052955946097618e-10, 
    2.9962827212436957e-10, 2.9879093910832666e-10, 2.9800933332640773e-10, 
    2.972720488753814e-10, 2.9656515904238442e-10, 2.9587302333319613e-10, 
    2.9517916522287142e-10, 2.9446716787613186e-10, 2.9372151454828491e-10, 
    2.9292833839941595e-10, 2.9207600679875835e-10, 2.9115555393319918e-10, 
    2.9016091012037606e-10, 2.8908896965655538e-10, 2.879394794399233e-10, 
    2.8671482150530106e-10, 2.8541967987169633e-10, 2.8406067680695744e-10, 
    2.8264596614438589e-10, 2.8118484602172339e-10, 2.7968737628742725e-10, 
    2.7816404270752009e-10, 2.7662541537916083e-10, 2.7508186002984546e-10, 
    2.7354321834279662e-10, 2.7201853457992227e-10, 2.705157527828538e-10, 
    2.6904146504155274e-10, 2.6760066392854406e-10, 2.6619658653898329e-10, 
    2.6483063070097536e-10, 2.6350240922350168e-10, 2.6220992203686037e-10, 
    2.6094989823993955e-10, 2.5971825290769264e-10, 2.585106744453259e-10, 
    2.5732324363599398e-10, 2.5615307430498148e-10, 2.5499886222250913e-10, 
    2.5386130718285179e-10, 2.5274330097494476e-10, 2.516499023425004e-10, 
    2.5058801600309505e-10, 2.4956584138986715e-10, 2.4859209484568671e-10, 
    2.4767511825623259e-10, 2.4682191660352031e-10, 2.4603728504213582e-10, 
    2.4532306693273107e-10, 2.446776823901914e-10, 2.4409593923957258e-10, 
    2.4356920350234819e-10, 2.4308586814035363e-10, 2.4263212919095609e-10, 
    2.4219293588989048e-10, 2.4175308069548285e-10, 2.4129824488074126e-10, 
    2.408159786280924e-10, 2.4029644271608342e-10, 2.3973291656006999e-10, 
    2.3912198173366564e-10, 2.3846343113271818e-10, 2.3775987850245831e-10, 
    2.3701618523296124e-10, 2.3623873104151731e-10, 2.3543465283210286e-10, 
    2.3461108640821275e-10, 2.3377454433146419e-10, 2.3293040557617564e-10, 
    2.3208262782533022e-10, 2.3123361220322654e-10, 2.3038427197456383e-10, 
    2.2953420859724033e-10, 2.2868201598716932e-10, 2.2782560624390233e-10, 
    2.2696256618144246e-10, 2.2609044943907487e-10, 2.2520704801207872e-10, 
    2.2431055274582679e-10, 2.2339967693570324e-10, 2.2247369929264084e-10, 
    2.2153248196392935e-10, 2.2057644687240139e-10, 2.1960658216514101e-10, 
    2.1862442480782398e-10, 2.176321113574033e-10, 2.166323997731955e-10, 
    2.1562874799092346e-10, 2.1462534796965815e-10, 2.1362716676971319e-10, 
    2.126398951447474e-10, 2.1166987160064483e-10, 2.1072388595580256e-10, 
    2.0980893465952208e-10, 2.0893187758125391e-10, 2.0809908450184533e-10, 
    2.0731602850143683e-10, 2.0658695939779988e-10, 2.0591459328383477e-10, 
    2.0529995849539769e-10, 2.0474232230589146e-10, 2.0423929641692704e-10, 
    2.0378702768201713e-10, 2.033805322621737e-10, 2.0301403937301065e-10, 
    2.0268140503863489e-10, 2.0237644403499498e-10, 2.0209323573659088e-10, 
    2.0182629494918371e-10, 2.0157067683233486e-10, 2.0132194943339199e-10, 
    2.0107614072508376e-10, 2.0082960583804805e-10, 2.0057895165185768e-10, 
    2.0032095014379894e-10, 2.0005256294724936e-10, 1.9977100501940672e-10, 
    1.9947390215183402e-10, 1.9915946111350351e-10, 1.9882666818980506e-10, 
    1.9847542122549118e-10, 1.9810661178238502e-10, 1.9772206617974563e-10, 
    1.9732439423578371e-10, 1.9691667412174006e-10, 1.9650208824968962e-10, 
    1.960834644556566e-10, 1.956628584228742e-10, 1.9524116267688027e-10, 
    1.9481788814241597e-10, 1.9439106705535422e-10, 1.9395741045675172e-10, 
    1.9351262764755354e-10, 1.9305197638591194e-10, 1.9257090547033478e-10, 
    1.9206581187881696e-10, 1.9153475139278037e-10, 1.9097808377795642e-10, 
    1.9039890945814907e-10, 1.8980330467227259e-10, 1.8920023191819027e-10, 
    1.8860120678221351e-10, 1.8801963586125827e-10, 1.8746996650762e-10, 
    1.8696664165749787e-10, 1.8652300471133686e-10, 1.8615017539010562e-10, 
    1.858560796749515e-10, 1.8564461934325687e-10, 1.8551513932052767e-10, 
    1.8546215475973359e-10, 1.8547543971544242e-10, 1.8554039391723463e-10, 
    1.8563874074795652e-10, 1.8574943158500089e-10, 1.8584976745800074e-10, 
    1.8591657489001575e-10, 1.8592744520357589e-10, 1.8586188259148269e-10, 
    1.8570235968849565e-10, 1.8543513788561799e-10, 1.8505091607736019e-10, 
    1.8454518276010823e-10, 1.8391835933198091e-10, 1.8317566042915258e-10, 
    1.8232678019172747e-10, 1.8138535400666948e-10, 1.8036831583077165e-10, 
    1.792951043012603e-10, 1.7818683617552717e-10, 1.7706540292856003e-10, 
    1.7595260164321892e-10, 1.7486923809915962e-10, 1.7383433490326584e-10, 
    1.7286437696659172e-10, 1.7197270821238233e-10, 1.7116904066234485e-10, 
    1.704591690136353e-10, 1.6984483390557042e-10, 1.6932383147110103e-10, 
    1.6889027680061049e-10, 1.6853509819982111e-10, 1.6824663102493729e-10, 
    1.6801137649097746e-10, 1.6781478655464559e-10, 1.6764211075766096e-10, 
    1.6747915462871627e-10, 1.6731302039314744e-10, 1.6713270140373988e-10, 
    1.6692958091907418e-10, 1.666977411387814e-10, 1.6643417341467062e-10, 
    1.6613879719507176e-10, 1.6581437372057971e-10, 1.6546626301059098e-10, 
    1.6510209766134524e-10, 1.6473131750842598e-10, 1.6436466535839912e-10, 
    1.6401357887479868e-10, 1.6368958561293604e-10, 1.6340364036947346e-10, 
    1.6316552073868078e-10, 1.6298322868182835e-10, 1.628625017647182e-10, 
    1.6280639508962721e-10, 1.6281502388589582e-10, 1.6288542251773826e-10, 
    1.6301159246939028e-10, 1.6318467524244645e-10, 1.633933169627165e-10, 
    1.6362413574417217e-10, 1.6386234047293881e-10, 1.6409238578819065e-10, 
    1.6429871830584353e-10, 1.6446648951408307e-10, 1.6458227217752083e-10, 
    1.6463466046633311e-10, 1.6461480791926818e-10, 1.6451678248331419e-10, 
    1.6433780528585722e-10, 1.6407827864232091e-10, 1.6374167825788451e-10, 
    1.6333423259054932e-10, 1.6286449899933444e-10, 1.6234277215652773e-10, 
    1.6178044704956587e-10, 1.6118929486701133e-10, 1.6058078456690204e-10, 
    1.5996541856751458e-10, 1.5935220629889532e-10, 1.5874823163371975e-10, 
    1.5815843241191746e-10, 1.5758552550402745e-10, 1.5703015061438728e-10, 
    1.5649113774133656e-10, 1.5596595188216036e-10, 1.5545118852562223e-10, 
    1.5494313456280242e-10, 1.5443828496887833e-10, 1.5393382238567397e-10, 
    1.5342793412001159e-10, 1.5292003080782043e-10, 1.5241077768808667e-10, 
    1.5190200184383212e-10, 1.5139642531140177e-10, 1.508973504008525e-10, 
    1.5040824735980713e-10, 1.4993237974504417e-10, 1.4947242821052559e-10, 
    1.4903024651960296e-10, 1.4860667756700047e-10, 1.4820155126822005e-10, 
    1.4781375471602808e-10, 1.4744145498094499e-10, 1.4708237227981054e-10, 
    1.4673412133771832e-10, 1.4639451980028804e-10, 1.4606188599536484e-10, 
    1.4573523298681442e-10, 1.4541438691315141e-10, 1.4509996094813706e-10, 
    1.4479326137275311e-10, 1.4449605832737596e-10, 1.4421033414861273e-10, 
    1.4393798088573773e-10, 1.4368054483848628e-10, 1.434389703573029e-10, 
    1.4321347418434686e-10, 1.4300347113047057e-10, 1.4280764000632584e-10, 
    1.4262402349704502e-10, 1.4245025402164123e-10, 1.4228378506368772e-10, 
    1.4212216777476413e-10, 1.4196328002871015e-10, 1.4180555828876124e-10, 
    1.4164813323993661e-10, 1.4149093886817959e-10, 1.4133470360490358e-10, 
    1.4118090805430524e-10, 1.4103164190593249e-10, 1.4088942929966584e-10, 
    1.4075697716769414e-10, 1.4063692053949099e-10, 1.4053150294211705e-10, 
    1.4044229628839948e-10, 1.4036989649394668e-10, 1.4031368259180906e-10, 
    1.4027160354454054e-10, 1.4024006708638071e-10, 1.4021388476338376e-10, 
    1.4018636284130257e-10, 1.4014944504140446e-10, 1.4009400214796121e-10, 
    1.4001016921387014e-10, 1.3988777728164587e-10, 1.3971678025191541e-10, 
    1.3948771742096785e-10, 1.3919212108077862e-10, 1.3882288566843121e-10, 
    1.3837453706103146e-10, 1.3784343397239744e-10, 1.3722785490758452e-10, 
    1.3652801794462375e-10, 1.3574600394185674e-10, 1.348856440838588e-10, 
    1.3395234679086398e-10, 1.3295292692014862e-10, 1.318954024782156e-10, 
    1.3078882474257654e-10, 1.2964309445818451e-10, 1.2846881556109738e-10, 
    1.2727712701869178e-10, 1.2607957475731463e-10, 1.2488794162918621e-10, 
    1.2371409695720608e-10, 1.2256979906479842e-10, 1.2146650912647557e-10, 
    1.2041513321634341e-10, 1.1942578415145206e-10, 1.1850750227751365e-10, 
    1.1766799452947152e-10, 1.1691336087937645e-10, 1.1624788212382676e-10, 
    1.1567384297133298e-10, 1.1519144388986564e-10, 1.1479878759301346e-10, 
    1.1449198378431822e-10, 1.1426531550805016e-10, 1.1411151403842109e-10, 
    1.1402208449287452e-10, 1.1398766473384314e-10, 1.1399837408004602e-10, 
    1.1404415673003791e-10, 1.141150446725353e-10, 1.1420138578078005e-10, 
    1.142939858032215e-10, 1.1438422287215774e-10, 1.1446409724431806e-10, 
    1.1452630101039689e-10, 1.1456428393017128e-10, 1.145723567326953e-10, 
    1.1454581994178404e-10, 1.1448113937735586e-10, 1.1437610471290099e-10, 
    1.1422999705195274e-10, 1.1404368797453657e-10, 1.1381966999746654e-10, 
    1.135619798005732e-10, 1.1327601725801324e-10, 1.1296824038028697e-10, 
    1.1264579119120851e-10, 1.1231605348576698e-10, 1.1198621362992346e-10, 
    1.116628336968179e-10, 1.1135151833273504e-10, 1.1105667082481783e-10, 
    1.107813937202354e-10, 1.1052749272447791e-10, 1.1029561866686222e-10, 
    1.1008547382639908e-10, 1.0989609584944723e-10, 1.0972613175377596e-10, 
    1.0957409979164936e-10, 1.0943859951694305e-10, 1.0931845175552865e-10, 
    1.0921273682777271e-10, 1.0912078581666887e-10, 1.0904208264496692e-10, 
    1.0897615212846183e-10, 1.0892240155912438e-10, 1.0887999530305989e-10, 
    1.0884773529361498e-10, 1.0882399100552815e-10, 1.0880665974035919e-10, 
    1.0879317434945138e-10, 1.08780531175077e-10, 1.0876534447526769e-10, 
    1.0874390148772783e-10, 1.0871222472045376e-10, 1.0866611759742276e-10, 
    1.0860122617683496e-10, 1.085130983291722e-10, 1.0839727569460014e-10, 
    1.0824940941801111e-10, 1.0806543988527161e-10, 1.0784181631723197e-10, 
    1.075757665909889e-10, 1.0726560404122208e-10, 1.0691103839900607e-10, 
    1.0651345046915419e-10, 1.0607611972868819e-10, 1.0560432325425861e-10, 
    1.0510532551205161e-10, 1.0458820233486973e-10, 1.0406352060332466e-10, 
    1.0354286740738403e-10, 1.0303827943176567e-10, 1.0256160279915376e-10, 
    1.0212382962576535e-10, 1.0173448911800912e-10, 1.0140111692680841e-10, 
    1.0112884217137624e-10, 1.0092014355549042e-10, 1.0077476247151072e-10, 
    1.0068978817534732e-10, 1.0065987428041534e-10, 1.0067759947798381e-10, 
    1.0073392188235609e-10, 1.0081869904063416e-10, 1.0092125627853631e-10, 
    1.0103096985921264e-10, 1.0113784904111534e-10, 1.0123308773701021e-10, 
    1.0130956162396969e-10, 1.0136225039340851e-10, 1.0138854764295334e-10, 
    1.0138843539240533e-10, 1.013644779311828e-10, 1.013216345463949e-10, 
    1.0126686119296447e-10, 1.0120852407866281e-10, 1.0115563160333026e-10, 
    1.0111696284171694e-10, 1.0110014308286489e-10, 1.0111075493915724e-10, 
    1.0115158545984697e-10, 1.0122209045427505e-10, 1.0131814351004791e-10, 
    1.0143212799100405e-10, 1.0155337611927867e-10, 1.0166893631891372e-10, 
    1.0176460099091216e-10, 1.0182611475218964e-10, 1.0184043257113846e-10, 
    1.0179691950588055e-10, 1.0168836435748927e-10, 1.0151170639255734e-10, 
    1.0126840707366637e-10, 1.0096442530483822e-10, 1.0060981066485563e-10, 
    1.0021794444972593e-10, 9.9804519844241702e-11, 9.9386358376081824e-11, 
    9.8980156290869677e-11, 9.8601300594727081e-11, 9.8262836991615757e-11, 
    9.7974672215928695e-11, 9.7743055391458445e-11, 9.7570365958517148e-11, 
    9.7455209389829904e-11, 9.7392756074862276e-11, 9.737530241887168e-11, 
    9.7392970864055686e-11, 9.7434467206718219e-11, 9.7487860255570139e-11, 
    9.7541294830429743e-11, 9.7583610369224258e-11, 9.7604836543654846e-11, 
    9.7596554452688283e-11, 9.7552119273808457e-11, 9.7466770023468416e-11, 
    9.7337649218751044e-11, 9.7163742285319427e-11, 9.6945754181432209e-11, 
    9.6685956488142127e-11, 9.6387994598824591e-11, 9.6056654804462313e-11, 
    9.5697598030580026e-11, 9.5317041622595484e-11, 9.4921405982685834e-11, 
    9.4516914387205225e-11, 9.4109167368883807e-11, 9.3702724448747323e-11, 
    9.3300717697468441e-11, 9.2904533437687897e-11, 9.2513605601693716e-11, 
    9.2125342303670264e-11, 9.1735222696197499e-11, 9.1337051830549992e-11, 
    9.0923368573496571e-11, 9.0485985640329939e-11, 9.0016614424688666e-11, 
    8.9507532122060716e-11, 8.8952223426425317e-11, 8.8345959413561779e-11, 
    8.7686267825157103e-11, 8.697324734672505e-11, 8.6209721636591872e-11, 
    8.5401227761087965e-11, 8.4555828870563727e-11, 8.3683806277282408e-11, 
    8.2797230105590618e-11, 8.1909453473574089e-11, 8.1034576831755111e-11, 
    8.0186895699044475e-11, 7.9380363987337446e-11, 7.8628102149193895e-11, 
    7.7941951136244699e-11, 7.7332094150591578e-11, 7.6806719911558842e-11, 
    7.6371774403926943e-11, 7.6030751113977341e-11, 7.5784558075315599e-11, 
    7.5631458915595961e-11, 7.5567088283175062e-11, 7.5584540086117098e-11, 
    7.5674569669046559e-11, 7.5825865644986724e-11, 7.6025436406033142e-11, 
    7.6259064700842054e-11, 7.651183150273673e-11, 7.6768690819908729e-11, 
    7.7015050397452473e-11, 7.7237340930436637e-11, 7.7423541073057714e-11, 
    7.7563617286919475e-11, 7.7649877257712138e-11, 7.767718967092181e-11, 
    7.7643082125857105e-11, 7.7547706877866131e-11, 7.7393676593236868e-11, 
    7.7185773548829906e-11, 7.6930572678504365e-11, 7.6635973742917535e-11, 
    7.6310696492139488e-11, 7.5963746789696347e-11, 7.5603907455129833e-11, 
    7.5239270376273238e-11, 7.4876855621164164e-11, 7.4522321315464824e-11, 
    7.4179814203596373e-11, 7.385193316998137e-11, 7.3539831415981322e-11, 
    7.324343457810362e-11, 7.2961753071345514e-11, 7.2693250161854752e-11, 
    7.2436241875002398e-11, 7.2189292145843306e-11, 7.1951545388118495e-11, 
    7.1722989724203966e-11, 7.1504612618053985e-11, 7.1298441638733373e-11, 
    7.1107467573865473e-11, 7.0935456818472226e-11, 7.0786680460605654e-11, 
    7.0665575460756906e-11, 7.0576386051739758e-11, 7.0522806775907444e-11, 
    7.0507672988794913e-11, 7.0532710968307062e-11, 7.0598390769309294e-11, 
    7.0703863082092001e-11, 7.084700735089117e-11, 7.1024561253010012e-11, 
    7.1232326664496334e-11, 7.1465403952995458e-11, 7.1718465374056461e-11, 
    7.1985995846606662e-11, 7.2262514295050822e-11, 7.2542741814234436e-11, 
    7.2821708237146792e-11, 7.3094810913671122e-11, 7.3357820530398032e-11, 
    7.3606847317248103e-11, 7.3838309749483176e-11, 7.4048888050353208e-11, 
    7.4235513126031392e-11, 7.4395390259504831e-11, 7.452606288063521e-11, 
    7.4625520255910324e-11, 7.4692344689452351e-11, 7.4725870260198325e-11, 
    7.4726356493942915e-11, 7.4695120705469062e-11, 7.4634638604765091e-11, 
    7.4548560548949198e-11, 7.4441650570509544e-11, 7.4319633736356553e-11, 
    7.4188943310140483e-11, 7.4056403266584219e-11, 7.3928851920166918e-11, 
    7.3812740178618053e-11, 7.3713748987083661e-11, 7.3636445585751601e-11, 
    7.3584018789534226e-11, 7.3558098199698981e-11, 7.3558678734034184e-11, 
    7.3584145072131779e-11, 7.3631381108113809e-11, 7.3695929365420746e-11, 
    7.3772210951572515e-11, 7.3853746145837112e-11, 7.3933386436628618e-11, 
    7.4003536110414319e-11, 7.4056359809215386e-11, 7.4083996915072363e-11, 
    7.4078785595017052e-11, 7.4033505970103776e-11, 7.3941676445268225e-11, 
    7.3797871003949747e-11, 7.3598088251333004e-11, 7.3340122625382801e-11, 
    7.3023919433190911e-11, 7.2651885038105392e-11, 7.2229089747766947e-11, 
    7.1763328940112378e-11, 7.1265025382675549e-11, 7.0746931606013901e-11, 
    7.022365455943898e-11, 6.971099191490377e-11, 6.922516225116206e-11, 
    6.8781925670724324e-11, 6.839570317473875e-11, 6.8078749982794774e-11, 
    6.78404370220281e-11, 6.7686690328365245e-11, 6.7619658308917054e-11, 
    6.7637598574509772e-11, 6.7735005402229545e-11, 6.7902955960972035e-11, 
    6.8129651501660472e-11, 6.8401101188752405e-11, 6.8701912873704337e-11, 
    6.9016122679938232e-11, 6.9328020086926358e-11, 6.9622908267870266e-11, 
    6.9887773830583457e-11, 7.0111814364398203e-11, 7.0286811692819311e-11, 
    7.0407345833576856e-11, 7.0470844001623871e-11, 7.0477465115316062e-11, 
    7.0429878713740756e-11, 7.0332936892545645e-11, 7.0193290579024275e-11, 
    7.0018982287654903e-11, 6.9819049816900229e-11, 6.9603168762888417e-11, 
    6.9381347569299553e-11, 6.9163680928342813e-11, 6.896016285634261e-11, 
    6.8780526161952529e-11, 6.8634118590135773e-11, 6.8529758615167033e-11, 
    6.8475579133024142e-11, 6.8478841805003721e-11, 6.854570667758005e-11, 
    6.8680985982959811e-11, 6.8887882223143175e-11, 6.9167746352189474e-11, 
    6.9519873189006887e-11, 6.9941367121131683e-11, 7.042709881245928e-11, 
    7.0969745252986292e-11, 7.1559951709015446e-11, 7.2186587760497175e-11, 
    7.2837099698663554e-11, 7.3497929573866326e-11, 7.4155014355543989e-11, 
    7.479431172884e-11, 7.5402362239506927e-11, 7.5966846491727569e-11, 
    7.6477119850288215e-11, 7.6924691844404947e-11, 7.730362030967537e-11, 
    7.7610784846458694e-11, 7.7846012546727216e-11, 7.8012018812502964e-11, 
    7.8114163488620998e-11, 7.8160015377225541e-11, 7.8158746883757276e-11, 
    7.8120399861233016e-11, 7.8055078169679664e-11, 7.7972141301113626e-11, 
    7.7879476495384201e-11, 7.7782915910317897e-11, 7.7685875119997691e-11, 
    7.7589246589513067e-11, 7.7491567206071618e-11, 7.7389445509821552e-11, 
    7.7278202943104353e-11, 7.7152658275871904e-11, 7.7007968069618885e-11, 
    7.6840411743909091e-11, 7.6648039176532092e-11, 7.6431099157880069e-11, 
    7.6192181755618577e-11, 7.5936069544914532e-11, 7.5669298680732761e-11, 
    7.5399513251964193e-11, 7.5134654927245713e-11, 7.4882117214031657e-11, 
    7.4647968060337189e-11, 7.4436321268633075e-11, 7.4248949633851672e-11, 
    7.4085166032501982e-11, 7.3941976142740324e-11, 7.381448249403241e-11, 
    7.369645359242381e-11, 7.3580983507226749e-11, 7.3461150731790431e-11, 
    7.3330588319223962e-11, 7.3183901048049393e-11, 7.301690531353379e-11, 
    7.282667173447302e-11, 7.2611410982766508e-11, 7.2370246381812151e-11, 
    7.2102942491616231e-11, 7.1809653806383943e-11, 7.149072779791428e-11, 
    7.1146628314960857e-11, 7.0777974199261276e-11, 7.0385674703788761e-11, 
    6.9971144252476506e-11, 6.9536541186347597e-11, 6.9084979886758756e-11, 
    6.8620675648828065e-11, 6.8148974148576586e-11, 6.7676257601225149e-11, 
    6.720972240101344e-11, 6.6757047507239629e-11, 6.6325973184987558e-11, 
    6.5923848166886004e-11, 6.5557192089532193e-11, 6.5231306635925477e-11, 
    6.4949968428252096e-11, 6.4715250166755665e-11, 6.452747379981226e-11, 
    6.4385286799668511e-11, 6.4285849222571962e-11, 6.4225125534224069e-11, 
    6.4198221250910682e-11, 6.4199745816101934e-11, 6.4224169782504841e-11, 
    6.4266130245872965e-11, 6.4320665690572284e-11, 6.4383372643506847e-11, 
    6.4450466240363466e-11, 6.4518753896143149e-11, 6.4585533315220934e-11, 
    6.4648435129766659e-11, 6.4705232830687693e-11, 6.4753651013631294e-11, 
    6.4791196536683036e-11, 6.4815040411237425e-11, 6.4821961314355998e-11, 
    6.4808373939298888e-11, 6.4770445971689639e-11, 6.4704288450831813e-11, 
    6.4606219124548629e-11, 6.4473078285000638e-11, 6.4302551632666732e-11, 
    6.4093497768610762e-11, 6.3846223949976533e-11, 6.3562688392870827e-11, 
    6.3246603533718062e-11, 6.2903415969286181e-11, 6.2540156312958961e-11, 
    6.2165166688675789e-11, 6.1787708866615358e-11, 6.1417492331573803e-11, 
    6.1064158832115136e-11, 6.0736754726616364e-11, 6.0443248326615962e-11, 
    6.0190133444489709e-11, 5.9982147373582735e-11, 5.9822134461638602e-11, 
    5.9711061524025178e-11, 5.9648173645788532e-11, 5.9631285561671162e-11, 
    5.9657158666055049e-11, 5.9721932278443617e-11, 5.9821559517568753e-11, 
    5.9952213235702364e-11, 6.0110601513305344e-11, 6.0294188611560211e-11, 
    6.0501276995880296e-11, 6.0730955152071257e-11, 6.0982919348381375e-11, 
    6.1257185014217749e-11, 6.1553715090148317e-11, 6.1872012039494837e-11, 
    6.2210710270152361e-11, 6.2567224368992189e-11, 6.2937485373659203e-11, 
    6.3315800329096482e-11, 6.3694863781627735e-11, 6.4065931042026218e-11, 
    6.4419133718928732e-11, 6.4743924130064372e-11, 6.5029608861141095e-11, 
    6.5265929357212048e-11, 6.54436301603677e-11, 6.5554978755610891e-11, 
    6.5594187266190453e-11, 6.5557696478116461e-11, 6.5444321835227105e-11, 
    6.5255244620438112e-11, 6.499385835205743e-11, 6.4665499431393095e-11, 
    6.4277084260865798e-11, 6.3836699247029952e-11, 6.3353171724478948e-11, 
    6.2835658983051581e-11, 6.2293295134270239e-11, 6.1734909493910629e-11, 
    6.1168828667265794e-11, 6.0602777436318951e-11, 6.0043850693239682e-11, 
    5.9498556175858748e-11, 5.897288790110556e-11, 5.8472403511900777e-11, 
    5.8002274421515247e-11, 5.756727619474918e-11, 5.7171706751402161e-11, 
    5.6819225239667869e-11, 5.6512630238829719e-11, 5.6253592823208102e-11, 
    5.6042404895773937e-11, 5.5877769830757784e-11, 5.5756706603805899e-11, 
    5.5674591559525349e-11, 5.5625370086017318e-11, 5.5601941025850722e-11, 
    5.5596678730985436e-11, 5.5602070249533675e-11, 5.5611374733779411e-11, 
    5.5619250987708398e-11, 5.5622270376047243e-11,
  // Sqw-Na(9, 0-1999)
    0.018573651683116414, 0.018571529519307125, 0.018565225972342767, 
    0.018554925079295993, 0.018540917979938565, 0.01852358089764412, 
    0.0185033469246495, 0.018480673960643155, 0.018456011468086054, 
    0.018429768788430771, 0.018402287596522484, 0.018373820664056125, 
    0.018344518488991119, 0.018314424581573219, 0.01828347935427567, 
    0.01825153173108179, 0.018218356863664208, 0.01818367780356488, 
    0.018147188696917456, 0.018108577078703142, 0.018067543147379968, 
    0.018023814458942491, 0.017977155216630927, 0.017927370145620278, 
    0.017874303714420142, 0.017817836083166241, 0.017757877531392588, 
    0.017694363188717928, 0.017627249652501686, 0.017556514568016251, 
    0.017482159554618345, 0.017404216102541458, 0.0173227533681929, 
    0.017237886280474766, 0.017149782125732805, 0.0170586638478239, 
    0.016964808672643432, 0.016868541282345374, 0.016770221522618558, 
    0.016670227404411889, 0.016568934837217074, 0.016466696003359503, 
    0.016363818487993401, 0.016260547199917364, 0.01615705078194719, 
    0.016053413681790508, 0.015949634423513898, 0.015845629980075954, 
    0.015741245583105613, 0.01563626887868667, 0.015530447079838286, 
    0.015423505680612478, 0.015315167361556026, 0.015205169893592076, 
    0.015093282092099477, 0.014979317141650685, 0.014863142868970846, 
    0.014744688762976764, 0.014623949714035141, 0.014500986568364758, 
    0.01437592367458207, 0.014248943650068924, 0.014120279630194077, 
    0.013990205298809847, 0.013859023047087827, 0.013727050678407673, 
    0.013594607171738635, 0.013461998128503024, 0.013329501643137938, 
    0.013197355432564065, 0.013065746106946219, 0.012934801436210919, 
    0.012804586342870615, 0.012675103123304434, 0.012546296075219092, 
    0.012418060315680214, 0.012290254155706603, 0.012162714008895334, 
    0.012035270510300199, 0.01190776435771455, 0.011780060393458407, 
    0.011652058629568446, 0.01152370126470858, 0.011394975203704352, 
    0.011265910108019733, 0.011136572506455196, 0.011007056911173371, 
    0.010877475160022141, 0.010747945309744409, 0.010618581331086164, 
    0.010489484628348944, 0.010360738067425268, 0.010232402806693252, 
    0.010104517846697608, 0.0099771019023780286, 0.0098501569945862229, 
    0.009723673072810456, 0.0095976330123745384, 0.0094720174508321365, 
    0.0093468091004471811, 0.009221996352674169, 0.0090975761373334255, 
    0.0089735560871219127, 0.0088499560778328816, 0.0087268091748362586, 
    0.0086041619406171301, 0.0084820739787774321, 0.0083606165399307993, 
    0.0082398700202039998, 0.0081199202561320263, 0.0080008536566503075, 
    0.0078827513938109547, 0.0077656830669629532, 0.0076497004231275423, 
    0.0075348318238341334, 0.0074210781693730965, 0.007308410912874732, 
    0.0071967726226562822, 0.0070860803011088347, 0.0069762313731591549, 
    0.0068671119548443004, 0.0067586067413839095, 0.0066506096482638064, 
    0.0065430342233523666, 0.0064358228366745377, 0.0063289537487225683, 
    0.0062224453480724641, 0.0061163571147219873, 0.0060107871795055008, 
    0.0059058666798670507, 0.0058017514239558513, 0.0056986116354963848, 
    0.0055966207327508522, 0.0054959441754985836, 0.0053967293842343885, 
    0.0052990975981855254, 0.0052031383087394831, 0.005108906609763644, 
    0.0050164234821300909, 0.0049256787167163175, 0.0048366359169796326, 
    0.004749238840630496, 0.0046634182600132747, 0.004579098548062239, 
    0.0044962033215537704, 0.0044146596729835686, 0.0043344007645421869, 
    0.0042553668059782711, 0.0041775046577169472, 0.0041007664630827575, 
    0.0040251078007913828, 0.003950485855172498, 0.003876858033157498, 
    0.0038041813304877867, 0.0037324125884835363, 0.0036615096137255615, 
    0.0035914329817636533, 0.0035221482334521653, 0.0034536281124293556, 
    0.0033858544896563539, 0.0033188196721723397, 0.003252526887175635, 
    0.0031869898527321365, 0.0031222314737903833, 0.0030582818179925972, 
    0.0029951756142051682, 0.0029329495668797886, 0.0028716397865361787, 
    0.0028112796023822546, 0.0027518979545608203, 0.0026935184721985097, 
    0.0026361592432201254, 0.0025798331870689837, 0.0025245488648330716, 
    0.002470311512517353, 0.0024171240678589447, 0.0023649879799977382, 
    0.002313903640733085, 0.0022638703482792677, 0.0022148857987579771, 
    0.0021669451850325917, 0.0021200400549094664, 0.0020741571308869654, 
    0.0020292773142510309, 0.0019853750841505083, 0.0019424184585985717, 
    0.0019003696147731456, 0.0018591861798256588, 0.001818823112348561, 
    0.0017792350112038793, 0.0017403786241393156, 0.001702215292519213, 
    0.001664713065736804, 0.0016278482500549142, 0.0015916062177074792, 
    0.00155598138501185, 0.0015209763620506471, 0.0014866003689547581, 
    0.0014528670931663475, 0.0014197922185815001, 0.0013873908848283476, 
    0.0013556753309357328, 0.0013246529443577066, 0.0012943248795881383, 
    0.0012646853390140761, 0.0012357215321748989, 0.001207414258041224, 
    0.0011797389966247056, 0.0011526673569390495, 0.0011261687106899759, 
    0.0011002118445281397, 0.001074766484972316, 0.0010498045839891516, 
    0.001025301293587421, 0.0010012355986499613, 0.00097759061357868783, 
    0.00095435357672085674, 0.00093151559533892752, 0.000909071203135418, 
    0.00088701779344130109, 0.00086535498631665295, 0.00084408397944652402, 
    0.00082320692304920407, 0.00080272634968611689, 0.00078264468177612696, 
    0.0007629638329822283, 0.00074368491412563336, 0.00072480804928067976, 
    0.00070633230257458133, 0.00068825571052796722, 0.00067057540843892414, 
    0.00065328783265567077, 0.00063638897427315097, 0.00061987465473738017, 
    0.00060374079100753342, 0.00058798361813062225, 0.00057259984081249843, 
    0.00055758669284116031, 0.00054294189350844173, 0.00052866350244116188, 
    0.00051474968703538388, 0.00050119842831807546, 0.00048800719989567406, 
    0.00047517265934599208, 0.00046269039114838048, 0.00045055473489928654, 
    0.00043875872272971931, 0.00042729413680044195, 0.00041615168324472552, 
    0.00040532126491585801, 0.00039479232363577311, 0.00038455421481860925, 
    0.00037459657425148435, 0.00036490963865711917, 0.00035548448795626257, 
    0.000346313186854132, 0.00033738881509077427, 0.00032870538789542096, 
    0.00032025767943775395, 0.00031204097122381424, 0.00030405075367019097, 
    0.00029628241215951358, 0.00028873092876771877, 0.00028139062790914906, 
    0.00027425498892830099, 0.00026731654185864609, 0.00026056685488234352, 
    0.00025399661415337251, 0.0002475957892137217, 0.00024135387076977479, 
    0.00023526016251624457, 0.00022930410527949722, 0.00022347561013292075, 
    0.00021776537730054966, 0.00021216517945508856, 0.00020666809116892462, 
    0.0002012686504515131, 0.00019596294314311695, 0.00019074860608603276, 
    0.00018562475016352484, 0.00018059180923761235, 0.00017565132553003842, 
    0.00017080568588992784, 0.00016605782648556179, 0.000161410925529271, 
    0.00015686810446769681, 0.00015243215743753575, 0.00014810532657491795, 
    0.00014388913698576764, 0.00013978430003854154, 0.00013579068753755242, 
    0.00013190737287161258, 0.00012813272912235419, 0.00012446456909665345, 
    0.00012090030895549687, 0.00011743713598299612, 0.0001140721622195113, 
    0.00011080254899985052, 0.00010762559241325724, 0.00010453876562926048, 
    0.00010153972007778546, 9.8626252805244716e-05, 9.5796251247843903e-05, 
    9.3047628700063654e-05, 9.0378263730763174e-05, 8.7785954844341575e-05, 
    8.5268398204677021e-05, 8.2823191845835567e-05, 8.0447865193906343e-05, 
    7.8139928619710633e-05, 7.5896934714604321e-05, 7.3716541419720889e-05, 
    7.1596567183921178e-05, 6.9535029871851592e-05, 6.753016386310261e-05, 
    6.558041319875751e-05, 6.368440219027049e-05, 6.1840888076751939e-05, 
    6.0048702662475919e-05, 5.8306691106044118e-05, 5.6613656064732171e-05, 
    5.4968314305407865e-05, 5.3369270909233987e-05, 5.181501366162247e-05, 
    5.0303927514642364e-05, 4.8834326510714144e-05, 4.7404498572870437e-05, 
    4.6012757312524857e-05, 4.465749457536403e-05, 4.3337227821356393e-05, 
    4.2050637491535443e-05, 4.0796591055929345e-05, 3.9574152221186432e-05, 
    3.8382575557049685e-05, 3.7221288354230455e-05, 3.6089862684781283e-05, 
    3.4987981298475382e-05, 3.3915401133430579e-05, 3.2871917893119162e-05, 
    3.1857334453120882e-05, 3.0871434950433759e-05, 2.9913965433038492e-05, 
    2.8984621049277115e-05, 2.8083039049520049e-05, 2.7208796423041724e-05, 
    2.6361410821998179e-05, 2.5540343504390164e-05, 2.4745003299256292e-05, 
    2.3974750975916745e-05, 2.3228903798618294e-05, 2.2506740387778065e-05, 
    2.1807506232144941e-05, 2.1130420269716539e-05, 2.0474682878474329e-05, 
    1.9839485414206664e-05, 1.9224021148709067e-05, 1.8627497153322937e-05, 
    1.8049146401358772e-05, 1.7488239179179865e-05, 1.6944092838221024e-05, 
    1.6416079003518994e-05, 1.5903627572597967e-05, 1.5406227161467094e-05, 
    1.4923422036952653e-05, 1.4454805959512629e-05, 1.4000013693174675e-05, 
    1.3558711170071816e-05, 1.3130585396559753e-05, 1.2715335144050498e-05, 
    1.2312663293766036e-05, 1.1922271429726035e-05, 1.1543856943965542e-05, 
    1.1177112579740738e-05, 1.0821728040071984e-05, 1.0477393065125705e-05, 
    1.0143801256039234e-05, 9.8206538992221374e-06, 9.5076631169227976e-06, 
    9.2045538157966707e-06, 8.9110641010568937e-06, 8.6269440404336843e-06, 
    8.3519528758795684e-06, 8.0858549694727413e-06, 7.8284149195421687e-06, 
    7.5793923825429798e-06, 7.3385371820585949e-06, 7.1055852759013179e-06, 
    6.8802560893143681e-06, 6.6622516106297133e-06, 6.451257495397682e-06, 
    6.2469462463950398e-06, 6.0489823463195509e-06, 5.857029032938683e-06, 
    5.6707562423497427e-06, 5.4898491201112745e-06, 5.3140164273748424e-06, 
    5.1429981571266574e-06, 4.9765717277620708e-06, 4.8145562317083777e-06, 
    4.6568143757346437e-06, 4.503251939560973e-06, 4.3538147821038718e-06, 
    4.2084836187184424e-06, 4.0672669609681608e-06, 3.9301927367302762e-06, 
    3.7972991850068245e-06, 3.6686256423377577e-06, 3.5442038101783338e-06, 
    3.42405002186322e-06, 3.3081589260068371e-06, 3.1964988818829381e-06, 
    3.0890092348245542e-06, 2.9855995150071586e-06, 2.8861504896725927e-06, 
    2.7905169003655071e-06, 2.6985316360515039e-06, 2.610011029607379e-06, 
    2.5247609199361012e-06, 2.4425830942626433e-06, 2.363281716885933e-06, 
    2.2866693623128958e-06, 2.2125723047958757e-06, 2.1408347719630815e-06, 
    2.0713219469098e-06, 2.0039215952650621e-06, 1.938544295293383e-06, 
    1.8751223498096738e-06, 1.8136075495709706e-06, 1.753968028540361e-06, 
    1.6961844963247518e-06, 1.6402461477906356e-06, 1.5861465367287912e-06, 
    1.5338796632857365e-06, 1.4834364729875113e-06, 1.4348019067067439e-06, 
    1.3879525857956328e-06, 1.3428551702751444e-06, 1.2994653949924493e-06, 
    1.2577277674338421e-06, 1.217575899407445e-06, 1.1789334367896761e-06, 
    1.1417155426151482e-06, 1.1058308739882915e-06, 1.0711839719968153e-06, 
    1.0376779564385895e-06, 1.0052173887600349e-06, 9.7371114192173804e-07, 
    9.430751019593922e-07, 9.1323452667315644e-07, 8.8412590552512833e-07, 
    8.5569819994547061e-07, 8.279133921168586e-07, 8.0074632606384027e-07, 
    7.7418388147719572e-07, 7.4822357015584998e-07, 7.2287168306764297e-07, 
    6.98141138369048e-07, 6.7404918803523831e-07, 6.5061513347711281e-07, 
    6.2785818330431161e-07, 6.0579556202281195e-07, 5.8444095193927321e-07, 
    5.6380332363513918e-07, 5.4388618563296661e-07, 5.2468726077522275e-07, 
    5.0619857587448935e-07, 4.8840693060681684e-07, 4.7129469231829154e-07, 
    4.5484084449462913e-07, 4.3902220076722864e-07, 4.2381468411909916e-07, 
    4.091945659936117e-07, 3.9513956290954787e-07, 3.8162970106411958e-07, 
    3.6864788084689339e-07, 3.5618010239165131e-07, 3.4421534618887808e-07, 
    3.3274513641739163e-07, 3.217628441028598e-07, 3.1126280982069109e-07, 
    3.0123937806359331e-07, 2.9168593764943331e-07, 2.8259405420650164e-07, 
    2.7395276482920519e-07, 2.6574808330182181e-07, 2.5796274110074023e-07, 
    2.5057616680479414e-07, 2.4356468787968702e-07, 2.3690192470852678e-07, 
    2.3055933855072449e-07, 2.2450689143173401e-07, 2.1871377681715464e-07, 
    2.1314918284000405e-07, 2.0778305453513065e-07, 2.0258682585854186e-07, 
    1.9753409655254649e-07, 1.926012318569753e-07, 1.8776786580595866e-07, 
    1.830172906880838e-07, 1.7833671764439037e-07, 1.7371739582011114e-07, 
    1.6915458131395975e-07, 1.6464735149410826e-07, 1.6019826631798615e-07, 
    1.558128848143172e-07, 1.5149915277593495e-07, 1.4726668549638244e-07, 
    1.4312597759346736e-07, 1.3908757889308963e-07, 1.3516128127287298e-07, 
    1.3135536434474985e-07, 1.2767594819253809e-07, 1.241264973490926e-07, 
    1.207075125482074e-07, 1.1741643466034001e-07, 1.1424777021758932e-07, 
    1.1119343044929549e-07, 1.082432582652965e-07, 1.053857012259198e-07, 
    1.0260857608693409e-07, 9.9899862590339285e-08, 9.7248462933443417e-08, 
    9.464486791643964e-08, 9.208168158540747e-08, 8.9553970896384243e-08, 
    8.7059424458694627e-08, 8.4598321601577596e-08, 8.2173328732937824e-08, 
    7.9789151508784441e-08, 7.7452078857938009e-08, 7.5169457238948861e-08, 
    7.2949132297169521e-08, 7.0798890675546371e-08, 6.8725929439268146e-08, 
    6.6736374961081662e-08, 6.4834869010397368e-08, 6.3024236733698991e-08, 
    6.130524986228704e-08, 5.9676497131588303e-08, 5.8134372505271017e-08, 
    5.667318834264116e-08, 5.5285415436933758e-08, 5.3962043829481883e-08, 
    5.2693049002801826e-08, 5.1467937500676044e-08, 5.027633690161188e-08, 
    4.9108587813614457e-08, 4.7956292719735671e-08, 4.6812777709054247e-08, 
    4.5673429706154589e-08, 4.4535882081717713e-08, 4.3400035229102401e-08, 
    4.2267913224235509e-08, 4.1143372192371664e-08, 4.0031687991958035e-08, 
    3.8939059881915813e-08, 3.7872071506318877e-08, 3.6837151586205879e-08, 
    3.5840073527293318e-08, 3.4885527616075945e-08, 3.3976791330040581e-08, 
    3.3115514661225385e-08, 3.2301627833800351e-08, 3.1533370266566914e-08, 
    3.0807431364216241e-08, 3.0119187287115658e-08, 2.9463012260434138e-08, 
    2.8832639613638695e-08, 2.8221545672543839e-08, 2.7623329953085645e-08, 
    2.7032066767797602e-08, 2.6442607236570463e-08, 2.5850815449840784e-08, 
    2.5253728702321036e-08, 2.4649637692290473e-08, 2.4038088788427169e-08, 
    2.3419815368963758e-08, 2.2796609340512549e-08, 2.2171146116947381e-08, 
    2.1546777564003296e-08, 2.0927306800649262e-08, 2.0316757824765786e-08, 
    1.9719150936636732e-08, 1.9138293398173327e-08, 1.8577592924595729e-08, 
    1.8039900592759721e-08, 1.7527388555266447e-08, 1.7041467381066107e-08, 
    1.6582746584069364e-08, 1.6151040737078604e-08, 1.5745421260550225e-08, 
    1.536431152481292e-08, 1.5005619466139234e-08, 1.4666898849574e-08, 
    1.4345527105676912e-08, 1.4038885884604646e-08, 1.3744529497691806e-08, 
    1.3460327557448924e-08, 1.3184570452316471e-08, 1.2916030437544096e-08, 
    1.2653975675490239e-08, 1.239813983699082e-08, 1.214865412427083e-08, 
    1.1905952240809932e-08, 1.1670660475646635e-08, 1.1443485471145738e-08, 
    1.1225110635611341e-08, 1.1016109768056177e-08, 1.0816882907382628e-08, 
    1.0627616299498926e-08, 1.0448265058022614e-08, 1.0278555166389012e-08, 
    1.011799996473709e-08, 9.9659263090868266e-09, 9.8215058759526898e-09, 
    9.6837884359742383e-09, 9.5517349827878157e-09, 9.4242500448944411e-09, 
    9.3002131595846458e-09, 9.1785101716197939e-09, 9.0580648071092616e-09, 
    8.9378708112736501e-09, 8.8170240880207256e-09, 8.694753814465318e-09, 
    8.5704506120209291e-09, 8.4436896218252379e-09, 8.3142459562034648e-09, 
    8.1821003932115312e-09, 8.0474334605106607e-09, 7.9106071558625865e-09, 
    7.7721343443581955e-09, 7.6326373551331212e-09, 7.492798234637647e-09, 
    7.3533044172447115e-09, 7.2147940772053939e-09, 7.0778060087027308e-09, 
    6.9427385049351034e-09, 6.809821286320999e-09, 6.6791031568837685e-09, 
    6.5504569080204813e-09, 6.4236010410895421e-09, 6.2981365312478032e-09, 
    6.1735951612602165e-09, 6.0494950997473376e-09, 5.9253985809089666e-09, 
    5.8009666794412765e-09, 5.6760064115067335e-09, 5.5505064648853784e-09, 
    5.4246588271238514e-09, 5.2988651325369774e-09, 5.1737276468898536e-09, 
    5.050026165437272e-09, 4.9286828279747839e-09, 4.8107176781298916e-09, 
    4.6971978814267364e-09, 4.5891837737839387e-09, 4.4876745625946841e-09, 
    4.3935564686256726e-09, 4.3075555532902062e-09, 4.2301974288504878e-09, 
    4.1617755395204156e-09, 4.1023296866861733e-09, 4.0516359575161752e-09, 
    4.0092090981489412e-09, 3.9743176736304599e-09, 3.9460120133939557e-09, 
    3.9231639537720949e-09, 3.9045168509585583e-09, 3.8887432621008816e-09, 
    3.8745071874362639e-09, 3.8605269820018994e-09, 3.8456349964880257e-09, 
    3.8288298404715273e-09, 3.8093177848122997e-09, 3.7865403964786658e-09, 
    3.7601867786182582e-09, 3.7301897812175848e-09, 3.6967071155524134e-09, 
    3.6600892369624859e-09, 3.6208371497932764e-09, 3.5795537385923022e-09, 
    3.5368927601230589e-09, 3.4935093643937157e-09, 3.4500158175785024e-09, 
    3.4069451474437871e-09, 3.3647247280546425e-09, 3.3236606596435862e-09, 
    3.2839329882291541e-09, 3.2456007821312215e-09, 3.2086156150873962e-09, 
    3.1728413500944884e-09, 3.1380781145177384e-09, 3.1040881338589364e-09, 
    3.0706214692496513e-09, 3.037439793191491e-09, 3.0043368814250528e-09, 
    2.9711547035122195e-09, 2.9377945955310929e-09, 2.9042231388496139e-09, 
    2.8704729229761951e-09, 2.8366384453963984e-09, 2.8028678525239419e-09, 
    2.7693512235664428e-09, 2.7363064631659118e-09, 2.7039637444123244e-09, 
    2.6725497204241235e-09, 2.6422724743539758e-09, 2.61330830188809e-09, 
    2.5857910905867607e-09, 2.5598050286874295e-09, 2.5353809818180402e-09, 
    2.5124967715331954e-09, 2.4910811406366228e-09, 2.47102111878723e-09, 
    2.4521720516697117e-09, 2.4343695526928e-09, 2.4174423228749393e-09, 
    2.4012248453456925e-09, 2.3855688310082505e-09, 2.3703525466331071e-09, 
    2.3554871651774271e-09, 2.3409197110777882e-09, 2.3266323175864394e-09, 
    2.3126380489850384e-09, 2.2989736733584161e-09, 2.2856902662521782e-09, 
    2.2728425239187713e-09, 2.2604779814168021e-09, 2.2486271108458824e-09, 
    2.237295329666847e-09, 2.2264575645824235e-09, 2.216055896915962e-09, 
    2.2060003184847782e-09, 2.1961725290064665e-09, 2.1864322323201366e-09, 
    2.1766253978131127e-09, 2.1665936399411785e-09, 2.1561839980844155e-09, 
    2.1452582885879714e-09, 2.1337014129160024e-09, 2.1214280161929352e-09, 
    2.1083871900511707e-09, 2.0945649224359119e-09, 2.0799843279230791e-09, 
    2.0647036743780347e-09, 2.0488125102933132e-09, 2.0324261337193619e-09, 
    2.0156788767670367e-09, 1.9987165337341956e-09, 1.9816884727732128e-09, 
    1.9647397541048461e-09, 1.9480037421922495e-09, 1.9315954792792217e-09, 
    1.9156062183668165e-09, 1.9000992879263385e-09, 1.8851075815808992e-09, 
    1.8706327291465574e-09, 1.8566461024998566e-09, 1.8430915563780532e-09, 
    1.829889873505827e-09, 1.8169446141243734e-09, 1.8041491143965561e-09, 
    1.7913941370684924e-09, 1.7785757469365467e-09, 1.7656028058301411e-09, 
    1.7524036296084542e-09, 1.7389312538440176e-09, 1.7251670114843707e-09, 
    1.7111221133534461e-09, 1.6968372188872664e-09, 1.6823800013641599e-09, 
    1.6678410380307929e-09, 1.6533282949918511e-09, 1.6389607279206975e-09, 
    1.6248614216567816e-09, 1.6111507978378279e-09, 1.5979402705939092e-09, 
    1.5853267602312245e-09, 1.5733882511679357e-09, 1.5621806361374684e-09, 
    1.5517358282195178e-09, 1.542061205764092e-09, 1.5331402363311905e-09, 
    1.5249342285366503e-09, 1.5173849700653493e-09, 1.5104181526814417e-09, 
    1.5039472996190901e-09, 1.497878048556284e-09, 1.4921124917530022e-09, 
    1.486553426720764e-09, 1.481108229371056e-09, 1.4756922246694776e-09, 
    1.4702313382086421e-09, 1.4646639955391535e-09, 1.4589421577942046e-09, 
    1.4530315739399043e-09, 1.4469112401361002e-09, 1.4405722550572065e-09, 
    1.4340161297480308e-09, 1.4272527709406468e-09, 1.4202982274299609e-09, 
    1.4131724024090427e-09, 1.4058968127507531e-09, 1.3984925606408667e-09, 
    1.3909785781752259e-09, 1.3833702821114128e-09, 1.375678639798617e-09, 
    1.3679097650103029e-09, 1.3600649871819072e-09, 1.3521414378484969e-09, 
    1.3441330419923169e-09, 1.3360318749675761e-09, 1.3278297236915633e-09, 
    1.3195197559493668e-09, 1.3110981101644681e-09, 1.3025653216155638e-09, 
    1.293927398092431e-09, 1.2851965358473874e-09, 1.2763913230517218e-09, 
    1.2675365017549055e-09, 1.2586622031957928e-09, 1.2498027822360844e-09, 
    1.2409952555327761e-09, 1.2322775010074779e-09, 1.223686286836166e-09, 
    1.2152553364484722e-09, 1.2070135243101504e-09, 1.1989834158540575e-09, 
    1.1911802347626436e-09, 1.1836114202362845e-09, 1.1762767776825614e-09, 
    1.169169280164335e-09, 1.1622763877915577e-09, 1.1555818317575453e-09, 
    1.1490676107144954e-09, 1.1427160682794455e-09, 1.1365117729931893e-09, 
    1.1304430770771349e-09, 1.1245031573734842e-09, 1.1186905059955632e-09, 
    1.1130087859580862e-09, 1.1074661736991118e-09, 1.1020742084915072e-09, 
    1.096846347622439e-09, 1.091796309834968e-09, 1.0869364285724172e-09, 
    1.0822760796989778e-09, 1.0778203683910509e-09, 1.0735690715863395e-09, 
    1.0695159784247283e-09, 1.0656485680945555e-09, 1.0619480923644065e-09, 
    1.0583899690476144e-09, 1.0549445322218714e-09, 1.0515779976707485e-09, 
    1.0482536758996031e-09, 1.0449332923257955e-09, 1.041578415413693e-09, 
    1.0381518596119778e-09, 1.0346190632764296e-09, 1.0309493255684117e-09, 
    1.0271168956707953e-09, 1.0231018206748013e-09, 1.0188905790668121e-09, 
    1.01447641514655e-09, 1.0098594302993211e-09, 1.0050463616868561e-09, 
    1.0000501515800559e-09, 9.9488923004565142e-10, 9.8958664650125024e-10, 
    9.8416900936476547e-10, 9.7866534972653291e-10, 9.7310591000900959e-10, 
    9.675209681829716e-10, 9.6193968628343507e-10, 9.5638910247613287e-10, 
    9.508932383585773e-10, 9.4547239683818936e-10, 9.4014261350781269e-10, 
    9.3491531009866497e-10, 9.2979709348301199e-10, 9.2478973548359204e-10, 
    9.1989027295049884e-10, 9.1509127687801389e-10, 9.1038124660444127e-10, 
    9.057451854439055e-10, 9.0116530326860083e-10, 8.9662192530530062e-10, 
    8.9209452833546609e-10, 8.8756292917430729e-10, 8.8300851517921316e-10, 
    8.7841550850703951e-10, 8.7377209468623643e-10, 8.6907138121359062e-10, 
    8.6431203848520563e-10, 8.5949859771488135e-10, 8.5464128436252757e-10, 
    8.4975546773739576e-10, 8.4486069041706859e-10, 8.3997939148526235e-10, 
    8.351353913657481e-10, 8.3035230056406184e-10, 8.2565193720523753e-10, 
    8.2105291102758229e-10, 8.1656942667843779e-10, 8.1221044018964824e-10, 
    8.0797915696678082e-10, 8.0387294439896449e-10, 7.9988359842683859e-10, 
    7.959979953802996e-10, 7.9219902256228396e-10, 7.8846678348278647e-10, 
    7.8477993913875795e-10, 7.8111716136949682e-10, 7.7745854645859472e-10, 
    7.7378693027816558e-10, 7.7008897483583232e-10, 7.6635597393180852e-10, 
    7.6258426419438755e-10, 7.5877525792005685e-10, 7.5493503138135757e-10, 
    7.5107355859283758e-10, 7.4720361327132584e-10, 7.4333949167222051e-10, 
    7.39495610103168e-10, 7.3568520562200737e-10, 7.3191917124821763e-10, 
    7.2820522761798615e-10, 7.2454742668210626e-10, 7.2094610221392448e-10, 
    7.1739819446119776e-10, 7.1389796423956554e-10, 7.1043795468025144e-10, 
    7.0701014682734283e-10, 7.0360711747832233e-10, 7.0022313842251354e-10, 
    6.9685504369173173e-10, 6.9350282971525117e-10, 6.9016986892646726e-10, 
    6.8686278324237369e-10, 6.835909398656954e-10, 6.8036567882140937e-10, 
    6.7719929823928049e-10, 6.7410396804953984e-10, 6.7109061337463296e-10, 
    6.6816793593888451e-10, 6.6534160469888518e-10, 6.6261372837919865e-10, 
    6.5998261162429504e-10, 6.5744282843247614e-10, 6.549855428695151e-10, 
    6.525991077304427e-10, 6.5026977052494265e-10, 6.4798252284104159e-10, 
    6.4572193260442669e-10, 6.4347294726758448e-10, 6.4122157136748677e-10, 
    6.3895542240362536e-10, 6.366640944511182e-10, 6.3433938309032075e-10, 
    6.3197532866983381e-10, 6.2956815008828381e-10, 6.2711606756393725e-10, 
    6.2461907459580251e-10, 6.2207866064508064e-10, 6.1949754281546967e-10, 
    6.1687938597352499e-10, 6.1422855387832255e-10, 6.1154984687839643e-10, 
    6.0884825658002489e-10, 6.0612870551910296e-10, 6.0339578625334225e-10, 
    6.0065347503666505e-10, 5.9790487153971694e-10, 5.9515196519379831e-10, 
    5.9239547200727569e-10, 5.8963475510702367e-10, 5.8686790762988969e-10, 
    5.8409195024504533e-10, 5.8130322387137176e-10, 5.7849788610816953e-10, 
    5.7567253450223482e-10, 5.7282484857888498e-10, 5.6995421306440196e-10, 
    5.6706222287618761e-10, 5.641530195137342e-10, 5.6123338443800689e-10, 
    5.5831259640779625e-10, 5.5540200436373144e-10, 5.5251441378583566e-10, 
    5.4966328644981827e-10, 5.4686188577476686e-10, 5.4412240418227793e-10, 
    5.4145520841403759e-10, 5.3886822507492372e-10, 5.3636655527322297e-10, 
    5.3395230290455302e-10, 5.3162464785311683e-10, 5.2938010721793689e-10, 
    5.2721297344265465e-10, 5.2511584599870886e-10, 5.2308024134605483e-10, 
    5.210972047911021e-10, 5.1915791514208503e-10, 5.1725421708028139e-10, 
    5.1537911806545072e-10, 5.1352714864816344e-10, 5.116946651269223e-10, 
    5.0987999861176036e-10, 5.0808348954161197e-10, 5.0630736822611774e-10, 
    5.0455548457772948e-10, 5.0283287556434686e-10, 5.011452138233557e-10, 
    4.9949813046314238e-10, 4.978965084473071e-10, 4.9634374954330957e-10, 
    4.9484114249311506e-10, 4.9338735315007404e-10, 4.9197812641362356e-10, 
    4.9060622447218583e-10, 4.8926163427562498e-10, 4.8793202306522291e-10, 
    4.8660341992705507e-10, 4.8526105350352675e-10, 4.8389028161930487e-10, 
    4.8247750434651917e-10, 4.8101101380940891e-10, 4.7948166853030641e-10, 
    4.7788336997243062e-10, 4.7621328657629596e-10, 4.744718531190798e-10, 
    4.7266252531917909e-10, 4.7079138696583562e-10, 4.6886661764363622e-10, 
    4.6689792243183785e-10, 4.6489595733276062e-10, 4.628718251411323e-10, 
    4.6083665077229914e-10, 4.5880128074894088e-10, 4.5677606820490601e-10, 
    4.5477076346485506e-10, 4.5279443382780603e-10, 4.5085542146568365e-10, 
    4.4896126643399847e-10, 4.4711859664664368e-10, 4.4533294970391779e-10, 
    4.4360855260784165e-10, 4.4194805258829416e-10, 4.4035225573697305e-10, 
    4.3881989110961638e-10, 4.3734746422448728e-10, 4.3592921755672142e-10, 
    4.3455724140101003e-10, 4.3322173429820162e-10, 4.3191141397947761e-10, 
    4.3061403631702219e-10, 4.2931700468060067e-10, 4.2800798556489805e-10, 
    4.2667550109284878e-10, 4.2530940975148187e-10, 4.2390128031824866e-10, 
    4.2244457876554995e-10, 4.2093471808551136e-10, 4.1936894715252617e-10, 
    4.1774614857404986e-10, 4.1606656409541233e-10, 4.143315324638503e-10, 
    4.1254325234167336e-10, 4.1070464503591329e-10, 4.0881929256305561e-10, 
    4.0689148013793036e-10, 4.0492628802024555e-10, 4.0292972024293588e-10, 
    4.0090878097460432e-10, 3.988715041524444e-10, 3.968268383475387e-10, 
    3.9478443121318299e-10, 3.9275426006019628e-10, 3.9074619130957167e-10, 
    3.8876946358099445e-10, 3.8683220560730887e-10, 3.8494100078500177e-10, 
    3.8310059516047791e-10, 3.8131374755389055e-10, 3.7958126991513367e-10, 
    3.7790220275460485e-10, 3.7627414044622565e-10, 3.746935842235415e-10, 
    3.7315633265589256e-10, 3.716577962848374e-10, 3.7019321869301835e-10, 
    3.687577687443095e-10, 3.673465216455507e-10, 3.6595434597342907e-10, 
    3.6457576764718657e-10, 3.6320485933358099e-10, 3.6183524997163959e-10, 
    3.6046026864051049e-10, 3.590733040193469e-10, 3.5766832947334617e-10, 
    3.5624059208746725e-10, 3.5478736892045883e-10, 3.5330871469923931e-10, 
    3.5180807026862802e-10, 3.5029265338096495e-10, 3.4877351172793222e-10, 
    3.4726521671202255e-10, 3.457851659119986e-10, 3.4435254001338383e-10, 
    3.4298698580499509e-10, 3.4170715763664151e-10, 3.4052922102674926e-10, 
    3.394655110629041e-10, 3.3852342006755581e-10, 3.3770467750138293e-10, 
    3.3700501805492569e-10, 3.364143331653818e-10, 3.3591721217111511e-10, 
    3.3549386214705722e-10, 3.3512126632543154e-10, 3.3477451137652357e-10, 
    3.344281347601271e-10, 3.3405742176815906e-10, 3.3363953866906e-10, 
    3.3315447863948237e-10, 3.3258575442982099e-10, 3.3192087315005047e-10, 
    3.3115157364027852e-10, 3.3027387536815796e-10, 3.2928795575881744e-10, 
    3.2819790207938525e-10, 3.270113406516635e-10, 3.25738988791091e-10, 
    3.2439412770233782e-10, 3.2299202315582927e-10, 3.2154928207625688e-10, 
    3.2008320970764498e-10, 3.1861112044575577e-10, 3.1714968956408037e-10, 
    3.157143198015603e-10, 3.1431857799288108e-10, 3.129736828403836e-10, 
    3.1168810702422549e-10, 3.1046723750386972e-10, 3.0931315845297529e-10, 
    3.0822452125256255e-10, 3.0719653355045609e-10, 3.0622105195375529e-10, 
    3.0528682601520203e-10, 3.0437987952884983e-10, 3.0348407097846368e-10, 
    3.0258181010532372e-10, 3.0165496308943626e-10, 3.0068587371678598e-10, 
    2.9965849387943181e-10, 2.9855951806815187e-10, 2.9737946651450138e-10, 
    2.9611358659960804e-10, 2.9476251273753603e-10, 2.933325739232893e-10, 
    2.9183573085314457e-10, 2.9028907441959446e-10, 2.8871396381893375e-10, 
    2.8713480087696732e-10, 2.8557760329239341e-10, 2.8406840607962581e-10, 
    2.8263171564247751e-10, 2.8128905813534244e-10, 2.8005779881852613e-10, 
    2.7895025736824384e-10, 2.7797323170305847e-10, 2.7712786980243869e-10, 
    2.7640994178920409e-10, 2.7581039496343748e-10, 2.7531615418387964e-10, 
    2.7491106528126278e-10, 2.745768926461591e-10, 2.7429428452002897e-10, 
    2.7404365869491298e-10, 2.7380591707522628e-10, 2.7356301847853123e-10, 
    2.7329834942694454e-10, 2.7299695381011668e-10, 2.7264559711961243e-10, 
    2.7223275843944663e-10, 2.7174853345523602e-10, 2.7118454560112329e-10, 
    2.7053384628764493e-10, 2.697908797981289e-10, 2.6895149292440855e-10, 
    2.6801302003961063e-10, 2.6697439389331128e-10, 2.6583632728702996e-10, 
    2.6460144482785417e-10, 2.632744299580135e-10, 2.6186206350056578e-10, 
    2.6037320347258687e-10, 2.5881862178058521e-10, 2.5721075234508497e-10, 
    2.5556331417932602e-10, 2.5389087776840658e-10, 2.5220834752269487e-10, 
    2.505304701649139e-10, 2.4887133505343643e-10, 2.4724395922409241e-10, 
    2.4565991728818086e-10, 2.4412909189781996e-10, 2.4265947483565695e-10, 
    2.4125708849453089e-10, 2.399259326004207e-10, 2.3866801941376095e-10, 
    2.3748343168236668e-10, 2.3637043678482638e-10, 2.353256201132741e-10, 
    2.3434408215051369e-10, 2.334196546097055e-10, 2.3254518345548934e-10, 
    2.3171282736300571e-10, 2.3091442026411088e-10, 2.3014180741842185e-10, 
    2.2938722647510133e-10, 2.286436208785471e-10, 2.2790495528348998e-10, 
    2.2716643941903082e-10, 2.2642471960954272e-10, 2.2567796065520715e-10, 
    2.2492588736257384e-10, 2.2416971414296678e-10, 2.2341202617243756e-10, 
    2.2265654880531064e-10, 2.2190787947341685e-10, 2.2117110468586088e-10, 
    2.2045139869479399e-10, 2.1975354615589957e-10, 2.19081488765606e-10, 
    2.1843785410234286e-10, 2.1782359826565412e-10, 2.1723770853941514e-10, 
    2.16677100009014e-10, 2.1613663798484117e-10, 2.1560938486029976e-10, 
    2.1508697034694051e-10, 2.1456014176568902e-10, 2.1401936174240177e-10, 
    2.1345546977036087e-10, 2.1286026018145447e-10, 2.1222701497435992e-10, 
    2.1155083267706579e-10, 2.1082883856643728e-10, 2.1006017835358575e-10, 
    2.0924589168899395e-10, 2.0838862699974381e-10, 2.0749232536674179e-10, 
    2.0656184003323773e-10, 2.0560263193076598e-10, 2.0462047397110171e-10, 
    2.0362128736075005e-10, 2.0261101829702636e-10, 2.015956239214153e-10, 
    2.0058106622648229e-10, 1.9957336302754615e-10, 1.9857858934541649e-10, 
    1.9760288533033132e-10, 1.9665238030529832e-10, 1.9573311004459817e-10, 
    1.9485085842457885e-10, 1.9401101479183145e-10, 1.9321838728266766e-10, 
    1.9247707109547876e-10, 1.9179029683403353e-10, 1.9116035208679954e-10, 
    1.9058848401583254e-10, 1.9007487129750054e-10, 1.8961855438132974e-10, 
    1.8921742314318283e-10, 1.888681537634031e-10, 1.8856620149154249e-10, 
    1.883057575805011e-10, 1.880797895985896e-10, 1.8788009418233438e-10, 
    1.8769745758816084e-10, 1.8752186878854774e-10, 1.8734286721253757e-10, 
    1.8714992534959294e-10, 1.869329450103043e-10, 1.8668274860010902e-10, 
    1.8639160349428931e-10, 1.8605366064615106e-10, 1.8566536130435172e-10, 
    1.8522566941519896e-10, 1.8473621892721826e-10, 1.8420126532560455e-10, 
    1.8362753279358127e-10, 1.8302386577518381e-10, 1.8240082442910237e-10, 
    1.8177013250387255e-10, 1.8114410263576648e-10, 1.8053498679689155e-10, 
    1.7995436274877292e-10, 1.7941248559823864e-10, 1.7891774816997637e-10, 
    1.7847615969215444e-10, 1.7809097855231006e-10, 1.7776243248329761e-10, 
    1.7748764210689176e-10, 1.772606847537353e-10, 1.7707289960506751e-10, 
    1.769133461515628e-10, 1.7676949571602897e-10, 1.7662803217302312e-10, 
    1.7647580462915047e-10, 1.7630076687613793e-10, 1.7609292347873041e-10, 
    1.7584511017351592e-10, 1.7555360778360251e-10, 1.7521843907997211e-10, 
    1.7484340201386701e-10, 1.7443572515773916e-10, 1.7400545710832396e-10, 
    1.7356454895489061e-10, 1.7312580099537924e-10, 1.7270167988374074e-10, 
    1.7230320067879566e-10, 1.7193890692831534e-10, 1.7161411877755624e-10, 
    1.7133042783911312e-10, 1.7108558470804762e-10, 1.708736923403297e-10, 
    1.7068576551731535e-10, 1.7051050424715533e-10, 1.7033530998399909e-10, 
    1.7014735065095889e-10, 1.6993465958177891e-10, 1.6968709605133275e-10, 
    1.6939716129115921e-10, 1.6906053067107741e-10, 1.6867633921611119e-10, 
    1.6824712648586867e-10, 1.6777853774949079e-10, 1.672787330358916e-10, 
    1.6675764983290331e-10, 1.6622609493227278e-10, 1.6569485505356862e-10, 
    1.6517380123831797e-10, 1.6467117093145717e-10, 1.6419299791149187e-10, 
    1.6374283241640388e-10, 1.6332168394247988e-10, 1.6292827034511738e-10, 
    1.625594696902267e-10, 1.6221099316802644e-10, 1.6187811181786776e-10, 
    1.6155645195196513e-10, 1.6124268007152145e-10, 1.6093507582997555e-10, 
    1.6063383418481882e-10, 1.6034116756962862e-10, 1.6006111012828028e-10, 
    1.5979911918701403e-10, 1.5956145483489215e-10, 1.5935449663440308e-10, 
    1.5918398913081686e-10, 1.5905438467952087e-10, 1.5896828127947486e-10, 
    1.5892607313967667e-10, 1.5892577277457149e-10, 1.5896308091040776e-10, 
    1.5903159872216623e-10, 1.5912322528485757e-10, 1.5922859333897028e-10, 
    1.593375869658666e-10, 1.5943978675199252e-10, 1.5952490109718603e-10, 
    1.595830700607724e-10, 1.5960511578225251e-10, 1.5958267352378939e-10, 
    1.595082981025763e-10, 1.5937549790510465e-10, 1.5917881118093036e-10, 
    1.5891386805530287e-10, 1.5857754530113374e-10, 1.5816812488026494e-10, 
    1.5768555115408839e-10, 1.5713167252442275e-10, 1.5651051384233256e-10, 
    1.5582846175302364e-10, 1.5509439441409793e-10, 1.5431962862305344e-10, 
    1.5351773144100441e-10, 1.5270410525005782e-10, 1.5189541471176854e-10, 
    1.5110880567898948e-10, 1.5036104429418202e-10, 1.4966756383545527e-10, 
    1.4904157334087571e-10, 1.4849323281419931e-10, 1.4802905827085198e-10, 
    1.4765152695855077e-10, 1.4735902814871565e-10, 1.4714605132891537e-10, 
    1.4700371448019486e-10, 1.4692048146417789e-10, 1.4688308490486247e-10, 
    1.4687748344044135e-10, 1.4688985040639495e-10, 1.4690742983141321e-10, 
    1.4691924343802267e-10, 1.4691655124349119e-10, 1.4689309243025784e-10, 
    1.4684502087481348e-10, 1.4677066221110185e-10, 1.4667005123404396e-10, 
    1.4654437691131619e-10, 1.463953337863823e-10, 1.462245381719484e-10, 
    1.4603298617137426e-10, 1.4582068630314736e-10, 1.4558642639985242e-10, 
    1.4532777189694533e-10, 1.4504120973772267e-10, 1.4472250281755438e-10, 
    1.4436713263025635e-10, 1.4397085792883087e-10, 1.4353027148185189e-10, 
    1.4304336470538924e-10, 1.425099635428252e-10, 1.4193209484912866e-10, 
    1.4131415673120473e-10, 1.4066295307925261e-10, 1.3998751922505723e-10, 
    1.3929881921660944e-10, 1.3860925312695953e-10, 1.3793208627235732e-10, 
    1.372807690948218e-10, 1.3666824719317806e-10, 1.3610623125256819e-10, 
    1.3560455495405705e-10, 1.3517059082051106e-10, 1.3480881648896741e-10, 
    1.3452050080938749e-10, 1.3430360973994834e-10, 1.3415287508830128e-10, 
    1.3406008829419045e-10, 1.3401454995417865e-10, 1.3400371725840884e-10, 
    1.3401395342330566e-10, 1.340313875107495e-10, 1.3404276960766495e-10, 
    1.3403632391294002e-10, 1.3400247341575106e-10, 1.3393443895620834e-10, 
    1.3382860017695289e-10, 1.3368465175249137e-10, 1.3350545647808007e-10, 
    1.3329668081959918e-10, 1.3306616393320612e-10, 1.3282312223945901e-10, 
    1.3257720774779926e-10, 1.3233753507372269e-10, 1.3211171824693592e-10, 
    1.3190505534645778e-10, 1.3171985934902973e-10, 1.3155507922219872e-10, 
    1.3140617798207178e-10, 1.3126534036297378e-10, 1.3112193087894206e-10, 
    1.3096323981376868e-10, 1.3077538691035342e-10, 1.305443576007309e-10, 
    1.3025703583565885e-10, 1.2990219132157726e-10, 1.2947128852317759e-10, 
    1.2895909643341235e-10, 1.2836400281240053e-10, 1.2768805549748428e-10, 
    1.2693668835602498e-10, 1.2611821681426714e-10, 1.2524309830848532e-10, 
    1.2432309214770485e-10, 1.2337035660260545e-10, 1.2239660697631448e-10, 
    1.2141238057260999e-10, 1.2042652110460626e-10, 1.1944586922334068e-10, 
    1.1847524150046014e-10, 1.1751762920212447e-10, 1.1657464164404701e-10, 
    1.156470633293507e-10, 1.1473553501733252e-10, 1.1384121542397223e-10, 
    1.1296638581306917e-10, 1.1211488939270261e-10, 1.1129240846333474e-10, 
    1.1050649283387763e-10, 1.0976637724922534e-10, 1.0908256835070687e-10, 
    1.0846627921619056e-10, 1.0792870553219081e-10, 1.0748027277855082e-10, 
    1.0712986931913312e-10, 1.0688415856706578e-10, 1.0674699286542199e-10, 
    1.0671901410398992e-10, 1.0679740881502057e-10, 1.0697587892807447e-10, 
    1.0724476561005383e-10, 1.0759135160989067e-10, 1.0800025168698659e-10, 
    1.0845391184044756e-10, 1.0893313232644648e-10, 1.0941762091715283e-10, 
    1.0988652504389876e-10, 1.1031897578440003e-10, 1.1069458966209081e-10, 
    1.1099401081446734e-10, 1.1119943072526723e-10, 1.1129516257336449e-10, 
    1.1126820978155551e-10, 1.1110887308997852e-10, 1.1081129942189184e-10, 
    1.1037399647916168e-10, 1.098002095339376e-10, 1.0909813521260261e-10, 
    1.0828088892829677e-10, 1.0736623376352072e-10, 1.0637600871038957e-10, 
    1.0533531130195564e-10, 1.0427142434251086e-10, 1.032126065049207e-10, 
    1.0218676813067779e-10, 1.0122018430229728e-10, 1.0033627980130943e-10, 
    9.9554618982240399e-11, 9.8890137246080147e-11, 9.8352680079342761e-11, 
    9.7946829385268385e-11, 9.7672063735392586e-11, 9.7523164317713359e-11, 
    9.7490866143982767e-11, 9.7562642511209907e-11, 9.7723608435821989e-11, 
    9.7957427667509174e-11, 9.8247209899175319e-11, 9.857629968997787e-11, 
    9.8928971017773018e-11, 9.9290954457974358e-11, 9.9649818048792423e-11, 
    9.9995174599877374e-11, 1.0031875110813497e-10, 1.0061428447324875e-10, 
    1.0087733779096358e-10, 1.0110499910688884e-10, 1.0129555034851466e-10, 
    1.0144809981514345e-10, 1.0156226730901736e-10, 1.0163790246925954e-10, 
    1.0167491980135333e-10, 1.0167322815149791e-10, 1.0163278620898335e-10, 
    1.0155374763263605e-10, 1.0143670539856831e-10, 1.0128294205825315e-10, 
    1.0109469720030904e-10, 1.0087534660782464e-10, 1.006294908042725e-10, 
    1.0036287987737727e-10, 1.0008219820818807e-10, 9.9794678945048355e-11, 
    9.9507601247886945e-11, 9.922770745357056e-11, 9.8960609332626497e-11, 
    9.8710214630150205e-11, 9.8478295788703864e-11, 9.8264200655779535e-11, 
    9.8064784045401208e-11, 9.7874537402986881e-11, 9.7685953543285555e-11, 
    9.7490077699349843e-11, 9.7277220350702824e-11, 9.703775742587788e-11, 
    9.6762993642971367e-11, 9.644599200872545e-11, 9.6082337427181702e-11, 
    9.5670751155424877e-11, 9.5213534958564951e-11, 9.4716777981710738e-11, 
    9.4190324953542151e-11, 9.3647462535173568e-11, 9.3104356784323649e-11, 
    9.2579229255835324e-11, 9.2091345646565813e-11, 9.1659829579721837e-11, 
    9.1302423148664164e-11, 9.1034238967568554e-11, 9.0866626519373972e-11, 
    9.0806226902098451e-11, 9.0854320165729811e-11, 9.1006502521582782e-11, 
    9.1252775644222647e-11, 9.1578022651678003e-11, 9.1962879890681665e-11, 
    9.2384911969690797e-11, 9.2820050435006761e-11, 9.3244124316356009e-11, 
    9.3634423243348515e-11, 9.39711106798882e-11, 9.4238411439921749e-11, 
    9.4425460464219479e-11, 9.4526764771124355e-11, 9.4542241250830267e-11, 
    9.4476867676933957e-11, 9.4339972906163272e-11, 9.4144278566211293e-11, 
    9.3904744731221489e-11, 9.3637377136108076e-11, 9.3358058297954985e-11, 
    9.3081514054513424e-11, 9.2820453024909399e-11, 9.2584952379641942e-11, 
    9.2382082654906338e-11, 9.2215769348685476e-11, 9.2086860649333161e-11, 
    9.1993383776553106e-11, 9.1930902157414374e-11, 9.1892989452484835e-11, 
    9.1871723975875783e-11, 9.1858210029524086e-11, 9.1843074326993343e-11, 
    9.1816944366921066e-11, 9.1770852957959015e-11, 9.1696616319397753e-11, 
    9.1587138889145571e-11, 9.1436675290622111e-11, 9.1241008200096851e-11, 
    9.0997601179112818e-11, 9.0705677572547105e-11, 9.0366260660405575e-11, 
    8.9982149010956836e-11, 8.9557847961681618e-11, 8.9099430922700653e-11, 
    8.8614352248758526e-11, 8.811116560472622e-11, 8.7599195400522553e-11, 
    8.7088117863538831e-11, 8.6587492831124488e-11, 8.6106236538887256e-11, 
    8.5652081099124377e-11, 8.5231043898548813e-11, 8.4846959010526434e-11, 
    8.4501080960935481e-11, 8.4191850852687596e-11, 8.3914809052087862e-11, 
    8.3662715297886165e-11, 8.3425844198126024e-11, 8.3192484807742681e-11, 
    8.294957828091485e-11, 8.2683484674394512e-11, 8.2380783568965092e-11, 
    8.2029102201922373e-11, 8.1617850147810504e-11, 8.1138872952195002e-11, 
    8.058693400601689e-11, 7.9960030856417226e-11, 7.9259533886397892e-11, 
    7.8490152164127706e-11, 7.7659730129115816e-11, 7.6778944056974976e-11, 
    7.5860884544750446e-11, 7.492058616619426e-11, 7.3974497656768167e-11, 
    7.3039946150879329e-11, 7.2134561089629146e-11, 7.127569682655102e-11, 
    7.0479845858628203e-11, 6.9762042094667425e-11, 6.9135257317716521e-11, 
    6.8609844152419812e-11, 6.8193006035563612e-11, 6.7888373825086316e-11, 
    6.7695701004231665e-11, 6.7610732842641583e-11, 6.7625273381314877e-11, 
    6.7727485090616948e-11, 6.7902398712895899e-11, 6.8132652651354075e-11, 
    6.8399377440742587e-11, 6.8683217546519166e-11, 6.8965365292107526e-11, 
    6.9228579336116147e-11, 6.9458078101089924e-11, 6.9642262177516713e-11, 
    6.9773200395734896e-11, 6.984687689460823e-11, 6.9863169466094735e-11, 
    6.9825600859736347e-11, 6.974087534769466e-11, 6.9618273426392961e-11, 
    6.9468925983943811e-11, 6.9305045485295808e-11, 6.9139135755405677e-11, 
    6.8983242872272646e-11, 6.8848239614527183e-11, 6.8743202529362841e-11, 
    6.8674871394944926e-11, 6.8647227687742207e-11, 6.8661187553528695e-11, 
    6.8714456643257896e-11, 6.880154737035066e-11, 6.8913994379088993e-11, 
    6.9040753412010175e-11, 6.9168823992015909e-11, 6.9284032418298935e-11, 
    6.9371980250180125e-11, 6.9419059600416697e-11, 6.9413496459813118e-11, 
    6.9346312631021027e-11, 6.9212132182457098e-11, 6.9009743542613411e-11, 
    6.8742372920551467e-11, 6.8417614351670694e-11, 6.8047041819267032e-11, 
    6.7645504215077476e-11, 6.7230188907885654e-11, 6.6819517757083887e-11, 
    6.6431985183847236e-11, 6.6085009698083461e-11, 6.5793922599878271e-11, 
    6.5571115823089574e-11, 6.5425445250738e-11, 6.5361866770066233e-11, 
    6.5381329139376039e-11, 6.5480897451558462e-11, 6.5654067139149527e-11, 
    6.5891216636656395e-11, 6.6180185046348036e-11, 6.6506895422826213e-11, 
    6.6856026003094168e-11, 6.7211679547514479e-11, 6.755804630912177e-11, 
    6.7880028733367144e-11, 6.8163843742099712e-11, 6.8397550329360584e-11, 
    6.8571531337269803e-11, 6.8678865536779665e-11, 6.8715620007790181e-11, 
    6.8680989405679201e-11, 6.8577311593540905e-11, 6.8409923829470494e-11, 
    6.818686497570522e-11, 6.7918427528289974e-11, 6.761659546438098e-11, 
    6.729437536467301e-11, 6.6965092714452994e-11, 6.6641673395636007e-11, 
    6.6335981361574437e-11, 6.6058238653401126e-11, 6.5816583393515341e-11, 
    6.5616783257333174e-11, 6.5462130808408939e-11, 6.5353486307577232e-11, 
    6.5289497819735782e-11, 6.5266930835073747e-11, 6.5281090429366556e-11, 
    6.5326283861065306e-11, 6.5396280171855742e-11, 6.5484732603279462e-11, 
    6.5585535986277098e-11, 6.5693091737397332e-11, 6.5802499935454157e-11, 
    6.5909661627575339e-11, 6.6011340381957199e-11, 6.6105187276191986e-11, 
    6.6189763097369942e-11, 6.6264586481758994e-11, 6.6330205659658367e-11, 
    6.6388285808862816e-11, 6.6441713321297829e-11, 6.6494665580092929e-11, 
    6.6552622240307064e-11, 6.6622265615583761e-11, 6.6711253251147971e-11, 
    6.6827826842598382e-11, 6.6980275333892457e-11, 6.717627062616528e-11, 
    6.7422129364997471e-11, 6.772204369587308e-11, 6.8077402720215198e-11, 
    6.8486247389643453e-11, 6.8942951266746839e-11, 6.9438170211435906e-11, 
    6.9959097890795854e-11, 7.0490011267571919e-11, 7.1013075343169093e-11, 
    7.1509337013768427e-11, 7.1959829028706735e-11, 7.2346664295448624e-11, 
    7.2654054208105294e-11, 7.2869143718157748e-11, 7.298260268505199e-11, 
    7.298895597030029e-11, 7.2886638802141717e-11, 7.2677785306312111e-11, 
    7.2367840550092321e-11, 7.1965030547000062e-11, 7.1479769283257697e-11, 
    7.0924076937768043e-11, 7.0311049460138156e-11, 6.9654428973102391e-11, 
    6.8968280208281465e-11, 6.8266765217435708e-11, 6.7564001006741625e-11, 
    6.6873944719310354e-11, 6.6210291375926269e-11, 6.5586317006895174e-11, 
    6.5014664414547698e-11, 6.4507046634783061e-11, 6.4073868106900365e-11, 
    6.3723793222034133e-11, 6.3463294589842767e-11, 6.3296226047787203e-11, 
    6.3223479765171394e-11, 6.3242764394440479e-11, 6.3348570146473687e-11, 
    6.3532314268302084e-11, 6.3782710749413459e-11, 6.408634091905479e-11, 
    6.4428388240946808e-11, 6.4793483323838719e-11, 6.5166617384468287e-11, 
    6.5534017176294359e-11, 6.5883928221763286e-11, 6.6207237378885127e-11, 
    6.64978617439816e-11, 6.675289106536863e-11, 6.6972461740485462e-11, 
    6.7159379090319115e-11, 6.7318538714772457e-11, 6.7456181660793017e-11, 
    6.7579084535809591e-11, 6.76937439960969e-11, 6.7805632715218235e-11, 
    6.7918600988124514e-11, 6.8034458352247081e-11, 6.8152782028690303e-11, 
    6.8270946681751989e-11, 6.8384367087851448e-11, 6.8486928495422287e-11, 
    6.8571552437475644e-11, 6.8630847439774674e-11, 6.8657783983686912e-11, 
    6.8646334100846313e-11, 6.8592023676928092e-11, 6.8492358773524655e-11, 
    6.8347073580735706e-11, 6.8158216306608948e-11, 6.7930045026712517e-11, 
    6.766876355957056e-11, 6.738211752193899e-11, 6.7078893259098795e-11, 
    6.6768376304965167e-11, 6.6459795737857489e-11, 6.6161817316256535e-11, 
    6.5882118576111668e-11, 6.5627066904204191e-11, 6.5401527008051619e-11, 
    6.5208791110215038e-11, 6.5050619885751617e-11, 6.4927390790674271e-11, 
    6.4838307576267036e-11, 6.4781656936059961e-11, 6.475507742050202e-11, 
    6.4755824972044273e-11, 6.4780998410288979e-11, 6.4827739416833349e-11, 
    6.4893369788345098e-11, 6.4975485674079475e-11, 6.5072000647051945e-11, 
    6.518115323734539e-11, 6.5301480345573479e-11, 6.5431760738204098e-11, 
    6.5570949425897498e-11, 6.5718105701429235e-11, 6.5872312197460851e-11, 
    6.6032610071131172e-11, 6.6197929728376242e-11, 6.6367042238762761e-11, 
    6.6538524282801702e-11, 6.6710739259866106e-11, 6.6881833138293713e-11, 
    6.7049768783510891e-11, 6.7212370367276223e-11, 6.7367395836023753e-11, 
    6.7512625132759197e-11, 6.7645973212659853e-11, 6.7765599253392552e-11, 
    6.7869994206828683e-11, 6.7958050739385836e-11, 6.8029092018879224e-11, 
    6.8082834112218999e-11, 6.8119286747695362e-11, 6.813859916017556e-11, 
    6.8140849596366398e-11, 6.8125810177296057e-11, 6.8092718644193074e-11, 
    6.8040083180518321e-11, 6.7965555513155308e-11, 6.7865902768623702e-11, 
    6.773710035204769e-11, 6.7574532502236536e-11, 6.7373304265623854e-11, 
    6.7128632498328708e-11, 6.6836277534276476e-11, 6.6492975495893704e-11, 
    6.6096822680165981e-11, 6.5647578506162323e-11, 6.5146848173718726e-11, 
    6.4598135039666055e-11, 6.4006763017751664e-11, 6.3379656834514138e-11, 
    6.2725029921052848e-11, 6.2051979312066287e-11, 6.1370039285466447e-11, 
    6.068871097436222e-11, 6.001701739695226e-11, 5.9363093480116641e-11, 
    5.8733855042401817e-11, 5.8134750969841053e-11, 5.7569632938343692e-11, 
    5.7040730114254444e-11, 5.6548752428729538e-11, 5.6093094325341844e-11, 
    5.5672148210103326e-11, 5.5283674353514159e-11, 5.4925216376647156e-11, 
    5.4594510027598999e-11, 5.4289854916323166e-11, 5.4010398593008922e-11, 
    5.3756313099935245e-11, 5.3528832086520254e-11, 5.333015186277112e-11, 
    5.3163194269159779e-11, 5.30312594720963e-11, 5.2937588467660522e-11, 
    5.288491052178186e-11, 5.2874972398981122e-11, 5.2908142396103219e-11, 
    5.2983096485677893e-11, 5.3096640844395768e-11, 5.32436756015086e-11, 
    5.341732608298934e-11, 5.3609216128879227e-11, 5.3809888645969373e-11, 
    5.4009318056696248e-11, 5.4197502827582697e-11, 5.4365075872789635e-11, 
    5.4503883287764411e-11, 5.4607493653467921e-11, 5.4671595983794595e-11, 
    5.4694239159261832e-11, 5.4675913564025726e-11, 5.4619444262055552e-11, 
    5.4529728123038808e-11, 5.4413316242536313e-11, 5.4277898115309463e-11, 
    5.4131711404244649e-11, 5.3982946577285374e-11, 5.3839177259509979e-11, 
    5.3706885291664853e-11, 5.3591079531000796e-11, 5.3495071266447019e-11, 
    5.3420382788349022e-11, 5.3366807634995929e-11, 5.3332583238511788e-11, 
    5.3314675529385962e-11, 5.3309115448332539e-11, 5.3311383892447294e-11, 
    5.331678465046273e-11, 5.33207999658054e-11, 5.3319392288688671e-11, 
    5.3309254132584952e-11, 5.3287976284631982e-11, 5.3254149361161047e-11, 
    5.3207388740689129e-11, 5.3148294483951869e-11, 5.3078335935553352e-11, 
    5.2999703020666223e-11, 5.2915091806290761e-11, 5.2827486897116067e-11, 
    5.2739919676190633e-11, 5.2655251148940468e-11, 5.2575979271501763e-11, 
    5.2504107801715753e-11, 5.2441074517218635e-11, 5.2387750131052951e-11, 
    5.2344503707706185e-11, 5.2311324111834069e-11, 5.2287969741104468e-11, 
    5.2274126665974234e-11, 5.2269543970698877e-11 ;

 Sqw-total =
  // Sqw-total(0, 0-1999)
    0.16264009699303753, 0.16163195674087402, 0.15864770764826069, 
    0.15380514226206929, 0.14729176699180579, 0.1393524593616951, 
    0.13027383547503818, 0.12036673358617973, 0.10994831686305906, 
    0.099325230216068719, 0.088779031953772916, 0.078554798247496838, 
    0.068853415111728225, 0.059827679980985565, 0.051581979507114198, 
    0.044175027791425736, 0.037624961515112652, 0.031916001741108611, 
    0.027005899224711735, 0.022833463190995908, 0.019325608911908092, 
    0.016403521530830373, 0.013987698987304252, 0.012001786890437873, 
    0.010375240235901299, 0.0090449347750758517, 0.0079559040427553355, 
    0.0070614001892050447, 0.0063224741406666899, 0.0057072506321317711, 
    0.0051900435683674487, 0.0047504232022174469, 0.0043723135084038555, 
    0.0040431689958580347, 0.0037532566795906012, 0.0034950514692314799, 
    0.0032627414297212894, 0.0030518323367845165, 0.0028588375838190083, 
    0.0026810387004511946, 0.002516302557979268, 0.0023629430095332788, 
    0.0022196167065938674, 0.0020852448078428963, 0.0019589540663330412, 
    0.0018400322726997479, 0.0017278942408673875, 0.0016220554797017899, 
    0.0015221114432420429, 0.0014277208361235822, 0.0013385919043727606, 
    0.0012544709905647779, 0.0011751328943861812, 0.0011003727679236609, 
    0.0010299993999876931, 0.00096382981529464715, 0.00090168514247112317, 
    0.00084338770023365201, 0.00078875922457802099, 0.00073762012192970378, 
    0.00068978959355591428, 0.00064508644322357179, 0.00060333035919526415, 
    0.00056434345695785743, 0.00052795188181945407, 0.00049398729947444024, 
    0.00046228814439681307, 0.00043270054539455439, 0.0004050788988143719, 
    0.00037928610665530839, 0.00035519353397137185, 0.00033268076375126738, 
    0.00031163523634836378, 0.00029195185512092783, 0.00027353262285206669, 
    0.00025628634884715059, 0.00024012843917202014, 0.00022498075703376627, 
    0.00021077152073033218, 0.00019743519547503466, 0.0001849123336900722, 
    0.00017314932544746538, 0.00016209803468846264, 0.00015171531490792761, 
    0.00014196241702854842, 0.00013280431926115537, 0.00012420902144364513, 
    0.00011614685309345094, 0.00010858984453757229, 0.00010151120426698478, 
    9.4884934141277144e-05, 8.8685598896624549e-05, 8.2888249582038017e-05, 
    7.746848418600925e-05, 7.2402614791630123e-05, 6.7667900743733359e-05, 
    6.3242802611001073e-05, 5.9107212617027603e-05, 5.5242623418463625e-05, 
    5.1632207690004791e-05, 4.8260794444064084e-05, 4.5114742545829798e-05, 
    4.2181725557956254e-05, 3.9450453127144967e-05, 3.6910361278759551e-05, 
    3.4551306494398493e-05, 3.2363296256155487e-05, 3.0336282465943761e-05, 
    2.8460034922837715e-05, 2.6724101345693431e-05, 2.5117849820743087e-05, 
    2.3630580454418935e-05, 2.2251686480606814e-05, 2.0970841705251976e-05, 
    1.9778191037523368e-05, 1.8664523562482037e-05, 1.7621412399844295e-05, 
    1.6641311521025419e-05, 1.5717605788553881e-05, 1.4844615899683309e-05, 
    1.4017564056517627e-05, 1.323250875086998e-05, 1.2486258032469446e-05, 
    1.1776270268796764e-05, 1.1100550096201904e-05, 1.0457545470862679e-05, 
    9.8460498786437113e-06, 9.2651121855560806e-06, 8.7139554864092156e-06, 
    8.1919056794496663e-06, 7.6983302669762918e-06, 7.232587895388389e-06, 
    6.7939892039644211e-06, 6.3817694885318663e-06, 5.9950733941937184e-06, 
    5.6329513146889761e-06, 5.2943664503859435e-06, 4.9782106895230769e-06, 
    4.6833267769536306e-06, 4.4085337715930874e-06, 4.1526526697021795e-06, 
    3.914529332846438e-06, 3.6930524733018869e-06, 3.4871653244232817e-06, 
    3.2958706151716795e-06, 3.1182294226927322e-06, 2.9533552481522464e-06, 
    2.8004051475483776e-06, 2.658569901438571e-06, 2.5270650410171868e-06, 
    2.4051241257678254e-06, 2.2919950955272868e-06, 2.1869399064744302e-06, 
    2.0892371162584257e-06, 1.9981866800487537e-06, 1.913116001606738e-06, 
    1.8333862486778917e-06, 1.7583980640223055e-06, 1.6875960287684708e-06, 
    1.6204715102440592e-06, 1.556563797802156e-06, 1.495459662571493e-06, 
    1.4367916454693882e-06, 1.3802354788153902e-06, 1.3255070816312443e-06, 
    1.2723595494199702e-06, 1.2205804959676965e-06, 1.169990009208814e-06, 
    1.1204393638710945e-06, 1.0718105014236026e-06, 1.0240161520648717e-06, 
    9.7700034960047608e-07, 9.307389909083374e-07, 8.852400359835092e-07, 
    8.4054293992036911e-07, 7.9671696490327747e-07, 7.538581301980822e-07, 
    7.120847124120026e-07, 6.7153138243369025e-07, 6.323422370902922e-07, 
    5.9466312474833546e-07, 5.5863375694660409e-07, 5.2438012853578543e-07, 
    4.9200773860070912e-07, 4.6159601964913039e-07, 4.3319426337242989e-07, 
    4.0681919558458935e-07, 3.8245422404722088e-07, 3.600502736625068e-07, 
    3.395280465000076e-07, 3.2078149700832794e-07, 3.0368229362981334e-07, 
    2.880850344162121e-07, 2.7383298767840642e-07, 2.6076412811954081e-07, 
    2.4871723202360531e-07, 2.3753777975405704e-07, 2.270833984563622e-07, 
    2.1722856835381526e-07, 2.0786832467366728e-07, 1.9892071998837551e-07, 
    1.9032787473557853e-07, 1.8205553330628256e-07, 1.7409115525487507e-07, 
    1.6644069104551518e-07, 1.5912430760131204e-07, 1.521714225283964e-07, 
    1.4561546715182782e-07, 1.3948881512332721e-07, 1.3381828542757102e-07, 
    1.2862155674261015e-07, 1.2390472530431626e-07, 1.1966111254990362e-07, 
    1.1587129963790379e-07, 1.1250424726477131e-07, 1.0951926714131329e-07, 
    1.0686855362755485e-07, 1.0449996654438956e-07, 1.0235977641773066e-07, 
    1.0039513619378529e-07, 9.8556117024003802e-08, 9.6797228609874412e-08, 
    9.507842226860117e-08, 9.336563813975157e-08, 9.1630996817749689e-08, 
    8.98527494971814e-08, 8.8015089385171374e-08, 8.6107898147843559e-08, 
    8.4126462207470493e-08, 8.207115642557085e-08, 7.9947063607756924e-08, 
    7.776348603563139e-08, 7.5533309912604098e-08, 7.3272204462592309e-08, 
    7.0997668445102167e-08, 6.8727970771953789e-08, 6.6481059857086977e-08, 
    6.427353324829148e-08, 6.2119758872742262e-08, 6.0031224204723994e-08, 
    5.8016160051446114e-08, 5.6079449834860776e-08, 5.4222797814281585e-08, 
    5.244509946237497e-08, 5.0742937734564743e-08, 4.9111124469619162e-08, 
    4.7543214975989895e-08, 4.6031944769243791e-08, 4.4569564104166545e-08, 
    4.314807426970975e-08, 4.1759392688198761e-08, 4.0395489139031617e-08, 
    3.904853878140664e-08, 3.7711131321618554e-08, 3.6376558745495753e-08, 
    3.5039183244026178e-08, 3.3694863305320859e-08, 3.2341396633279325e-08, 
    3.0978924576591942e-08, 2.9610238443436159e-08, 2.8240932443426995e-08, 
    2.6879361481171155e-08, 2.5536381349989782e-08, 2.4224872679464028e-08, 
    2.2959072741963391e-08, 2.1753760972366831e-08, 2.0623359218331514e-08, 
    1.9581017164809077e-08, 1.8637755206426554e-08, 1.7801731811922856e-08, 
    1.707769102572362e-08, 1.646662985234329e-08, 1.5965706314867019e-08, 
    1.5568389269712875e-08, 1.5264831862721146e-08, 1.504243423554221e-08, 
    1.4886547903772161e-08, 1.4781266288449447e-08, 1.4710242505367403e-08, 
    1.4657477585548713e-08, 1.4608028432608391e-08, 1.4548595141979929e-08, 
    1.4467959602713101e-08, 1.4357261267630455e-08, 1.4210108988011595e-08, 
    1.402254042645044e-08, 1.3792849573420946e-08, 1.3521310167752502e-08, 
    1.320982580452866e-08, 1.2861538740525176e-08, 1.2480426856455067e-08, 
    1.2070915482961523e-08, 1.1637525417995581e-08, 1.1184574518892066e-08, 
    1.0715944805818799e-08, 1.0234923657620377e-08, 9.7441232786787785e-09, 
    9.2454797547083461e-09, 8.7403287950687791e-09, 8.229551837206216e-09, 
    7.7137809733656414e-09, 7.1936468618066257e-09, 6.6700480325892063e-09, 
    6.14441664969951e-09, 5.618952436517326e-09, 5.0967970276758353e-09, 
    4.5821235550461233e-09, 4.0801228968857852e-09, 3.596876798916761e-09, 
    3.1391198349743586e-09, 2.7139036112065493e-09, 2.3281882389767958e-09, 
    1.9883945677197839e-09, 1.6999563861564507e-09, 1.4669123575637678e-09, 
    1.2915747098148083e-09, 1.1743040144234853e-09, 1.1134098678947398e-09, 
    1.1051852962104049e-09, 1.1440715018887631e-09, 1.2229384747157831e-09, 
    1.3334590036755268e-09, 1.4665473096171075e-09, 1.6128308564169154e-09, 
    1.7631232755882783e-09, 1.9088688013257988e-09, 2.0425322106948761e-09, 
    2.1579139095847618e-09, 2.2503754026443765e-09, 2.3169674792252354e-09, 
    2.3564589382032291e-09, 2.3692702396068182e-09, 2.3573208588279558e-09, 
    2.3238039034133746e-09, 2.2729041848242413e-09, 2.2094782350989174e-09, 
    2.1387155412086807e-09, 2.0658005833882428e-09, 1.9955938646877963e-09, 
    1.9323490752665879e-09, 1.8794805155672512e-09, 1.8393924762127332e-09, 
    1.8133781976211355e-09, 1.8015923527532859e-09, 1.803096338037675e-09, 
    1.815971396157338e-09, 1.8374899817420694e-09, 1.8643322386140754e-09, 
    1.8928310821695225e-09, 1.9192278651538685e-09, 1.939919860267953e-09, 
    1.9516821311788802e-09, 1.9518486648661582e-09, 1.9384417971550859e-09, 
    1.9102434926255869e-09, 1.8668074920096538e-09, 1.8084163590861711e-09, 
    1.7359922180894193e-09, 1.6509732295964594e-09, 1.5551702231342478e-09, 
    1.450618235232203e-09, 1.3394367044561273e-09, 1.2237098164890494e-09, 
    1.1053949767140613e-09, 9.8626347590683328e-10, 8.6787343349132908e-10, 
    7.5157133354798119e-10, 6.3851580088536469e-10, 5.2971507629912281e-10, 
    4.2606947975777507e-10, 3.2841011860193508e-10, 2.3752703416896936e-10, 
    1.5418188093576412e-10, 7.9103185979373793e-11, 1.2964612990191535e-11, 
    -4.3650426505494667e-11, -9.0293076172168685e-11, 
    -1.2669572537007282e-10, -1.5281464749026821e-10, 
    -1.6886225101689176e-10, -1.7532399090744604e-10, 
    -1.7295651922854481e-10, -1.6276598592075208e-10, 
    -1.4596740008209094e-10, -1.2392817718409306e-10, 
    -9.8100591144142323e-11, -6.9949106352393548e-11, 
    -4.0878756932196805e-11, -1.217069074035476e-11, 1.5070247724699991e-11, 
    3.9952305203130479e-11, 6.1816648240906107e-11, 8.0240423872788344e-11, 
    9.5025322826005158e-11, 1.0617495893983413e-10, 1.1386527019142008e-10, 
    1.1841191358004192e-10, 1.2023827198298552e-10, 1.1984649919820634e-10, 
    1.1779272869010747e-10, 1.146663104740917e-10, 1.1107211768016702e-10, 
    1.0761400156988608e-10, 1.0487795415341464e-10, 1.0341330235677738e-10, 
    1.0371167027000671e-10, 1.0618385184868827e-10, 1.1113609460734546e-10, 
    1.1874767755957613e-10, 1.2905243114605339e-10, 1.4192640499418064e-10, 
    1.5708400258007805e-10, 1.7408372167504765e-10, 1.9234416566697509e-10, 
    2.1116966671749655e-10, 2.2978429695948363e-10, 2.4737203477180735e-10, 
    2.6312060598860561e-10, 2.7626589614499734e-10, 2.8613431314650085e-10, 
    2.9218014512362219e-10, 2.940157384568808e-10, 2.9143263601285707e-10, 
    2.8441251793892431e-10, 2.7312744863212139e-10, 2.579297425278627e-10, 
    2.3933231182686089e-10, 2.1798118972960731e-10, 1.9462220838360088e-10, 
    1.7006437551861288e-10, 1.4514233049808431e-10, 1.2068036182191552e-10, 
    9.7460017201382479e-11, 7.6192835347540942e-11, 5.7499070664492243e-11, 
    4.1892816676253949e-11, 2.9773155453210296e-11, 2.1420763540925588e-11, 
    1.6999032555533814e-11, 1.6558769464833598e-11, 2.0045647313741482e-11, 
    2.7309750784179155e-11, 3.8116694527588084e-11, 5.216015679226297e-11, 
    6.9075493302114728e-11, 8.8454241746374671e-11, 1.0985909204466005e-10, 
    1.3283880724849485e-10, 1.5694238419833372e-10, 1.817316130646415e-10, 
    2.0679124971557803e-10, 2.3173617968946082e-10, 2.5621517624937425e-10, 
    2.799112735955954e-10, 3.025391300462388e-10, 3.2384022060977794e-10, 
    3.4357687597633224e-10, 3.6152649280062849e-10, 3.7747712055127619e-10, 
    3.9122556679967188e-10, 4.0257876439491087e-10, 4.1135881477239346e-10, 
    4.1741151499472314e-10, 4.2061774710479884e-10, 4.2090663849620035e-10, 
    4.1826905227336778e-10, 4.1276968841196044e-10, 4.045562510082202e-10, 
    3.9386409606150037e-10, 3.8101531919884857e-10, 3.6641162241295219e-10, 
    3.5052100151664021e-10, 3.338588351820303e-10, 3.1696458450784275e-10, 
    3.0037578025165509e-10, 2.8460113568306483e-10, 2.7009485516211718e-10, 
    2.5723404755564825e-10, 2.4630072232389819e-10, 2.3746970164068479e-10, 
    2.3080297253860586e-10, 2.2625078838896474e-10, 2.2365910342322366e-10, 
    2.2278272271560567e-10, 2.2330300162675549e-10, 2.2484897993751838e-10, 
    2.2702038700319693e-10, 2.2941116823846647e-10, 2.3163205316289344e-10, 
    2.3333092993851377e-10, 2.3420970583303347e-10, 2.3403708007838159e-10, 
    2.3265640946412775e-10, 2.2998863835788936e-10, 2.2603033504633583e-10, 
    2.2084745378649864e-10, 2.1456548991995141e-10, 2.0735712166577064e-10, 
    1.9942832309897787e-10, 1.9100414464328024e-10, 1.8231501421466477e-10, 
    1.7358446227347094e-10, 1.6501877881365739e-10, 1.5679904432493943e-10, 
    1.4907555760489733e-10, 1.4196472508393849e-10, 1.3554816665416757e-10, 
    1.298737544272242e-10, 1.2495830249643779e-10, 1.2079142786224628e-10, 
    1.1734033053443651e-10, 1.1455497725665843e-10, 1.1237340243388268e-10, 
    1.1072674577387924e-10, 1.0954373475657704e-10, 1.0875436077445398e-10, 
    1.0829258512004509e-10, 1.0809802754160149e-10, 1.0811662233794894e-10, 
    1.0830040410567209e-10, 1.0860656786362398e-10, 1.0899611442279478e-10, 
    1.0943231715674714e-10, 1.0987929704633846e-10, 1.1030094897143506e-10, 
    1.1066036064642543e-10, 1.1091987681499847e-10, 1.1104176716289592e-10, 
    1.1098935633506445e-10, 1.1072859491173772e-10, 1.10229724393218e-10, 
    1.0946890841557575e-10, 1.0842949790993147e-10, 1.0710283634098995e-10, 
    1.0548840127517143e-10, 1.0359330220203612e-10, 1.0143108573601271e-10, 
    9.9020028752620039e-11, 9.6381094877154295e-11, 9.3535753444403319e-11, 
    9.0503961375276324e-11, 8.7302511704619646e-11, 8.3943987061237128e-11, 
    8.0436449267980327e-11, 7.6783924025855775e-11, 7.2987690648177251e-11, 
    6.9048190021887624e-11, 6.4967426333893532e-11, 6.0751572997402349e-11, 
    5.6413465066549206e-11, 5.1974679654658921e-11, 4.7466953039728642e-11, 
    4.2932670586938829e-11, 3.8424321593929252e-11, 3.4002876389186486e-11, 
    2.9735157453625126e-11, 2.569038029074487e-11, 2.1936177844143157e-11, 
    1.8534353957734388e-11, 1.553687003778114e-11, 1.2982280616650186e-11, 
    1.0893090669097881e-11, 9.2741632009912224e-12, 8.1124712351308e-12, 
    7.3780436059274208e-12, 7.0262493132293825e-12, 7.0010521049389459e-12, 
    7.2390695060430575e-12, 7.6740081830218818e-12, 8.2411782861942397e-12, 
    8.8816419662283373e-12, 9.5457547353067008e-12, 1.0195778977842021e-11, 
    1.0807441723218453e-11, 1.1370366609777146e-11, 1.1887447730606325e-11, 
    1.2373221235620257e-11, 1.2851506469820422e-11, 1.3352431503911938e-11, 
    1.3909256757073961e-11, 1.4555040661297356e-11, 1.5319557032379725e-11, 
    1.6226524960992617e-11, 1.7291443132943038e-11, 1.8519990333714821e-11, 
    1.9907285532100459e-11, 2.143786833570549e-11, 2.3086557681399947e-11, 
    2.482000630979392e-11, 2.6598996439816264e-11, 2.8381141811251336e-11, 
    3.0123987512202116e-11, 3.1788049633815253e-11, 3.3339683235269284e-11, 
    3.4753381364766271e-11, 3.6013384809093878e-11, 3.7114340748373971e-11, 
    3.8061037436358821e-11, 3.8867125703007993e-11, 3.9553131573294784e-11, 
    4.0143821292139214e-11, 4.0665404775161683e-11, 4.1142698457938554e-11, 
    4.1596784206630772e-11, 4.2043207438778681e-11, 4.2491089351293158e-11, 
    4.2943037745299552e-11, 4.3395972177843607e-11, 4.3842595627319908e-11, 
    4.4273404528339812e-11, 4.467882527740554e-11, 4.5051348087443665e-11, 
    4.538724757957055e-11, 4.5687810392588968e-11, 4.595981080933407e-11, 
    4.6215331156556147e-11, 4.647079682641937e-11, 4.6745511401222657e-11, 
    4.705972527052527e-11, 4.7432568961205424e-11, 4.7879919076315333e-11, 
    4.841256310799379e-11, 4.9034675565215745e-11, 4.9742853834010953e-11, 
    5.0525666232294144e-11, 5.13638508064695e-11, 5.2231057099951736e-11, 
    5.309512620090787e-11, 5.391977092772754e-11, 5.4666597139081939e-11, 
    5.5297337001065247e-11, 5.5776127536758469e-11, 5.6071716601534442e-11, 
    5.6159454120395341e-11, 5.6022957477207357e-11, 5.5655299428651448e-11, 
    5.5059633718977036e-11, 5.4249255937429244e-11, 5.3246990444156295e-11, 
    5.208405459971305e-11, 5.0798360121516721e-11, 4.9432486099538764e-11, 
    4.8031359914982174e-11, 4.6639918871894964e-11, 4.5300803484571618e-11, 
    4.405233346664133e-11, 4.2926817900495632e-11, 4.1949341563300112e-11, 
    4.1137002090067394e-11, 4.0498694151123298e-11, 4.0035355463324649e-11, 
    3.974065653140022e-11, 3.9601979257132844e-11, 3.9601716225583177e-11, 
    3.9718647480212597e-11, 3.99294398067411e-11, 4.0209982579472711e-11, 
    4.0536683316211866e-11, 4.088746276066951e-11, 4.1242552442546162e-11, 
    4.1584910136251495e-11, 4.1900430143018101e-11, 4.2177795792795138e-11, 
    4.2408200293164642e-11, 4.2584830194154282e-11, 4.2702348878096252e-11, 
    4.2756394079087749e-11, 4.2743168889273454e-11, 4.2659188393620765e-11, 
    4.2501234953513617e-11, 4.2266530270521451e-11, 4.1953074704955118e-11, 
    4.1560080815931645e-11, 4.1088484251043927e-11, 4.0541356273523184e-11, 
    3.9924242556551708e-11, 3.9245229984057431e-11, 3.8514826486345661e-11, 
    3.7745543949603173e-11, 3.6951282223233373e-11, 3.6146506184155528e-11, 
    3.5345378614986865e-11, 3.4560827661933437e-11, 3.3803762548655623e-11, 
    3.3082447983010358e-11, 3.2402094361509489e-11, 3.1764737094568687e-11, 
    3.116936230202798e-11, 3.0612267760639795e-11, 3.008761875568432e-11, 
    2.9588105458979331e-11, 2.9105655829706767e-11, 2.8632110598173675e-11, 
    2.8159825157324009e-11, 2.7682133695068875e-11, 2.7193683740889126e-11, 
    2.6690601977870523e-11, 2.6170514357076666e-11, 2.5632490841449309e-11, 
    2.5076864379353183e-11, 2.4505033617796704e-11, 2.3919247912889169e-11, 
    2.3322399246239776e-11, 2.2717856397256843e-11, 2.2109329990596953e-11, 
    2.1500787234865423e-11, 2.0896382570807403e-11, 2.0300420062381574e-11, 
    1.9717312940802319e-11, 1.915156243143213e-11, 1.8607670932113191e-11, 
    1.8090086478664121e-11, 1.7603091411205997e-11, 1.7150722874943979e-11, 
    1.6736609485217022e-11, 1.6363880625282791e-11, 1.6035050048904762e-11, 
    1.575191742747786e-11, 1.551548304116458e-11, 1.5325913460558833e-11, 
    1.5182478678570373e-11, 1.5083585712414698e-11, 1.5026758839851848e-11, 
    1.5008706006410648e-11, 1.5025356567075572e-11, 1.5071967143489328e-11, 
    1.5143182590117157e-11, 1.5233191227203814e-11, 1.533584011939349e-11, 
    1.5444831665175995e-11, 1.5553908835888867e-11, 1.5657116945694007e-11, 
    1.5749062535375176e-11, 1.5825229962197075e-11, 1.5882253506337877e-11, 
    1.5918223453409634e-11, 1.5932905094093876e-11, 1.592789390642949e-11, 
    1.590663590923658e-11, 1.5874318128278556e-11, 1.5837588811691159e-11, 
    1.5804144923305835e-11, 1.5782157068794292e-11, 1.5779637877317975e-11, 
    1.5803736680629341e-11, 1.5860124129530934e-11, 1.5952403009087837e-11, 
    1.6081738926849992e-11, 1.6246683701473148e-11, 1.6443255977854772e-11, 
    1.6665185178913623e-11, 1.6904432800387244e-11, 1.7151861080044063e-11, 
    1.7397976836957636e-11, 1.7633695865604873e-11, 1.7851059833623092e-11, 
    1.8043808996502149e-11, 1.8207783654404662e-11, 1.8341108264062319e-11, 
    1.8444172294749382e-11, 1.8519369293714266e-11, 1.8570709242567444e-11, 
    1.8603260866721972e-11, 1.8622574273223423e-11, 1.8634062594976817e-11, 
    1.8642485460856912e-11, 1.8651458965712789e-11, 1.8663169288321645e-11, 
    1.8678213673073617e-11, 1.8695632523685276e-11, 1.8713029907880104e-11, 
    1.8726902854743341e-11, 1.8733018120144879e-11, 1.8726861751851136e-11, 
    1.8704125448258593e-11, 1.8661156834877543e-11, 1.8595319668563209e-11, 
    1.850533686773011e-11, 1.8391431531516302e-11, 1.8255406904017369e-11, 
    1.8100595855054003e-11, 1.7931656395545894e-11, 1.7754333582392983e-11, 
    1.7575089106822338e-11, 1.7400730954803121e-11, 1.7238005556350182e-11, 
    1.7093198532658759e-11, 1.6971772392994216e-11, 1.6878032899024592e-11, 
    1.6814886343996168e-11, 1.6783616285449553e-11, 1.6783753211374523e-11, 
    1.681304879793137e-11, 1.6867489302460866e-11, 1.6941428211837199e-11, 
    1.7027793959511921e-11, 1.7118408194318252e-11, 1.7204384919933393e-11, 
    1.7276587490729953e-11, 1.7326184605530702e-11, 1.7345160211250701e-11, 
    1.7326872597050995e-11, 1.7266481614532778e-11, 1.7161344393329049e-11, 
    1.7011192258739971e-11, 1.6818193945906706e-11, 1.6586791589936815e-11, 
    1.6323404448557065e-11, 1.6035933348335021e-11, 1.5733193797155422e-11, 
    1.5424293985128295e-11, 1.511800189855663e-11, 1.4822207676690789e-11, 
    1.4543473827660186e-11, 1.4286755330880799e-11, 1.4055273692330189e-11, 
    1.3850545754198569e-11, 1.3672571520588539e-11, 1.3520090565529866e-11, 
    1.3390901263454994e-11, 1.3282199847642559e-11, 1.3190863087288425e-11, 
    1.3113687487462491e-11, 1.3047536693469843e-11, 1.2989420350806325e-11, 
    1.2936496174760061e-11, 1.2886059830087327e-11, 1.2835476845711026e-11, 
    1.2782166084349486e-11, 1.2723589110654456e-11, 1.2657300220149046e-11, 
    1.2581034756477367e-11, 1.2492847780687421e-11, 1.2391260554753297e-11, 
    1.227544057481037e-11, 1.2145339092117633e-11, 1.2001812673808122e-11, 
    1.1846688242483701e-11, 1.1682761125248407e-11, 1.1513727713229477e-11, 
    1.1344073804758184e-11, 1.1178859279356311e-11, 1.1023500182759332e-11, 
    1.0883482137993776e-11, 1.0764066958923544e-11, 1.0669973458315546e-11, 
    1.0605102283919696e-11, 1.0572262548896099e-11, 1.0572959857909997e-11, 
    1.0607232499485136e-11, 1.067361685933314e-11, 1.0769137421710583e-11, 
    1.0889439838474654e-11, 1.1028988046055073e-11, 1.1181351369145083e-11, 
    1.1339514913442484e-11, 1.1496255659111547e-11, 1.1644470809428725e-11, 
    1.177751654647732e-11, 1.188942411047694e-11, 1.1975113267168643e-11, 
    1.2030470153316393e-11, 1.2052373625682131e-11, 1.2038629007425133e-11, 
    1.1987930870767825e-11, 1.1899738019859407e-11, 1.1774213255632624e-11, 
    1.161216488585716e-11, 1.1415058771292432e-11, 1.1185044301167691e-11, 
    1.0925023515449977e-11, 1.0638738702649759e-11, 1.0330814400564392e-11, 
    1.0006805791278431e-11, 9.6731359822525264e-12, 9.3369870625011007e-12, 
    9.0061093799443545e-12, 8.6885482689504638e-12, 8.3923078217590641e-12, 
    8.1250011880098733e-12, 7.8934681453520479e-12, 7.7034590717444213e-12, 
    7.5593145951733036e-12, 7.4637635938953543e-12, 7.4177719318229388e-12, 
    7.4205263788624597e-12, 7.4694381323483113e-12, 7.5602888348880141e-12, 
    7.6873924730578553e-12, 7.8438591998380863e-12, 8.0218310222129471e-12, 
    8.2127884318853671e-12, 8.4078566020278027e-12, 8.5981356726869286e-12, 
    8.7749855124185625e-12, 8.9303827508717382e-12, 9.0571885046644889e-12, 
    9.149485921536548e-12, 9.202802206095195e-12, 9.2143646992311314e-12, 
    9.1832507430590678e-12, 9.1104934833945434e-12, 8.9990594163189514e-12, 
    8.85377490576721e-12, 8.6810883443453537e-12, 8.488785530672293e-12, 
    8.2855818647591027e-12, 8.080670336742607e-12, 7.8832221063380727e-12, 
    7.7019079069202668e-12, 7.5444358232955908e-12, 7.4171694103267502e-12, 
    7.3248467512661017e-12, 7.2704062248920139e-12, 7.2549425174506158e-12, 
    7.2777699371887672e-12, 7.3365908206352939e-12, 7.4277497218683519e-12, 
    7.5465276405778841e-12, 7.6874474321361296e-12, 7.8445997707261539e-12, 
    8.011901118646721e-12, 8.1833389179881535e-12, 8.3531416279011347e-12, 
    8.515918900444976e-12, 8.6667226990536561e-12, 8.8011304754587463e-12, 
    8.9152676073954536e-12, 9.0058365435034353e-12, 9.0701630399365703e-12, 
    9.1062293152030248e-12, 9.1127221746140072e-12, 9.0890953881895886e-12, 
    9.035629303193758e-12, 8.9534356288008438e-12, 8.8445004308687313e-12, 
    8.7116425099695811e-12, 8.5584830614850189e-12, 8.3893296187969802e-12, 
    8.2090722581995223e-12, 8.0230108987916683e-12, 7.8367081180937521e-12, 
    7.6557543200241161e-12, 7.4855954682594871e-12, 7.331305726651625e-12, 
    7.1974213296611888e-12, 7.0877183860524815e-12, 7.0050964379779461e-12, 
    6.9513901134175776e-12, 6.9273154311815379e-12, 6.93237292215663e-12, 
    6.9648897896989911e-12, 7.0220090910061025e-12, 7.0998448539674217e-12, 
    7.1936044198232352e-12, 7.2978485397384598e-12, 7.4067030163436834e-12, 
    7.5141806943574793e-12, 7.6144525966269158e-12, 7.7021558279503735e-12, 
    7.7726262666480907e-12, 7.8221437623966006e-12, 7.8480621573209394e-12, 
    7.8489225796957992e-12, 7.8244620481065843e-12, 7.7756057010968877e-12, 
    7.7043436618795123e-12, 7.6136207741506395e-12, 7.5071508405174342e-12, 
    7.3892412687942766e-12, 7.2645644181791018e-12, 7.1379723850309413e-12, 
    7.0142604458437542e-12, 6.8979527495183822e-12, 6.7931206543305829e-12, 
    6.7031800731479206e-12, 6.6307194944460969e-12, 6.5773462935598483e-12, 
    6.5435930365784305e-12, 6.5288490181857308e-12, 6.5313362396328983e-12, 
    6.5481774322284888e-12, 6.5754798438894695e-12, 6.6085066633530976e-12, 
    6.6419235990944041e-12, 6.6700383116710959e-12, 6.6871216685270145e-12, 
    6.6877226244403651e-12, 6.6669878786565229e-12, 6.6209665358805829e-12, 
    6.5468822590271466e-12, 6.4433549842370448e-12, 6.310536932969349e-12, 
    6.1501905007720919e-12, 5.9656860676219051e-12, 5.7618791341781404e-12, 
    5.5449384731373536e-12, 5.3220645321817213e-12, 5.1011580734869309e-12, 
    4.8904337092845582e-12, 4.6980019685070942e-12, 4.5314505573943516e-12, 
    4.397412229856104e-12, 4.3012315974361068e-12, 4.2466426207430358e-12, 
    4.2355562393031419e-12, 4.267911725426792e-12, 4.3416674108180128e-12, 
    4.4528834261853977e-12, 4.5959088899859949e-12, 4.7636905299700349e-12, 
    4.948148137095372e-12, 5.1406331445333773e-12, 5.3324340436800861e-12, 
    5.5152880706659126e-12, 5.6818762225379153e-12, 5.8262650367839584e-12, 
    5.9442769511971481e-12, 6.033686626214804e-12, 6.0943252812268969e-12, 
    6.1280077533165049e-12, 6.1382955220860568e-12, 6.1301182813925604e-12, 
    6.1092974919150297e-12, 6.0819846103743742e-12, 6.054097319802684e-12, 
    6.030781508819728e-12, 6.0159712292955293e-12, 6.0120819135457524e-12, 
    6.0198793056568414e-12, 6.0384949551453523e-12, 6.0656526902139356e-12, 
    6.0979782013583828e-12, 6.131460554668015e-12, 6.1619093309234088e-12, 
    6.1854403613183395e-12, 6.1988537361991354e-12, 6.1999360745277991e-12, 
    6.1876090967229499e-12, 6.1619326779090324e-12, 6.1239941169998387e-12, 
    6.0756509028350492e-12, 6.019239048222968e-12, 5.9572260624771441e-12, 
    5.8918959744224527e-12, 5.8250893098086243e-12, 5.7580366554057106e-12, 
    5.6912955608078256e-12, 5.6248195803774567e-12, 5.5580801177641218e-12, 
    5.4903215956373009e-12, 5.4208364186501122e-12, 5.3491840831294749e-12, 
    5.2754479051654708e-12, 5.2003768011740818e-12, 5.1254264588925655e-12, 
    5.052702594339435e-12, 4.9848077892425266e-12, 4.9245822356767284e-12, 
    4.8748180388501087e-12, 4.8379314451899999e-12, 4.8156998138998114e-12, 
    4.8089967553089275e-12, 4.8176843189529852e-12, 4.8405562015345218e-12, 
    4.875431795071547e-12, 4.9192914350730579e-12, 4.9685588303849402e-12, 
    5.0193509119421948e-12, 5.0678038454511275e-12, 5.1103366410810683e-12, 
    5.1438915248805502e-12, 5.1661040327351726e-12, 5.1754042544876559e-12, 
    5.1710350468511121e-12, 5.1530338277271705e-12, 5.1221237016948904e-12, 
    5.0795923651766413e-12, 5.0271715803071682e-12, 4.9668687494602011e-12, 
    4.900837862915663e-12, 4.8312469399957064e-12, 4.7601554874969946e-12, 
    4.68941468546465e-12, 4.6205715404250448e-12, 4.5547821256275968e-12, 
    4.4927596618580587e-12, 4.4347199379587887e-12, 4.3803534684246121e-12, 
    4.3288409045032263e-12, 4.2789036137818476e-12, 4.2288840692816972e-12, 
    4.1768936934547417e-12, 4.1209489682447725e-12, 4.0592043340392508e-12, 
    3.9901161132729641e-12, 3.9126607758792353e-12, 3.8264889803241791e-12, 
    3.7320357581929076e-12, 3.6305813045878143e-12, 3.5242466519584609e-12, 
    3.4158870224948728e-12, 3.3089748200796552e-12, 3.2073876318079735e-12, 
    3.1151951579997186e-12, 3.0364135117374816e-12, 2.974778582232652e-12, 
    2.9335311093764854e-12, 2.9152542454681373e-12, 2.9217453162690083e-12, 
    2.9539173292100751e-12, 3.0117670807669095e-12, 3.0943865145118774e-12, 
    3.1999838573383462e-12, 3.3259711591977468e-12, 3.4690714924178217e-12, 
    3.6254409510745606e-12, 3.790830465796804e-12, 3.9607821364716501e-12, 
    4.1308242395994369e-12, 4.2966886051954539e-12, 4.454504335926659e-12, 
    4.6009938390544715e-12, 4.7336334944551255e-12, 4.8507199343473389e-12, 
    4.9513927924301713e-12, 5.0355970536131136e-12, 5.1039317908174069e-12, 
    5.1574612821293554e-12, 5.197467067407392e-12, 5.2251880257236695e-12, 
    5.2415707518238968e-12, 5.2470629439945716e-12, 5.2414863514106899e-12, 
    5.2239970893111401e-12, 5.1931470859376827e-12, 5.1470359608188014e-12, 
    5.0835721845450164e-12, 5.0007455673489593e-12, 4.8969455794185217e-12, 
    4.7712893605938527e-12, 4.6238495329859854e-12, 4.4558511781167092e-12, 
    4.2697236833650641e-12, 4.0690889522268681e-12, 3.8585436877807187e-12, 
    3.6434743411880463e-12, 3.4296607309056723e-12, 3.2229149647465471e-12, 
    3.0286434790517515e-12, 2.8515064810156785e-12, 2.6950452832425967e-12, 
    2.5615078963913729e-12, 2.4516855839435401e-12, 2.3649706503454951e-12, 
    2.2994489455527822e-12, 2.252198813290847e-12, 2.2195785476542964e-12, 
    2.1976484182014037e-12, 2.1825124825441154e-12, 2.1707345671958036e-12, 
    2.1595801544820927e-12, 2.1472443845579223e-12, 2.132897922986957e-12, 
    2.1166896913060904e-12, 2.09958346578162e-12, 2.0831408014060822e-12, 
    2.0692258676165686e-12, 2.0597182983331304e-12, 2.0561776233253091e-12, 
    2.0596234022310447e-12, 2.0703100612215644e-12, 2.0876459490612158e-12, 
    2.1101641423050537e-12, 2.1356302417285465e-12, 2.161200155086228e-12, 
    2.1837007291239656e-12, 2.1999211486309596e-12, 2.2069559662663821e-12, 
    2.2025417671285802e-12, 2.1853444076471714e-12, 2.1551803358275275e-12, 
    2.1131767660420813e-12, 2.061782935351254e-12, 2.0046887943575879e-12, 
    1.9466085875741739e-12, 1.8929985914809122e-12, 1.8496485910353137e-12, 
    1.8222813599937701e-12, 1.8160779518771326e-12, 1.8353213917583758e-12, 
    1.8830130154461405e-12, 1.9606610748674205e-12, 2.068143513329464e-12, 
    2.2037110112966334e-12, 2.3641033868153173e-12, 2.5447891371014646e-12, 
    2.7402702455422103e-12, 2.9444536207921885e-12, 3.1510340807764366e-12, 
    3.3538766316881207e-12, 3.5473356129671111e-12, 3.7265302357881905e-12, 
    3.8875307578151404e-12, 4.0274665210780007e-12, 4.1445162287965167e-12, 
    4.2378730582730426e-12, 4.3075802906834517e-12, 4.3543693727124088e-12, 
    4.3794264532479711e-12, 4.3841727955014149e-12, 4.3700234644509592e-12, 
    4.3381976895339888e-12, 4.2895666738372966e-12, 4.2245372417196124e-12, 
    4.1430235369910011e-12, 4.0445060364173816e-12, 3.9281152941223887e-12, 
    3.7928674774941135e-12, 3.6378605207917161e-12, 3.4625800310636798e-12, 
    3.2671668517624988e-12, 3.0526734459033962e-12, 2.8212483466444213e-12, 
    2.576254806411729e-12, 2.322263407748865e-12, 2.0649383433784565e-12, 
    1.81079358458647e-12, 1.5668685018520827e-12, 1.3403073776768712e-12, 
    1.1379238956257896e-12, 9.6575368972450183e-13, 8.2865994387036709e-13, 
    7.2999341924783879e-13, 6.7140777708949982e-13, 6.5278402417077786e-13, 
    6.7223260308834217e-13, 7.2631287741570212e-13, 8.102395108798034e-13, 
    9.1829380444518025e-13, 1.0441221995285594e-12, 1.1812175782496369e-12, 
    1.3232034338649508e-12, 1.4642464791956825e-12, 1.5992390598700657e-12, 
    1.7240849877687864e-12, 1.8357156742993345e-12, 1.9322358134209104e-12, 
    2.0128033665546709e-12, 2.0776369547550706e-12, 2.1278186752669695e-12, 
    2.1652011157958227e-12, 2.1921648740273812e-12, 2.2115071476374127e-12, 
    2.2261791053179918e-12, 2.239175616457159e-12, 2.2533177683379127e-12, 
    2.2711404048405549e-12, 2.2947418867992854e-12, 2.3257163684782381e-12, 
    2.3650273921759783e-12, 2.4129998843704008e-12, 2.4692623169632748e-12, 
    2.5327903126153234e-12, 2.6019174786594099e-12, 2.6744464252818547e-12, 
    2.7477446776203713e-12, 2.8189171854236343e-12, 2.8849883721401374e-12, 
    2.9431177210332582e-12, 2.9908071385307747e-12, 3.0261257668914624e-12, 
    3.0478799043511704e-12, 3.0557714244446634e-12, 3.0504463309218031e-12, 
    3.0335065945981331e-12, 3.0074197463871319e-12, 2.9753640928027103e-12, 
    2.9409817428123652e-12, 2.9081129467722107e-12, 2.8804676865941444e-12, 
    2.8613342084796905e-12, 2.8532759810666927e-12, 2.8579398601291757e-12, 
    2.875855695767151e-12, 2.9064230887512874e-12, 2.9478993912402216e-12, 
    2.9975602160590065e-12, 3.0518668826229175e-12, 3.1067618364581679e-12, 
    3.1579568297135536e-12, 3.2012816226305436e-12, 3.2329723205666474e-12, 
    3.2499883272038901e-12, 3.2502040568644653e-12, 3.2325993090280109e-12, 
    3.1972937477135853e-12, 3.145566161861142e-12, 3.079712875582437e-12, 
    3.0029037263305238e-12, 2.9188968837461048e-12, 2.8317739559853824e-12, 
    2.745626316628045e-12, 2.6642573333638819e-12, 2.5908980293115043e-12, 
    2.5279995274962948e-12, 2.4770638580020933e-12, 2.4385896415578446e-12, 
    2.412058323082664e-12, 2.3960393576023678e-12, 2.3883424907037365e-12, 
    2.3862373138172433e-12, 2.3866954308225046e-12, 2.3866613013360532e-12, 
    2.3832891094267356e-12, 2.3741852330795941e-12, 2.3575510167829388e-12, 
    2.3323077848869487e-12, 2.2981216525792922e-12, 2.2553965545250716e-12, 
    2.2051727580770596e-12, 2.1490098999842479e-12, 2.0888305970536788e-12, 
    2.0267571886485218e-12, 1.9649505917001254e-12, 1.9055080266256645e-12, 
    1.8503160241528821e-12, 1.8010195059817009e-12, 1.7589633501517094e-12, 
    1.725204816484429e-12, 1.7004984467184881e-12, 1.6853416499973657e-12, 
    1.6799696873435992e-12, 1.68440009238395e-12, 1.6984484751098129e-12, 
    1.7216942304605919e-12, 1.7535475579876538e-12, 1.7932532276498459e-12, 
    1.839893231226281e-12, 1.8924357624287517e-12, 1.9497424919343274e-12, 
    2.0106253335296256e-12, 2.0738460757702439e-12, 2.1381551619237127e-12, 
    2.2022782382933296e-12, 2.2649042905060675e-12, 2.324652342010281e-12, 
    2.3800585695104755e-12, 2.4295126706627485e-12, 2.4712616882008917e-12, 
    2.503407664414554e-12, 2.5239552411780135e-12, 2.5308953646676189e-12, 
    2.5223350757117484e-12, 2.4966462119089691e-12, 2.4526486031033531e-12, 
    2.3897798940796219e-12, 2.3082480495387968e-12, 2.2091284953600594e-12, 
    2.0944060065300254e-12, 1.9669204017256216e-12, 1.8302542278685107e-12, 
    1.6885086915259039e-12, 1.5460435705904649e-12, 1.4071689532106805e-12, 
    1.2758415304475056e-12, 1.1553573240412804e-12, 1.0481351847427423e-12, 
    9.5555063879870655e-13, 8.7788658131485174e-13, 8.1437285393784755e-13, 
    7.6332590568561624e-13, 7.2236514031396787e-13, 6.8869627339412745e-13, 
    6.5940511480371731e-13, 6.3176587309358677e-13, 6.0351935333954539e-13, 
    5.7309137465965306e-13, 5.3974850251252187e-13, 5.0369433489048935e-13, 
    4.6604413317320095e-13, 4.2877793219437726e-13, 3.9458691341872788e-13, 
    3.6668572640423192e-13, 3.4859810196893605e-13, 3.4390027121216174e-13, 
    3.5597756931712755e-13, 3.877860343187298e-13, 4.416365062191617e-13, 
    5.1903644583726481e-13, 6.2055714906004313e-13, 7.4576922983987175e-13, 
    8.9325054010782387e-13, 1.0606194946510116e-12, 1.2446711950666941e-12, 
    1.4415206380042719e-12, 1.6467961944606124e-12, 1.8558293839353086e-12, 
    2.0638786175313845e-12, 2.2662978744978102e-12, 2.4587054005931288e-12, 
    2.6370958365622855e-12, 2.7979268616126179e-12, 2.9381669490089117e-12, 
    3.055311250647731e-12, 3.1473785844853179e-12, 3.2129210764941732e-12, 
    3.2510036968501022e-12, 3.2612457313558402e-12, 3.2438300564442846e-12, 
    3.1995600062086139e-12, 3.1299056187405093e-12, 3.0370538679031862e-12, 
    2.9239214653990923e-12, 2.794165864755896e-12, 2.6521322645261099e-12, 
    2.5027409577813103e-12, 2.35133899068643e-12, 2.2034802578707067e-12, 
    2.0646901242194649e-12, 1.9401633719637887e-12, 1.8345333596272451e-12, 
    1.751549456275454e-12, 1.6938866591954513e-12, 1.6629988461959901e-12, 
    1.6590320552994815e-12, 1.6808216057390235e-12, 1.7259833186922543e-12, 
    1.7911019479863191e-12, 1.8719711959002025e-12, 1.9638482918712377e-12, 
    2.0617872725161583e-12, 2.1609112851825581e-12, 2.2566847809810724e-12, 
    2.3451329945167751e-12, 2.4230129818025099e-12, 2.4878881880464901e-12, 
    2.5381695658423824e-12, 2.5730896493069871e-12, 2.5926434100076326e-12, 
    2.597461950356781e-12, 2.5887176317336219e-12, 2.5679781905009861e-12, 
    2.5370965255759251e-12, 2.4980784127704724e-12, 2.4529852792652972e-12, 
    2.403828872267795e-12, 2.3524936863983573e-12, 2.3006505969369775e-12, 
    2.2496937677361216e-12, 2.2006948721607457e-12, 2.1543373190356432e-12, 
    2.1109228781505594e-12, 2.0703656772330085e-12, 2.0322066592878505e-12, 
    1.9956818096780278e-12, 1.9597886814827042e-12, 1.9233977376083606e-12, 
    1.8853515346388343e-12, 1.8445859718933334e-12, 1.800231175338067e-12, 
    1.7517083474885725e-12, 1.6987824281753761e-12, 1.6415894557255394e-12, 
    1.5806385933602925e-12, 1.5167793245257985e-12, 1.4511223570975317e-12, 
    1.3849735237394516e-12, 1.3197410854605931e-12, 1.2568646336212748e-12, 
    1.197735530325273e-12, 1.1436491265188587e-12, 1.095781177277712e-12, 
    1.0551824345784241e-12, 1.0227696741832899e-12, 9.9933281698978344e-13, 
    9.8554461702072047e-13, 9.819345311626319e-13, 9.8885116056899617e-13, 
    1.006407386696178e-12, 1.0343792340114862e-12, 1.0721286176520046e-12, 
    1.1185107604170498e-12, 1.1717954898260211e-12, 1.2296548703173815e-12, 
    1.2891715495166791e-12, 1.3469330766480729e-12, 1.3991955924331325e-12, 
    1.4420810226051744e-12, 1.471847808367423e-12, 1.4851621447190281e-12, 
    1.4793820817780968e-12, 1.4527956670832207e-12, 1.4048303737476368e-12, 
    1.3361281055411171e-12, 1.248569958656025e-12, 1.1452116256519276e-12, 
    1.0301069650223316e-12, 9.0804486931504566e-13, 7.8425272543825212e-13, 
    6.6406154891765758e-13, 5.5255676880392484e-13, 4.5426452909238012e-13, 
    3.7287103442232201e-13, 3.1101042723855612e-13, 2.7014334340343148e-13, 
    2.5047397725288175e-13, 2.5101552025216046e-13, 2.6965966937015059e-13, 
    3.0338836266545641e-13, 3.484694614556176e-13, 4.0073568701497035e-13, 
    4.5586164035042822e-13, 5.0967257914126223e-13, 5.5837924576694114e-13, 
    5.9884672532466521e-13, 6.2876633415593977e-13, 6.4679851320332251e-13, 
    6.5263250889163102e-13, 6.4698981572796616e-13, 6.3152740243864038e-13, 
    6.0870966066339686e-13, 5.8158763417666274e-13, 5.5356979954617382e-13, 
    5.2813580267575885e-13, 5.0855928330848075e-13, 4.976710147309753e-13, 
    4.9763128102698961e-13, 5.0978229512208017e-13, 5.3455980331515883e-13, 
    5.7150038492613842e-13, 6.1930060034250633e-13, 6.7599206317669757e-13, 
    7.3910424759479171e-13, 8.059377634916164e-13, 8.7378602206513873e-13, 
    9.4019339734636562e-13, 1.0031299838918862e-12, 1.061180789353115e-12, 
    1.1136071119242004e-12, 1.160379547354624e-12, 1.2021177837561105e-12, 
    1.2399773751470247e-12, 1.2754774638152639e-12, 1.3102973798668539e-12, 
    1.3460315168833574e-12, 1.3839973783458513e-12, 1.4250214016946486e-12, 
    1.4692920712016245e-12, 1.5162740073452926e-12, 1.5646853194118596e-12, 
    1.6125588114512259e-12, 1.6573852832037479e-12, 1.6963057801325887e-12, 
    1.726362263956804e-12, 1.744772659592448e-12, 1.7492043347541658e-12, 
    1.7380175868310992e-12, 1.7104660608824746e-12, 1.6668196443499301e-12, 
    1.6083873850229528e-12, 1.5374952134057104e-12, 1.4573077293453157e-12, 
    1.371641510678742e-12, 1.2846846985218818e-12, 1.2007087975835624e-12, 
    1.123773256738747e-12, 1.0574649892345035e-12, 1.0046571185200366e-12, 
    9.6738215283170974e-13, 9.467360369276514e-13, 9.4289507298289659e-13, 
    9.5516872033303601e-13, 9.8213804073617226e-13, 1.0218265089967004e-12, 
    1.071918337882032e-12, 1.1299092599666816e-12, 1.1933187850618818e-12, 
    1.2598281353367232e-12, 1.3273897862522283e-12, 1.394287596388224e-12, 
    1.4591429713514019e-12, 1.5208958511396878e-12, 1.5787405576697141e-12, 
    1.6320556935910547e-12, 1.6803264361173992e-12, 1.7230842551653683e-12, 
    1.7598609567523796e-12, 1.7901945057762727e-12, 1.8136428143340326e-12, 
    1.8298690008519847e-12, 1.8387188427393804e-12, 1.8403204109646145e-12, 
    1.8351759429193989e-12, 1.8242463039664574e-12, 1.8089527694636883e-12, 
    1.7911898401181283e-12, 1.7732420141951053e-12, 1.7576279946232831e-12, 
    1.7469439607493586e-12, 1.7436421659237293e-12, 1.7498009608513598e-12, 
    1.7669242411226936e-12, 1.7957745222480738e-12, 1.8362521221738231e-12, 
    1.8873621571709953e-12, 1.9472322286229207e-12, 2.0132336913291834e-12, 
    2.0821541942244254e-12, 2.1504146204358773e-12, 2.2143312466510626e-12, 
    2.2703634553455162e-12, 2.3153414209012039e-12, 2.3466667368027912e-12, 
    2.362458753202446e-12, 2.361606977118691e-12, 2.3438157460500425e-12, 
    2.3095541140628248e-12, 2.2599528366781031e-12, 2.1966760152788418e-12, 
    2.1217896046673652e-12, 2.0375753426119718e-12, 1.9464071685054011e-12, 
    1.8506136120605009e-12, 1.7523564345596801e-12, 1.6535511428709936e-12, 
    1.5558266111812755e-12, 1.4604853162927975e-12, 1.3685169116176729e-12, 
    1.2806101181092414e-12, 1.1972010579441477e-12, 1.1185135854346151e-12, 
    1.0446257917271982e-12, 9.7553068991655361e-13, 9.1118316127995501e-13, 
    8.5156014781491309e-13, 7.966964736724242e-13, 7.4671925186346086e-13, 
    7.0184570051062411e-13, 6.62380463640591e-13, 6.2869372410315451e-13, 
    6.0117214693370153e-13, 5.8017245220972278e-13, 5.6596653672551477e-13, 
    5.5867350734269255e-13, 5.5820862682574131e-13, 5.6426418306056886e-13, 
    5.7628561616425972e-13, 5.9349475451769028e-13, 6.149090891712086e-13, 
    6.3944137130308219e-13, 6.6596718142894115e-13, 6.9343012208529934e-13, 
    7.2094674484201423e-13, 7.4789355134298234e-13, 7.7395996620873904e-13, 
    7.9919721519107942e-13, 8.2398830924062318e-13, 8.4898588744066075e-13, 
    8.7501728842746323e-13, 9.0293384664749683e-13, 9.3345985160666249e-13, 
    9.6703920035208776e-13, 1.0036731313157181e-12, 1.0428413355810589e-12, 
    1.0834327114657725e-12, 1.1237665490415812e-12, 1.1616636597669177e-12, 
    1.1945646217080376e-12, 1.2197265188624698e-12, 1.2344184476724008e-12, 
    1.23611715095237e-12, 1.2227334833611044e-12, 1.1927339565021541e-12, 
    1.145281822283943e-12, 1.0802915198910636e-12, 9.9842274851489079e-13, 
    9.0104187497620234e-13, 7.9013615118884615e-13, 6.6820352770411808e-13, 
    5.3813197035284699e-13, 4.0305888769189254e-13, 2.6627605508129421e-13, 
    1.3109711430074868e-13, 7.7768015992495243e-16, -1.2156312415052461e-13, 
    -2.3304305452064568e-13, -3.310634490818556e-13, -4.1339604549319411e-13, 
    -4.7824830084169316e-13, -5.2432000363033206e-13, 
    -5.5087112246727192e-13, -5.5775654519327988e-13, 
    -5.4544027778135604e-13, -5.1499737304274762e-13, 
    -4.6809568323881667e-13, -4.0688610689574798e-13, 
    -3.3393068327964198e-13, -2.5207216547268446e-13, 
    -1.6429728529840527e-13, -7.3572362743409782e-14, 1.727981248582551e-14, 
    1.0574904136824208e-13, 1.8971846020412635e-13, 2.6757696703969006e-13, 
    3.3826241651464713e-13, 4.012984973017782e-13, 4.5674738189501019e-13, 
    5.0521695947779375e-13, 5.4776927645357321e-13, 5.8583060838049201e-13, 
    6.2108389439192744e-13, 6.5535865478595522e-13, 6.9050214302373013e-13, 
    7.2826314175825245e-13, 7.7016848761707905e-13, 8.1741311507976118e-13, 
    8.7079798558632062e-13, 9.3064929870205959e-13, 9.9679752950697085e-13, 
    1.0685806020426468e-12, 1.1448816707121292e-12, 1.2241924437055756e-12, 
    1.3047164227284286e-12, 1.38448143462852e-12, 1.4614862664068107e-12, 
    1.5338186743612878e-12, 1.5998019661323755e-12, 1.6580869724960289e-12, 
    1.7077486546861338e-12, 1.7483141234418153e-12, 1.77977517324923e-12, 
    1.8025337235580355e-12, 1.8173294137873739e-12, 1.8251115009858096e-12, 
    1.8268980944752477e-12, 1.823623850019339e-12, 1.8159717279587578e-12, 
    1.8042764154976559e-12, 1.7884192309232291e-12, 1.7677992982428418e-12, 
    1.7413517068715473e-12, 1.7076481485014307e-12, 1.665039384232949e-12, 
    1.6118542435462953e-12, 1.5466164034408151e-12, 1.4682836664644402e-12, 
    1.3764481620182505e-12, 1.2715129869401266e-12, 1.15477818637589e-12, 
    1.0284890654402356e-12, 8.9575022912146357e-13, 7.6039984099785881e-13, 
    6.2677682027833802e-13, 4.9946463450942061e-13, 3.8297337074817055e-13, 
    2.8145737069964768e-13, 1.9839810780258624e-13, 1.3640501609357858e-13, 
    9.7052316892504682e-14, 8.0755004902766682e-14, 8.6787847633217959e-14, 
    1.1337199398267643e-13, 1.5781114571520533e-13, 2.1670393658429097e-13, 
    2.8618824323258895e-13, 3.6219135690963299e-13, 4.4068441655859148e-13, 
    5.17898890421018e-13, 5.9051531584059588e-13, 6.5577355874815843e-13, 
    7.1155638744738324e-13, 7.5638843918352366e-13, 7.8940544006952455e-13, 
    8.1028259017935901e-13, 8.1912768024737878e-13, 8.1638184086715092e-13, 
    8.0273379577111164e-13, 7.7902463429346596e-13, 7.4620420900198052e-13, 
    7.0530740942008515e-13, 6.5748485443680275e-13, 6.0399521632045525e-13, 
    5.4623829695944404e-13, 4.8580170314526237e-13, 4.2446158766306378e-13, 
    3.6415467604196287e-13, 3.069266863544022e-13, 2.5486053143772475e-13, 
    2.0997003481014265e-13, 1.7406532309736452e-13, 1.4863903989377513e-13, 
    1.3475558428003339e-13, 1.3296319309656957e-13, 1.4324838064085683e-13, 
    1.6502438034380111e-13, 1.9717990897842187e-13, 2.3816240281229013e-13, 
    2.8608569526646166e-13, 3.3887184857725511e-13, 3.9440437937103356e-13, 
    4.5069427811174559e-13, 5.0600031342911976e-13, 5.5897320126832155e-13, 
    6.0871985370029268e-13, 6.5488107175374508e-13, 6.9763180865061855e-13, 
    7.3765338996260991e-13, 7.7606289967635426e-13, 8.1430557958811879e-13, 
    8.5400631732515838e-13, 8.9680106705893414e-13, 9.4415253925749851e-13, 
    9.9719711180601302e-13, 1.0565418024470223e-12, 1.1221446358771877e-12, 
    1.1932393900599066e-12, 1.2682875295199607e-12, 1.3450083633257514e-12, 
    1.4204592817036809e-12, 1.4911733467221802e-12, 1.553371570722351e-12, 
    1.6031556721542139e-12, 1.6367742409521494e-12, 1.6508519165125545e-12, 
    1.6426234537852929e-12, 1.6101347533781744e-12, 1.5524137740752373e-12, 
    1.4695666729760359e-12, 1.3628567843886452e-12, 1.2346991539653882e-12, 
    1.0886112111209126e-12, 9.291079423117711e-13, 7.6155841807272945e-13, 
    5.9195877987758956e-13, 4.2668663302023204e-13, 2.7223659038075736e-13, 
    1.3491489608082387e-13, 2.0522101096431011e-14, -6.5936755874051375e-14, 
    -1.205229736359843e-13, -1.4058947858066674e-13, -1.2493833695198822e-13, 
    -7.3905441878030755e-14, 1.0649531713558037e-14, 1.2541773462145442e-13, 
    2.658494288174259e-13, 4.2637636675718051e-13, 6.007266455220634e-13, 
    7.8226322235681724e-13, 9.6433270727945448e-13, 1.1405948981166005e-12, 
    1.3053249564159216e-12, 1.4536386102269102e-12, 1.5816847039739377e-12, 
    1.6867238578723596e-12, 1.7671726494300945e-12, 1.8225495235256276e-12, 
    1.853403576820571e-12, 1.8611497121903362e-12, 1.8479559680948415e-12, 
    1.8165592813008672e-12, 1.7701123823734714e-12, 1.7120388987214179e-12, 
    1.6459172597356637e-12, 1.5753629875376955e-12, 1.5039333273668149e-12, 
    1.4350512424746409e-12, 1.3718887100253529e-12, 1.3173019665149836e-12, 
    1.27371826958711e-12, 1.2430251456676169e-12, 1.2264731887824867e-12, 
    1.2245497689174586e-12, 1.236930450482782e-12, 1.2624052686811362e-12, 
    1.2989025229474764e-12, 1.343516342343444e-12, 1.3926534320235129e-12, 
    1.4422169321966023e-12, 1.4878205152139751e-12, 1.5250728350488913e-12, 
    1.5498816191932811e-12, 1.5587131056416102e-12, 1.5488584896485347e-12, 
    1.5186197503396256e-12, 1.4674145574038874e-12, 1.3958143182113713e-12, 
    1.3054666023396963e-12, 1.1989319822862563e-12, 1.0795037810784983e-12, 
    9.5093157391773511e-13, 8.171434969723687e-13, 6.8198901344263122e-13, 
    5.4901457961646139e-13, 4.2127048676728621e-13, 3.0121273989885346e-13, 
    1.9064141452365217e-13, 9.0708673976656228e-14, 1.9677528315253666e-15, 
    -7.5525194957727274e-14, -1.4212262930220883e-13, 
    -1.9844955955814427e-13, -2.4531437790212798e-13, -2.835923260509743e-13, 
    -3.141643401693155e-13, -3.3781313194614382e-13, -3.5519734619083851e-13, 
    -3.6677419911548443e-13, -3.7280451900700565e-13, 
    -3.7329284016573572e-13, -3.6800541675109886e-13, 
    -3.5648404747038311e-13, -3.3809513570356138e-13, 
    -3.1207273032465946e-13, -2.7765147811560165e-13, 
    -2.3414072872774039e-13, -1.8109141723538449e-13, 
    -1.1836951924165498e-13, -4.6340231910532714e-14, 3.4127440626731854e-14, 
    1.2159567804848452e-13, 2.1404918639105187e-13, 3.0897514056813177e-13, 
    4.0350412440720292e-13, 4.9453976681334733e-13, 5.789922844600597e-13, 
    6.5397211484945093e-13, 7.1701388271102746e-13, 7.6625681236635609e-13, 
    8.0061302846107109e-13, 8.1984108837160632e-13, 8.2461983275477116e-13, 
    8.1648720584107166e-13, 7.9775606919412327e-13, 7.7133813098479789e-13, 
    7.4055778044275135e-13, 7.088817506374907e-13, 6.7968603094507402e-13, 
    6.5599708519460206e-13, 6.4029044175943807e-13, 6.3431163869781608e-13, 
    6.3900574006369412e-13, 6.5448120194637985e-13, 6.8008240975480166e-13, 
    7.1450976619903216e-13, 7.5600291466281373e-13, 8.0255139024161788e-13, 
    8.5211416259232482e-13, 9.0280863081680049e-13, 9.5307690006182957e-13, 
    1.0017759595701902e-12, 1.0482204676628125e-12, 1.0921265507161536e-12, 
    1.1335526430043747e-12, 1.1727602935704294e-12, 1.2100498094102786e-12, 
    1.2456219506703493e-12, 1.2794578569494423e-12, 1.3112298716486535e-12, 
    1.3402611268478811e-12, 1.3655475887319143e-12, 1.3858305874514077e-12, 
    1.3997085587566077e-12, 1.4057732921534409e-12, 1.4027680948969009e-12, 
    1.3897262285857337e-12, 1.3660949432660736e-12, 1.3318254725726589e-12, 
    1.2873981274161288e-12, 1.2338389050022624e-12, 1.1726481821861027e-12, 
    1.1057154606628045e-12, 1.0351794227862826e-12, 9.6329099777170932e-13, 
    8.9225221353855881e-13, 8.2406338294110509e-13, 7.6037062547110387e-13, 
    7.0238053464909909e-13, 6.5075153459669006e-13, 6.0557835173562656e-13, 
    5.6637896763879277e-13, 5.3215900316775334e-13, 5.0149745554559985e-13, 
    4.7268158739193244e-13, 4.4387299914721518e-13, 4.1328815783416356e-13, 
    3.7938764326345015e-13, 3.4105200511301767e-13, 2.9772455495352558e-13, 
    2.4951574184239397e-13, 1.9723903700746597e-13, 1.423883148695847e-13, 
    8.7042484973550757e-14, 3.3700294324783376e-14, -1.4923605422824563e-14, 
    -5.6137716561588187e-14, -8.753475067965298e-14, -1.0719905754295663e-13, 
    -1.1390146174311039e-13,
  // Sqw-total(1, 0-1999)
    0.11872223080445742, 0.11819878894488221, 0.11664584873709521, 
    0.11411453152502088, 0.11068667929133567, 0.10647011566303145, 
    0.10159257945337803, 0.096194822911686365, 0.090423410694380368, 
    0.084423745282931228, 0.07833378487368324, 0.072278820993778387, 
    0.066367559390134542, 0.060689614797853793, 0.055314403068853941, 
    0.050291305347961196, 0.045650897226846295, 0.041406985410920805, 
    0.037559175472832357, 0.034095703251311976, 0.030996293397835155, 
    0.028234854188561111, 0.025781870559140951, 0.023606410707497194, 
    0.021677710262214461, 0.01996633835086048, 0.018444980061602209, 
    0.017088889427685928, 0.015876077009235309, 0.014787298012823604, 
    0.013805902684514417, 0.012917602512763212, 0.012110195482933879, 
    0.011373282802086278, 0.01069799932283097, 0.010076771089459518, 
    0.0095031063910774212, 0.0089714215211182235, 0.0084768989826606855, 
    0.0080153738846563197, 0.0075832434246572945, 0.0071773943222284958, 
    0.0067951435589651129, 0.00643418855382576, 0.0060925637744397489, 
    0.005768601631936523, 0.005460896253501186, 0.0051682693360487943, 
    0.0048897377456499436, 0.0046244828474642195, 0.004371821746761503, 
    0.0041311807149462367, 0.0039020710887662951, 0.0036840678890072772, 
    0.0034767913278346122, 0.003279891279420283, 0.0030930346906689007, 
    0.0029158958178301031, 0.0027481490967576879, 0.0025894643925479985, 
    0.0024395043289416529, 0.0022979233686374473, 0.0021643683015587314, 
    0.002038479798291339, 0.0019198946997170069, 0.0018082487405910793, 
    0.0017031794431628918, 0.0016043289646492757, 0.0015113467359653546, 
    0.0014238917841188502, 0.0013416346821293454, 0.0012642591136331066, 
    0.0011914630710194534, 0.0011229597243962895, 0.0010584780043826462, 
    0.00099776293714196529, 0.00094057575907589678, 0.00088669382567531287, 
    0.00083591031834089524, 0.00078803374764010439, 0.00074288725298039533, 
    0.00070030770687951765, 0.00066014464523526451, 0.00062225906057044157, 
    0.00058652211007346382, 0.00055281380149482036, 0.00052102172538563143, 
    0.0004910399005578983, 0.00046276779085294883, 0.00043610953619607144, 
    0.00041097342116339439, 0.00038727158212533905, 0.00036491993193643607, 
    0.00034383826156492603, 0.00032395046313263721, 0.00030518481017415884, 
    0.00028747422940616731, 0.00027075650398528778, 0.00025497436033098352, 
    0.00024007540754182485, 0.00022601191808972978, 0.00021274045838405155, 
    0.00020022139550986788, 0.00018841831987680477, 0.00017729743121213038, 
    0.00016682693667978291, 0.00015697650518309094, 0.00014771681221719592, 
    0.00013901919669510421, 0.00013085543703303135, 0.00012319764048611699, 
    0.00011601822901301305, 0.00010928999798393325, 0.00010298622132142881, 
    9.7080777949313827e-05, 9.154827891282167e-05, 8.636418099867254e-05, 
    8.1504879759535157e-05, 7.6947781244361325e-05, 7.2671356469947333e-05, 
    6.8655185172024428e-05, 6.4879995557743191e-05, 6.1327704974891984e-05, 
    5.7981463274944224e-05, 5.4825696991097221e-05, 5.1846149112683306e-05, 
    4.9029906901243523e-05, 4.6365409321843531e-05, 4.3842426417106504e-05, 
    4.1452005208103028e-05, 3.9186380088285648e-05, 3.7038849642529909e-05, 
    3.5003625751132216e-05, 3.3075664137763445e-05, 3.1250487709610315e-05, 
    2.9524014823762942e-05, 2.7892403916184042e-05, 2.6351923894651388e-05, 
    2.4898856654265266e-05, 2.3529434488032505e-05, 2.223981154343705e-05, 
    2.1026065302273441e-05, 1.9884221706987324e-05, 1.8810296244249144e-05, 
    1.7800343066374932e-05, 1.6850504964437275e-05, 1.5957058452237794e-05, 
    1.5116450063534991e-05, 1.4325321877291519e-05, 1.3580525992384534e-05, 
    1.2879128978369068e-05, 1.2218408145984863e-05, 1.1595841813388926e-05, 
    1.1009095678319269e-05, 1.0456007066488882e-05, 9.9345683544611543e-06, 
    9.442910383521956e-06, 8.9792862823540578e-06, 8.5420558510071354e-06, 
    8.1296705421732491e-06, 7.7406590899207701e-06, 7.3736139470421466e-06, 
    7.0271788529215407e-06, 6.7000380181823466e-06, 6.3909075357808975e-06, 
    6.0985296756733271e-06, 5.8216706648367931e-06, 5.5591223862085018e-06, 
    5.3097081501875757e-06, 5.0722923258655581e-06, 4.8457932023371394e-06, 
    4.6291980404456378e-06, 4.4215789309882399e-06, 4.2221078600483731e-06, 
    4.0300693398454562e-06, 3.8448691213428615e-06, 3.6660378542338019e-06, 
    3.4932290645952239e-06, 3.326211412254759e-06, 3.1648557879001722e-06, 
    3.0091183247547154e-06, 2.8590207603657603e-06, 2.714629740631492e-06, 
    2.5760366010235933e-06, 2.4433389110083155e-06, 2.3166246860966892e-06, 
    2.195959730851687e-06, 2.0813781589384501e-06, 1.972875809630503e-06, 
    1.870406091460321e-06, 1.7738777441688582e-06, 1.6831541031782239e-06, 
    1.5980536293374071e-06, 1.5183516727985653e-06, 1.4437836097416038e-06, 
    1.3740495772540062e-06, 1.3088210042538446e-06, 1.2477489971251706e-06, 
    1.1904744101198494e-06, 1.1366391600305464e-06, 1.0858980860563117e-06, 
    1.0379304641864542e-06, 9.924502020239287e-07, 9.4921378846220395e-07, 
    9.0802525001162853e-07, 8.68737650995e-07, 8.3125102463573104e-07, 
    7.9550698869984349e-07, 7.6148062908657827e-07, 7.291704870912384e-07, 
    6.985876294644794e-07, 6.6974480635081535e-07, 6.4264661457361526e-07, 
    6.1728140688442659e-07, 5.9361545139337741e-07, 5.715895870928241e-07, 
    5.51118373755214e-07, 5.3209152634991886e-07, 5.1437727093209213e-07, 
    4.9782716861664867e-07, 4.8228192130372768e-07, 4.6757768703563349e-07, 
    4.5355247754943901e-07, 4.4005227126362265e-07, 4.2693653748307016e-07, 
    4.1408292533707362e-07, 4.0139092101822696e-07, 3.8878432248589915e-07, 
    3.7621242711180466e-07, 3.6364988184254213e-07, 3.5109521019432657e-07, 
    3.3856810725237385e-07, 3.261056771398554e-07, 3.1375786944126771e-07, 
    3.0158243962806142e-07, 2.8963980314099956e-07, 2.7798816305168603e-07, 
    2.6667926423872965e-07, 2.5575506204473079e-07, 2.4524549927679796e-07, 
    2.3516747235802796e-07, 2.2552495130101485e-07, 2.1631011252101237e-07, 
    2.0750526218311087e-07, 1.9908527795048623e-07, 1.9102028351626999e-07, 
    1.8327828973720882e-07, 1.7582758350776732e-07, 1.6863870986576287e-07, 
    1.6168596477750945e-07, 1.5494838363944858e-07, 1.4841026675842788e-07, 
    1.4206132099525917e-07, 1.3589651507504945e-07, 1.2991574452978524e-07, 
    1.2412338565582791e-07, 1.1852779045153493e-07, 1.1314074371018464e-07, 
    1.0797687457796056e-07, 1.0305299459829305e-07, 9.8387325015129101e-08, 
    9.3998580838477907e-08, 8.9904896316705397e-08, 8.6122604349711623e-08, 
    8.2664915084356291e-08, 7.9540572676980899e-08, 7.6752596191852767e-08, 
    7.4297226769717043e-08, 7.2163203803040866e-08, 7.0331476658918671e-08, 
    6.8775425165182091e-08, 6.7461616006827452e-08, 6.6351067562327652e-08, 
    6.5400940692210517e-08, 6.4566523804230932e-08, 6.3803345556908572e-08, 
    6.3069231738436161e-08, 6.2326128361906102e-08, 6.1541539274307389e-08, 
    6.0689471872560095e-08, 5.9750841068355634e-08, 5.8713343604314714e-08, 
    5.7570872008175806e-08, 5.6322583706487566e-08, 5.4971768804483117e-08, 
    5.3524668051477896e-08, 5.1989378861059639e-08, 5.0374957136534017e-08, 
    4.8690779435267879e-08, 4.6946183131848657e-08, 4.5150357120408091e-08, 
    4.3312420963488866e-08, 4.1441608654649572e-08, 3.9547469032147273e-08, 
    3.7640004939774968e-08, 3.5729697144069639e-08, 3.3827389043288986e-08, 
    3.1944041145205437e-08, 3.0090391830000818e-08, 2.8276581162306482e-08, 
    2.6511801669571451e-08, 2.4804036441753103e-08, 2.3159928982343258e-08, 
    2.158480695343335e-08, 2.0082854757870519e-08, 1.8657405052366756e-08, 
    1.7311298345834818e-08, 1.6047248369647171e-08, 1.4868148208357173e-08, 
    1.3777260652105318e-08, 1.2778251952743638e-08, 1.1875050909920013e-08, 
    1.1071539273772649e-08, 1.0371103671863278e-08, 9.7760981460314852e-09, 
    9.2872800516163753e-09, 8.903286692380458e-09, 8.6202177855240965e-09, 
    8.4313782872289081e-09, 8.3272207276870337e-09, 8.2955061040307817e-09, 
    8.3216819853977438e-09, 8.3894556407137664e-09, 8.4815227020219565e-09, 
    8.5803980333975041e-09, 8.6692873523615472e-09, 8.7329349270367526e-09, 
    8.758385707523059e-09, 8.7356076150176181e-09, 8.6579320697333608e-09, 
    8.5222852102678906e-09, 8.3291992332743116e-09, 8.082609323656965e-09, 
    7.7894574794080944e-09, 7.459136871091518e-09, 7.1028202173248601e-09, 
    6.7327208016758846e-09, 6.3613366558474833e-09, 6.0007257346417282e-09, 
    5.6618547300085829e-09, 5.354055884824982e-09, 5.084616799650723e-09, 
    4.8585176416914389e-09, 4.6783200445790802e-09, 4.5442021102014406e-09, 
    4.4541257334923495e-09, 4.4041152163775868e-09, 4.3886214556887003e-09, 
    4.4009423674640681e-09, 4.433669459219219e-09, 4.4791308051458073e-09, 
    4.5298037394426791e-09, 4.5786742359933023e-09, 4.6195259059298018e-09, 
    4.6471473402964526e-09, 4.6574536504733349e-09, 4.6475240707738132e-09, 
    4.6155639375695042e-09, 4.5608036648279079e-09, 4.4833513808277284e-09, 
    4.3840174472643486e-09, 4.2641297189612438e-09, 4.1253569823476193e-09, 
    3.9695556752110282e-09, 3.7986508802245908e-09, 3.6145584237228103e-09, 
    3.4191495657163187e-09, 3.2142551412015939e-09, 3.0017012368709927e-09, 
    2.7833652334566576e-09, 2.5612385343823148e-09, 2.3374818852847115e-09, 
    2.1144599757094891e-09, 1.8947449045680643e-09, 1.6810818246138029e-09, 
    1.476315255913111e-09, 1.283279459012293e-09, 1.1046614511199151e-09, 
    9.4284897279261538e-10, 7.9977846283853724e-10, 6.7679881613988277e-10, 
    5.7456585404618822e-10, 4.9297960107716438e-10, 4.3117268775694629e-10, 
    3.875529513293638e-10, 3.5989845460567154e-10, 3.4549769105478411e-10, 
    3.4132402633832959e-10, 3.4422988839610898e-10, 3.5114509639091014e-10, 
    3.5926324594939142e-10, 3.6620209454577229e-10, 3.7012617142077203e-10, 
    3.6982398871663394e-10, 3.6473621471713118e-10, 3.5493586449352269e-10, 
    3.4106508781307683e-10, 3.2423692488919384e-10, 3.0591206983238767e-10, 
    2.87762098681596e-10, 2.715301194230208e-10, 2.5889895900036694e-10, 
    2.5137465731019394e-10, 2.5019100957771741e-10, 2.5623805891538142e-10, 
    2.700154626102557e-10, 2.9160960443756685e-10, 3.2069235177984269e-10, 
    3.5653852877373644e-10, 3.9805930658207006e-10, 4.4384873979947058e-10, 
    4.9224129592464526e-10, 5.4137834326409357e-10, 5.8928187355592384e-10, 
    6.339334260997767e-10, 6.7335599321826928e-10, 7.0569600167208835e-10, 
    7.2930207243114552e-10, 7.4279675442974259e-10, 7.4513758180378742e-10, 
    7.3566383315486512e-10, 7.1412640863714273e-10, 6.8069900878225145e-10, 
    6.359703327656866e-10, 5.8091810891823424e-10, 5.1686729541184872e-10, 
    4.4543540656430728e-10, 3.6846888822020334e-10, 2.8797430125324709e-10, 
    2.0604821240678339e-10, 1.2480886371777241e-10, 4.6332268868286507e-11, 
    -2.7405560162848099e-11, -9.4579140072907433e-11, 
    -1.5355638524547754e-10, -2.0293350870637735e-10, 
    -2.4156219043784161e-10, -2.6856893851912493e-10, 
    -2.8336688319223901e-10, -2.8565995353374237e-10, 
    -2.7543971746815449e-10, -2.5297508066782736e-10, -2.187955416266235e-10, 
    -1.7366869418886269e-10, -1.1857327207468263e-10, 
    -5.4668898899083398e-11, 1.6735945677050682e-11, 9.4216619468711908e-11, 
    1.7626459862000395e-10, 2.6131873128768251e-10, 3.4779521458680841e-10, 
    4.3411641559398248e-10, 5.1873876823214247e-10, 6.0018024839988183e-10, 
    6.770475460516895e-10, 7.4806306418479149e-10, 8.1209126248577066e-10, 
    8.6816378776846818e-10, 9.1550220727367258e-10, 9.5353728118918926e-10, 
    9.8192336087905449e-10, 1.0005468944326794e-09, 1.0095280130445114e-09, 
    1.009214769066878e-09, 1.0001698076959954e-09, 9.8314985862781454e-10, 
    9.5907870659893545e-10, 9.2901474802849126e-10, 8.9411439165458461e-10, 
    8.5559290476950763e-10, 8.146841813358109e-10, 7.7260113266317505e-10, 
    7.3049814699493735e-10, 6.894370470026749e-10, 6.5035772426720392e-10, 
    6.1405437539203399e-10, 5.8115805223824464e-10, 5.521259605410384e-10, 
    5.2723752985122287e-10, 5.0659728615326606e-10, 4.901439587972466e-10, 
    4.7766539075794374e-10, 4.6881829115755673e-10, 4.6315203091488207e-10, 
    4.6013518476017049e-10, 4.5918386028488642e-10, 4.5969037580905808e-10, 
    4.6105123422262326e-10, 4.6269311678779678e-10, 4.6409595726597139e-10, 
    4.6481207214723228e-10, 4.6448086606706946e-10, 4.6283842779180647e-10, 
    4.5972199159607939e-10, 4.5506907898432762e-10, 4.4891167909005541e-10, 
    4.4136577640787318e-10, 4.3261694500177657e-10, 4.2290272132881926e-10, 
    4.1249284975243711e-10, 4.0166843663544994e-10, 3.9070139114670486e-10, 
    3.798353622099266e-10, 3.69269634073856e-10, 3.5914699627978748e-10, 
    3.4954666735052282e-10, 3.4048275968617619e-10, 3.3190847135739501e-10, 
    3.2372556534151741e-10, 3.1579829765073376e-10, 3.0797044024582698e-10, 
    3.0008376319760605e-10, 2.919961698883584e-10, 2.835978020013848e-10, 
    2.7482354332947087e-10, 2.6566093827609552e-10, 2.5615287903788953e-10, 
    2.4639513620721172e-10, 2.365291906728278e-10, 2.2673141720655203e-10, 
    2.1719973337190927e-10, 2.0813922940834883e-10, 1.9974798121029082e-10, 
    1.9220426745906214e-10, 1.8565599365881574e-10, 1.8021288761988929e-10, 
    1.7594172625046196e-10, 1.7286444757243545e-10, 1.7095888731963032e-10, 
    1.701617460961022e-10, 1.7037321695226756e-10, 1.7146281723305639e-10, 
    1.7327585617662233e-10, 1.7564018590125487e-10, 1.7837282393085365e-10, 
    1.812862173267379e-10, 1.8419389797434037e-10, 1.8691549293339742e-10, 
    1.8928097658502999e-10, 1.9113425972287187e-10, 1.923361325404728e-10, 
    1.9276670594595276e-10, 1.9232743986670819e-10, 1.9094287412609208e-10, 
    1.8856205104695627e-10, 1.8515968534290465e-10, 1.8073692565805339e-10, 
    1.7532163150659964e-10, 1.6896801833772853e-10, 1.6175548235330387e-10, 
    1.5378650680726454e-10, 1.4518364920737903e-10, 1.3608559352769033e-10, 
    1.2664248958832515e-10, 1.1701073024183317e-10, 1.0734752655485819e-10, 
    9.780557005201844e-11, 8.8528112646313189e-11, 7.9644728244720348e-11, 
    7.1268024412257266e-11, 6.349136313219018e-11, 5.6387696787254472e-11, 
    5.0009425461365507e-11, 4.4389193627009186e-11, 3.9541365423182577e-11, 
    3.5464068654033004e-11, 3.2141490592800051e-11, 2.9546313549208166e-11, 
    2.7642018532523271e-11, 2.6385106707633082e-11, 2.5727029441610845e-11, 
    2.5616000225599892e-11, 2.5998594140551276e-11, 2.6821286424577601e-11, 
    2.8031914721213838e-11, 2.9581098687750735e-11, 3.1423515900483187e-11, 
    3.3519012810138698e-11, 3.583328325368573e-11, 3.833814403886695e-11, 
    4.1011098915471199e-11, 4.3834351307329434e-11, 4.6793105746170424e-11, 
    4.9873517599057408e-11, 5.3060313341336579e-11, 5.6334615761187151e-11, 
    5.9672089666928466e-11, 6.3041887797940237e-11, 6.64064138719134e-11, 
    6.9722189747149217e-11, 7.2941569960427341e-11, 7.6015296236008366e-11, 
    7.8895387659342564e-11, 8.1538202684177104e-11, 8.3907064381881742e-11, 
    8.5974303835200346e-11, 8.772231946389524e-11, 8.9143665093950028e-11, 
    9.0240032835015818e-11, 9.1020499071006434e-11, 9.1499085195327757e-11, 
    9.1692208145352284e-11, 9.1616214185661607e-11, 9.1285497943838095e-11, 
    9.0711381568727622e-11, 8.9902037462686617e-11, 8.8863390019564058e-11, 
    8.7601023765819788e-11, 8.6122763321000795e-11, 8.4441699708771362e-11, 
    8.2579155507708672e-11, 8.0567291808750078e-11, 7.845081914872737e-11, 
    7.6287632330287304e-11, 7.4148033413559913e-11, 7.2112574629513963e-11, 
    7.0268536751573359e-11, 6.8705310876104554e-11, 6.7509034606949958e-11, 
    6.675692293738178e-11, 6.6511782135733494e-11, 6.6817166882909296e-11, 
    6.7693631902094415e-11, 6.9136373123905051e-11, 7.1114436147892167e-11, 
    7.3571605734126309e-11, 7.6428828662160882e-11, 7.9588064588603423e-11, 
    8.2937145909376697e-11, 8.6355456726315126e-11, 8.9719914041732739e-11, 
    9.2910993188988491e-11, 9.5818336405651965e-11, 9.8345758346856601e-11, 
    1.004153244478684e-10, 1.0197037529638877e-10, 1.0297732075044983e-10, 
    1.0342625324643318e-10, 1.0333028368544176e-10, 1.0272378980043071e-10, 
    1.0165963098977786e-10, 1.0020556774577628e-10, 9.8440102948125229e-11, 
    9.6448011194010853e-11, 9.4315796891929138e-11, 9.2127409320052793e-11, 
    8.9960389301770742e-11, 8.7882721537128178e-11, 8.5950440407502703e-11, 
    8.4206182616911629e-11, 8.267862916927107e-11, 8.1382838450033252e-11, 
    8.0321290243923124e-11, 7.9485615288472256e-11, 7.8858725237681929e-11, 
    7.8417213491785964e-11, 7.8133747980542164e-11, 7.7979376449903367e-11, 
    7.7925468595140764e-11, 7.7945258633090969e-11, 7.8014818929740501e-11, 
    7.8113548900118525e-11, 7.8224081691049392e-11, 7.8331837933724044e-11, 
    7.8424200802179654e-11, 7.84896011043333e-11, 7.851659321495968e-11, 
    7.8493128267976134e-11, 7.8406103753349893e-11, 7.8241319552586077e-11, 
    7.7983849306369272e-11, 7.7618810260384731e-11, 7.7132402598001228e-11, 
    7.6513178071061537e-11, 7.5753280183296687e-11, 7.4849620369648293e-11, 
    7.3804693599640423e-11, 7.2627071755664484e-11, 7.1331359617006585e-11, 
    6.9937702136060145e-11, 6.8470772415928387e-11, 6.6958425448598034e-11, 
    6.5430007370271062e-11, 6.3914607581703966e-11, 6.2439291153215774e-11, 
    6.1027546380970827e-11, 5.9698002972083096e-11, 5.8463584938802509e-11, 
    5.7331073728686268e-11, 5.6301142885653566e-11, 5.5368783922841311e-11, 
    5.4524095609684316e-11, 5.375323995998204e-11, 5.3039623672159418e-11, 
    5.2365017643891414e-11, 5.1710703169814907e-11, 5.1058434326534345e-11, 
    5.0391315981167434e-11, 4.9694473270645705e-11, 4.8955603238854269e-11, 
    4.8165365390820189e-11, 4.73176842817365e-11, 4.6409908973845793e-11, 
    4.5442930257432842e-11, 4.4421127081551127e-11, 4.3352260747213744e-11, 
    4.2247185804085607e-11, 4.11194413130627e-11, 3.9984686044243446e-11, 
    3.8860015350844357e-11, 3.7763128798126188e-11, 3.6711486039785765e-11, 
    3.5721419065229297e-11, 3.4807346910060969e-11, 3.3981056238916842e-11, 
    3.3251208075874997e-11, 3.2623034418740365e-11, 3.2098272429051729e-11, 
    3.1675303369915807e-11, 3.1349511768794698e-11, 3.1113774250053349e-11, 
    3.0959066759860783e-11, 3.0875078944836944e-11, 3.0850840206806225e-11, 
    3.087525938126163e-11, 3.0937589778847858e-11, 3.1027753538737612e-11, 
    3.1136592485834315e-11, 3.1255999932178042e-11, 3.1378996331438109e-11, 
    3.1499764378686264e-11, 3.1613667489053882e-11, 3.1717281244960849e-11, 
    3.1808441110395844e-11, 3.1886287036770086e-11, 3.1951317649339037e-11, 
    3.2005429870921464e-11, 3.2051882342597972e-11, 3.2095201642354905e-11, 
    3.2140966497722653e-11, 3.2195512277511984e-11, 3.2265513249099499e-11, 
    3.2357479831667431e-11, 3.2477243307211757e-11, 3.2629379178659689e-11, 
    3.2816750662620559e-11, 3.3040100889428199e-11, 3.3297835391639009e-11, 
    3.3585971112831033e-11, 3.3898343889835144e-11, 3.422693560084628e-11, 
    3.4562484386397972e-11, 3.4895193426040338e-11, 3.5215546647430003e-11, 
    3.5515111205053459e-11, 3.5787312038162384e-11, 3.6028011058863451e-11, 
    3.6235907778140181e-11, 3.6412638245436266e-11, 3.6562617244510052e-11, 
    3.669252646181773e-11, 3.6810598565350829e-11, 3.6925669403784354e-11, 
    3.7046132556417728e-11, 3.7178887536172849e-11, 3.7328416584732862e-11, 
    3.7496024686250593e-11, 3.7679416244597202e-11, 3.7872609455940087e-11, 
    3.8066225570745578e-11, 3.8248101669502468e-11, 3.8404238761998401e-11, 
    3.8519916802648087e-11, 3.8580927893790284e-11, 3.8574790685050932e-11, 
    3.849183412117984e-11, 3.8326022422757383e-11, 3.8075546041035571e-11, 
    3.7742990854163365e-11, 3.7335234925325216e-11, 3.6862985424872022e-11, 
    3.6340069219348202e-11, 3.578250895733624e-11, 3.5207491413859838e-11, 
    3.4632297299007945e-11, 3.4073281871037928e-11, 3.3544935497089704e-11, 
    3.3059139524504706e-11, 3.2624562302143735e-11, 3.2246331665099115e-11, 
    3.1925856718896291e-11, 3.1660905827923262e-11, 3.1445865289255337e-11, 
    3.1272185398436429e-11, 3.1128946488118193e-11, 3.1003587491692763e-11, 
    3.0882671598873973e-11, 3.0752750714975347e-11, 3.0601183906843496e-11, 
    3.0416949493368231e-11, 3.0191355075758734e-11, 2.9918610249562682e-11, 
    2.9596208252858846e-11, 2.9225134151346084e-11, 2.8809769535920067e-11, 
    2.8357613420014309e-11, 2.7878739245783446e-11, 2.73850895613966e-11, 
    2.6889582129220916e-11, 2.6405202114097127e-11, 2.5944074067474918e-11, 
    2.5516629877107029e-11, 2.5130919382181869e-11, 2.4792175729878476e-11, 
    2.4502555204816968e-11, 2.4261215848051942e-11, 2.4064564705257447e-11, 
    2.3906762295860539e-11, 2.378033405896779e-11, 2.3676884550074881e-11, 
    2.3587813155400719e-11, 2.3504982100909643e-11, 2.3421251169438652e-11, 
    2.3330884437166665e-11, 2.3229760389420377e-11, 2.3115414037914714e-11, 
    2.2986916414084249e-11, 2.2844628575123033e-11, 2.2689851732351192e-11, 
    2.2524470236606492e-11, 2.2350587944784708e-11, 2.2170252267572377e-11, 
    2.1985233579253685e-11, 2.1796975154092381e-11, 2.1606616081577649e-11, 
    2.1415162025308529e-11, 2.1223709238976357e-11, 2.1033738261275556e-11, 
    2.0847367082723951e-11, 2.066760274512523e-11, 2.0498457807693315e-11, 
    2.0344970686361754e-11, 2.0213079018761582e-11, 2.0109348488931575e-11, 
    2.004055013226156e-11, 2.0013172597723579e-11, 2.0032828995560333e-11, 
    2.010369158047547e-11, 2.0227917999644792e-11, 2.0405202624813118e-11, 
    2.0632451670674975e-11, 2.0903639876799045e-11, 2.1209836024919775e-11, 
    2.1539477273453544e-11, 2.1878792183856081e-11, 2.2212431094684089e-11, 
    2.2524188301481378e-11, 2.279784740594495e-11, 2.3017998406873919e-11, 
    2.3170853858072704e-11, 2.3244955788325273e-11, 2.3231765983443811e-11, 
    2.3126046879102869e-11, 2.2926106413206992e-11, 2.2633814526458275e-11, 
    2.2254477850974095e-11, 2.1796513976840541e-11, 2.1271051346001111e-11, 
    2.0691407568348102e-11, 2.0072523025609739e-11, 1.9430356851535036e-11, 
    1.8781305347704439e-11, 1.8141612752535506e-11, 1.752685484993447e-11, 
    1.6951431609196723e-11, 1.6428160545306843e-11, 1.5967916160224542e-11, 
    1.5579366620682186e-11, 1.5268777347105339e-11, 1.5039909264707557e-11, 
    1.4894003782148393e-11, 1.4829857650381045e-11, 1.4843943858906772e-11, 
    1.4930617274742817e-11, 1.5082355585268447e-11, 1.5290045235761677e-11, 
    1.5543245497510349e-11, 1.5830508333313815e-11, 1.6139666292118959e-11, 
    1.6458152362037612e-11, 1.6773288447567043e-11, 1.7072603821152e-11, 
    1.734416839276071e-11, 1.7576932822229848e-11, 1.7761067265329705e-11, 
    1.7888310682879261e-11, 1.795229542744606e-11, 1.7948850265345681e-11, 
    1.7876225010421703e-11, 1.7735250199515475e-11, 1.7529396806924013e-11, 
    1.7264731471024934e-11, 1.6949720701278473e-11, 1.6594951921836751e-11, 
    1.6212707010790487e-11, 1.5816465623843289e-11, 1.5420315607561482e-11, 
    1.503833905410447e-11, 1.4683977235642883e-11, 1.4369447613772215e-11, 
    1.410520337224844e-11, 1.3899519991727927e-11, 1.3758185074515952e-11, 
    1.3684344885805126e-11, 1.3678481654009914e-11, 1.3738535219778868e-11, 
    1.3860148910281091e-11, 1.4036998046784461e-11, 1.4261195232725492e-11, 
    1.4523720264096643e-11, 1.4814847441808117e-11, 1.512456281965363e-11, 
    1.5442908949431599e-11, 1.576030675908635e-11, 1.6067781210306542e-11, 
    1.6357135594367947e-11, 1.6621074531689163e-11, 1.6853282278745361e-11, 
    1.7048440579528973e-11, 1.7202252012636787e-11, 1.7311424319631957e-11, 
    1.7373662942964312e-11, 1.7387659190952173e-11, 1.735311718419075e-11, 
    1.7270720301201746e-11, 1.7142177705956775e-11, 1.6970213394005804e-11, 
    1.6758587784417263e-11, 1.6512058885028589e-11, 1.6236332839562255e-11, 
    1.5937965212447107e-11, 1.5624226409226137e-11, 1.5302868794952909e-11, 
    1.4981906489417738e-11, 1.4669307504986487e-11, 1.4372706317601025e-11, 
    1.4099071523864799e-11, 1.3854438715900685e-11, 1.3643627042910617e-11, 
    1.3470076636767153e-11, 1.3335685852890654e-11, 1.3240818446288116e-11, 
    1.3184269631749545e-11, 1.316342260913713e-11, 1.3174378414818809e-11, 
    1.3212218221389443e-11, 1.3271223958912248e-11, 1.3345189805429155e-11, 
    1.3427690382805907e-11, 1.3512391279152641e-11, 1.3593298161439823e-11, 
    1.3665032604272864e-11, 1.3723033162553154e-11, 1.3763774915383471e-11, 
    1.3784891897143294e-11, 1.378533252736178e-11, 1.3765395887551558e-11, 
    1.3726783015043598e-11, 1.3672540443432673e-11, 1.3606985375709022e-11, 
    1.3535510606358231e-11, 1.3464372409689786e-11, 1.3400336222430331e-11, 
    1.3350282381598325e-11, 1.3320763150587985e-11, 1.3317492152069459e-11, 
    1.3344821791664458e-11, 1.3405259324953726e-11, 1.3499038973991546e-11, 
    1.3623810803763134e-11, 1.3774453422148735e-11, 1.3943102726771227e-11, 
    1.4119328942304685e-11, 1.4290536864345691e-11, 1.4442558860269579e-11, 
    1.456037640865114e-11, 1.4628969290227399e-11, 1.4634216091026269e-11, 
    1.4563774780051826e-11, 1.4407922609760731e-11, 1.4160259442980927e-11, 
    1.3818250640490503e-11, 1.3383557950861032e-11, 1.2862150822612663e-11, 
    1.2264193203589439e-11, 1.1603703654393132e-11, 1.0898004963487819e-11, 
    1.0167015262627459e-11, 9.4323884552193908e-12, 8.7165785727915005e-12, 
    8.041845739003774e-12, 7.4292800978183209e-12, 6.8978463439557655e-12, 
    6.4635704213861868e-12, 6.1388109892333989e-12, 5.9317364114874835e-12, 
    5.8459622284343254e-12, 5.8804345452022987e-12, 6.029515392957287e-12, 
    6.2832983728144741e-12, 6.6281395043007279e-12, 7.0473819476792447e-12, 
    7.522218447789009e-12, 8.0326960550988504e-12, 8.5587471331958982e-12, 
    9.0812521658980252e-12, 9.5829981875945894e-12, 1.0049550417806844e-11, 
    1.0469871721666535e-11, 1.0836753692944332e-11, 1.1146930757448125e-11, 
    1.1400933210893038e-11, 1.1602622677492087e-11, 1.1758520795387125e-11, 
    1.1876922863640576e-11, 1.1966927887803576e-11, 1.2037426043085449e-11, 
    1.209620793587319e-11, 1.214920019971786e-11, 1.2199990957155342e-11, 
    1.2249597071718887e-11, 1.229657678431343e-11, 1.2337390667151781e-11, 
    1.2367032106728965e-11, 1.2379774042281355e-11, 1.237002089127616e-11, 
    1.2333066937469641e-11, 1.2265770779181276e-11, 1.2166994463042968e-11, 
    1.2037794831511492e-11, 1.1881350555802473e-11, 1.1702641946241211e-11, 
    1.1507923619976485e-11, 1.1304095335311564e-11, 1.1098002007622472e-11, 
    1.0895813623542678e-11, 1.0702507165944317e-11, 1.0521541580485749e-11, 
    1.035474105456564e-11, 1.0202380069876447e-11, 1.0063463409322971e-11, 
    9.936157095509183e-12, 9.8182223900222416e-12, 9.7075175701934623e-12, 
    9.6024042127653707e-12, 9.5020267978026753e-12, 9.4064515994774043e-12, 
    9.3166534481993735e-12, 9.2343471530350247e-12, 9.1617194037763617e-12, 
    9.1010764015889838e-12, 9.0545131447120894e-12, 9.023567069419985e-12, 
    9.0089917345746561e-12, 9.0105892763095463e-12, 9.0271879933844022e-12, 
    9.0566736464222513e-12, 9.0961585989074756e-12, 9.1421676313063509e-12, 
    9.1908879878524471e-12, 9.2384002206856699e-12, 9.2809235967514833e-12, 
    9.3150048121222189e-12, 9.3376905375231678e-12, 9.3466440477788877e-12, 
    9.3402420684295172e-12, 9.3176014915835066e-12, 9.2785927107952364e-12, 
    9.2238166322544227e-12, 9.1545272891177425e-12, 9.0725256892606235e-12, 
    8.9800217123915151e-12, 8.8794450706026849e-12, 8.7732533870501288e-12, 
    8.6637215803939473e-12, 8.5527389838802386e-12, 8.4416436300927798e-12, 
    8.3311209543197677e-12, 8.2211321075173149e-12, 8.1109630703271963e-12, 
    7.9993250982005086e-12, 7.8845431717472779e-12, 7.7647868175540681e-12, 
    7.6383237030932571e-12, 7.5037932249915954e-12, 7.3604218449674401e-12, 
    7.2082157324360897e-12, 7.0480626783746502e-12, 6.8817433874671552e-12, 
    6.7119045351762613e-12, 6.5419287315867474e-12, 6.3757544956981131e-12, 
    6.217712840626976e-12, 6.0722984698177823e-12, 5.9439971930800289e-12, 
    5.8371144329428024e-12, 5.7556476463163106e-12, 5.7031693910942959e-12, 
    5.6827637171124896e-12, 5.6969637423089495e-12, 5.7476790413798772e-12, 
    5.8361490625696631e-12, 5.9628797733680514e-12, 6.1275629311810929e-12, 
    6.3290118032772158e-12, 6.5651218483419363e-12, 6.8328123220929484e-12, 
    7.1280351605846787e-12, 7.4458373244870311e-12, 7.7804598011144207e-12, 
    8.1254819987518068e-12, 8.4740302293044784e-12, 8.8190031536675618e-12, 
    9.1533295409937381e-12, 9.4701869924819868e-12, 9.7632233970295314e-12, 
    1.0026726476021888e-11, 1.0255730157995223e-11, 1.0446080284400546e-11, 
    1.0594419428462166e-11, 1.0698156179194498e-11, 1.0755387731380329e-11, 
    1.0764828891556981e-11, 1.072574711782465e-11, 1.0637936663358719e-11, 
    1.0501733611781601e-11, 1.0318066059421026e-11, 1.0088570943319132e-11, 
    9.8156885560308403e-12, 9.5027967723033452e-12, 9.1543114807169672e-12, 
    8.7757226859088882e-12, 8.3735649983704079e-12, 7.9553021557984229e-12, 
    7.529102210927383e-12, 7.1035148945372604e-12, 6.6871148308215608e-12, 
    6.288064998146446e-12, 5.9136952663145715e-12, 5.5700969242214269e-12, 
    5.261836741481431e-12, 4.9917265115830297e-12, 4.7607761696318923e-12, 
    4.568248850422471e-12, 4.4118803989167454e-12, 4.2881620536486542e-12, 
    4.1927551587120096e-12, 4.120869486699324e-12, 4.0676686835666793e-12, 
    4.0285761774908161e-12, 3.9995350156198329e-12, 3.9771212051292228e-12, 
    3.9585751472325759e-12, 3.9417139431644618e-12, 3.92482511512978e-12, 
    3.906484491186132e-12, 3.885404088871471e-12, 3.8602911668787102e-12, 
    3.829798117853688e-12, 3.7924878034213463e-12, 3.7469091558871528e-12, 
    3.6916792274682753e-12, 3.6256303211332998e-12, 3.5479373459127015e-12, 
    3.4582666018889497e-12, 3.3568707457489294e-12, 3.244683271339343e-12, 
    3.1233493685274757e-12, 2.9952525945361716e-12, 2.863508137257241e-12, 
    2.7319307372155699e-12, 2.6049911453815296e-12, 2.4877724188725815e-12, 
    2.385881480577445e-12, 2.3053422104838054e-12, 2.2524344250191278e-12, 
    2.2335135466778369e-12, 2.2547446473198036e-12, 2.321803813533701e-12, 
    2.4395303860725177e-12, 2.611585306777806e-12, 2.8400734319112612e-12, 
    3.1252509695659129e-12, 3.4652727529677259e-12, 3.8560438584073022e-12, 
    4.2911976617078235e-12, 4.762212495532177e-12, 5.2586647338729399e-12, 
    5.7686036985037514e-12, 6.2790510391604594e-12, 6.7765706863251245e-12, 
    7.2478792209692583e-12, 7.6804628135645214e-12, 8.0631537972668634e-12, 
    8.3866154281393829e-12, 8.643720657891254e-12, 8.8297959525497813e-12, 
    8.9426959123057599e-12, 8.9827282213803528e-12, 8.9524458292905046e-12, 
    8.8562894977100257e-12, 8.7001349323078895e-12, 8.4908120055464332e-12, 
    8.2355852839096857e-12, 7.9416542456416118e-12, 7.6157573777679074e-12, 
    7.2638540547347054e-12, 6.8909355420843044e-12, 6.5010001472853216e-12, 
    6.0971345550246073e-12, 5.6817415868133683e-12, 5.256844131390675e-12, 
    4.8244447225668445e-12, 4.3868991005289486e-12, 3.9472411417447887e-12, 
    3.5094358733836124e-12, 3.0785069741734679e-12, 2.660547709603961e-12, 
    2.2625617347222033e-12, 1.8922033965753074e-12, 1.5573801706533408e-12, 
    1.2658007208790368e-12, 1.0244741409472703e-12, 8.3923204575776093e-13, 
    7.1430254254614035e-13, 6.5199461380614168e-13, 6.5246115449094478e-13, 
    7.1366843220270591e-13, 8.3142726055015512e-13, 9.9966288390798965e-13, 
    1.2106841350395765e-12, 1.4556769311568559e-12, 1.725125369262991e-12, 
    2.0093856745636478e-12, 2.2991316049284728e-12, 2.5858826472076497e-12, 
    2.8623202922911012e-12, 3.1226550393466891e-12, 3.3627491541744484e-12, 
    3.5802358702497079e-12, 3.7744288296539712e-12, 3.9462069634563224e-12, 
    4.0977115296268658e-12, 4.2320889217955978e-12, 4.3530601544983614e-12, 
    4.4646006952236142e-12, 4.5705282016892616e-12, 4.6742065476225619e-12, 
    4.7782603340832688e-12, 4.8844230406580314e-12, 4.9933899605045192e-12, 
    5.1048577401062276e-12, 5.2175717440357674e-12, 5.3295116036127082e-12, 
    5.4380803553956389e-12, 5.5403998112944339e-12, 5.6335639572909225e-12, 
    5.7149558126410098e-12, 5.7824741683298071e-12, 5.8347799267151023e-12, 
    5.8714277674521038e-12, 5.8929589615351368e-12, 5.9008744401508285e-12, 
    5.897575194878376e-12, 5.8861453996371138e-12, 5.8701396114662917e-12, 
    5.8532746832326972e-12, 5.8391286112865745e-12, 5.8308098307099896e-12, 
    5.8306941552035946e-12, 5.840183719769113e-12, 5.8595701286464088e-12, 
    5.8879648813745534e-12, 5.9233717860718774e-12, 5.9627839451794434e-12, 
    6.0024371395504882e-12, 6.0380846222572398e-12, 6.0653549235791778e-12, 
    6.0800810416436024e-12, 6.0786833764980774e-12, 6.058457050882743e-12, 
    6.0178502492262464e-12, 5.9566203847598454e-12, 5.8759327155088016e-12, 
    5.7782990624136719e-12, 5.6674635160714902e-12, 5.5481312700544124e-12, 
    5.4256473376168499e-12, 5.3055721966316022e-12, 5.1932681465912169e-12, 
    5.0934183349913621e-12, 5.0096560899157322e-12, 4.9442173621111498e-12, 
    4.8977467483665828e-12, 4.869194921623249e-12, 4.8559068333217825e-12, 
    4.8538280441147354e-12, 4.8578723479806917e-12, 4.8623471897022082e-12, 
    4.8614937551650913e-12, 4.849997080631148e-12, 4.8234879539550976e-12, 
    4.7789205832328429e-12, 4.714858336726844e-12, 4.6315791260209241e-12, 
    4.5310282941997168e-12, 4.4165996855198385e-12, 4.2927809755338303e-12, 
    4.1647224661765378e-12, 4.0377422006608512e-12, 3.9168423546554903e-12, 
    3.8062901115394902e-12, 3.7093147493985835e-12, 3.6279207815750699e-12, 
    3.5628659106975163e-12, 3.5137968481153466e-12, 3.4794671242549698e-12, 
    3.458083374172021e-12, 3.4476579516287811e-12, 3.4463782967935074e-12, 
    3.452884023107227e-12, 3.4664849270285159e-12, 3.487233023880239e-12, 
    3.5158942678227113e-12, 3.5538002818686386e-12, 3.6025833132724632e-12, 
    3.6639084889358626e-12, 3.7391591501344838e-12, 3.829130132256206e-12, 
    3.9338129182913668e-12, 4.052210708552048e-12, 4.1822937141032683e-12, 
    4.3209935310109957e-12, 4.4643454434105494e-12, 4.6076284184705789e-12, 
    4.7456107646110688e-12, 4.8727922145642526e-12, 4.9836826264702537e-12, 
    5.0730312518187474e-12, 5.1360758024666349e-12, 5.168735267493475e-12, 
    5.1677886299570048e-12, 5.1309887958722636e-12, 5.0571638034201479e-12, 
    4.946254760393628e-12, 4.7993405130103356e-12, 4.6185777292473485e-12, 
    4.4071407382501027e-12, 4.1690902964565232e-12, 3.9092323910495815e-12, 
    3.6329057485125868e-12, 3.3457899501521301e-12, 3.0536579241996359e-12, 
    2.7621606247809983e-12, 2.4766087823471616e-12, 2.2017979143807221e-12, 
    1.9418535550770531e-12, 1.7001439768990735e-12, 1.4792344746680844e-12, 
    1.2809012346622523e-12, 1.1061805606610163e-12, 9.55469971292509e-13, 
    8.2863472690135428e-13, 7.2514141568007838e-13, 6.4418292348014929e-13, 
    5.8479795016322329e-13, 5.4598006178325426e-13, 5.2676267581155102e-13, 
    5.2630070474300808e-13, 5.4393162256291247e-13, 5.7921593217502088e-13, 
    6.3198493703535211e-13, 7.0235385590130352e-13, 7.9072202958503603e-13, 
    8.9776088017311879e-13, 1.0243544417348623e-12, 1.1715042889625814e-12, 
    1.3402240496693938e-12, 1.531371485918135e-12, 1.7454966112321315e-12, 
    1.9826540291304405e-12, 2.2422507327505463e-12, 2.522916572982481e-12, 
    2.8224248520168654e-12, 3.1376752916682194e-12, 3.4647479242788162e-12, 
    3.7990076226928695e-12, 4.135277436284073e-12, 4.4680391219796396e-12, 
    4.7916779207868772e-12, 5.1006859454611362e-12, 5.3898774643870956e-12, 
    5.6545553523224815e-12, 5.8906401359109385e-12, 6.0947290450486613e-12, 
    6.2641403203532921e-12, 6.3968970021276473e-12, 6.4917017359780932e-12, 
    6.5479043360912178e-12, 6.565480070411233e-12, 6.54500035150093e-12, 
    6.4876502390889876e-12, 6.3952517453209552e-12, 6.2702839857392783e-12, 
    6.115932075522866e-12, 5.9360847913710023e-12, 5.7353217413591607e-12, 
    5.51884736263112e-12, 5.2923641164272252e-12, 5.0619197419902362e-12, 
    4.8336625579398503e-12, 4.6136180767092762e-12, 4.407395240883399e-12, 
    4.2199248739843471e-12, 4.0552571904751128e-12, 3.9163793684580531e-12, 
    3.8051008379453258e-12, 3.722031147531508e-12, 3.6666490427046295e-12, 
    3.6374237252384641e-12, 3.6319879625189938e-12, 3.6473692768949795e-12, 
    3.6802235803527095e-12, 3.7270416061672603e-12, 3.7843689457607185e-12, 
    3.8489591235840632e-12, 3.9178763611142166e-12, 3.9885660321765398e-12, 
    4.058883007267763e-12, 4.1270876420536614e-12, 4.1917986691571791e-12, 
    4.2519565992377612e-12, 4.3067707164837518e-12, 4.3556705191353315e-12, 
    4.3982351672202457e-12, 4.4341601916376639e-12, 4.463191090115402e-12, 
    4.4850852715325174e-12, 4.499558725657348e-12, 4.5062512303132582e-12, 
    4.5047009886687034e-12, 4.4943341034646418e-12, 4.4744814802374223e-12, 
    4.4444378547257434e-12, 4.4035041904504963e-12, 4.3511050284878737e-12, 
    4.2868658895461398e-12, 4.2107392323258769e-12, 4.1230766764434236e-12, 
    4.0246934270890513e-12, 3.9168740172249121e-12, 3.8013645848012139e-12, 
    3.6802608899954573e-12, 3.5559022581833789e-12, 3.4307069957419673e-12, 
    3.3070226430592629e-12, 3.1869373452055479e-12, 3.0721741883912554e-12, 
    2.9639848275116976e-12, 2.8631503935715467e-12, 2.7700006898679238e-12, 
    2.6845218955329931e-12, 2.6064991064377861e-12, 2.5356970544544396e-12, 
    2.4720052841912087e-12, 2.4155860364998558e-12, 2.3669435175123026e-12, 
    2.3269293619064003e-12, 2.296637786146046e-12, 2.2772507456730665e-12, 
    2.2697662837864916e-12, 2.2747356114293564e-12, 2.291958113550901e-12, 
    2.3202430177966591e-12, 2.3572207928314755e-12, 2.3993002425109667e-12, 
    2.4417282324242139e-12, 2.4788149911824486e-12, 2.5042578514884663e-12, 
    2.5115962495559096e-12, 2.4946907938481457e-12, 2.4482434558147724e-12, 
    2.3682350725114716e-12, 2.2523334012893895e-12, 2.1000952817380978e-12, 
    1.9130924736077424e-12, 1.6948451343735412e-12, 1.4506385220399965e-12, 
    1.1871723429649311e-12, 9.1216911309643058e-13, 6.3389634314770434e-13, 
    3.6070235978176371e-13, 1.0053676876704814e-13, -1.3942645880628273e-13, 
    -3.5314649004260927e-13, -5.3593381569434706e-13, 
    -6.8462214561523058e-13, -7.9760301130368648e-13, 
    -8.7481940565158921e-13, -9.1763064619263988e-13, 
    -9.2867205374210864e-13, -9.116062238718111e-13, -8.708886512205401e-13, 
    -8.1144641154273947e-13, -7.3842107443721831e-13, 
    -6.5683550470969316e-13, -5.7134056527310219e-13, 
    -4.8593929740045542e-13, -4.0379050736622948e-13, -3.270291338372155e-13, 
    -2.5669440269658628e-13, -1.9268517447045954e-13, 
    -1.3382584806346002e-13, -7.797701624169636e-14, -2.2236944599920366e-14, 
    3.6817129076243476e-14, 1.028487410580455e-13, 1.7947323886743746e-13, 
    2.699519000010095e-13, 3.7694193109717082e-13, 5.0228993823508077e-13, 
    6.4688082549275644e-13, 8.1058805927762127e-13, 9.9227672365347943e-13, 
    1.1899116897047042e-12, 1.4007256987821342e-12, 1.6214083909094803e-12, 
    1.8483581712694713e-12, 2.0779148889393443e-12, 2.306567714696109e-12, 
    2.5311199559064462e-12, 2.7488002296468154e-12, 2.9572907224700966e-12, 
    3.1547071079182118e-12, 3.3395007922883778e-12, 3.510327676845036e-12, 
    3.6659121285735003e-12, 3.8048995467890886e-12, 3.9257359431587917e-12, 
    4.0266228766002755e-12, 4.1055007061338882e-12, 4.1601342759241675e-12, 
    4.1882432053744301e-12, 4.187712806753454e-12, 4.1568084409366808e-12, 
    4.0944491960751614e-12, 4.0004274877615045e-12, 3.8756217474301766e-12, 
    3.7221378061031737e-12, 3.5433761015967502e-12, 3.3439902789232622e-12, 
    3.1297850262598907e-12, 2.9074724742837728e-12, 2.6843993922976631e-12, 
    2.4681716743616598e-12, 2.2662812949458589e-12, 2.0856867532379863e-12, 
    1.932452603626461e-12, 1.8114148075430727e-12, 1.7259338705250457e-12, 
    1.6777464654302728e-12, 1.6669212085193183e-12, 1.6919137467243793e-12, 
    1.7497366933948347e-12, 1.836222416129075e-12, 1.9463573332265098e-12, 
    2.0746214972167795e-12, 2.2153899114463511e-12, 2.3632766059846203e-12, 
    2.513460821487664e-12, 2.6619196605822462e-12, 2.8055907084564661e-12, 
    2.9424259255940797e-12, 3.0713556880357637e-12, 3.1921613856511499e-12, 
    3.3052765322024068e-12, 3.4115508439278913e-12, 3.511988814143933e-12, 
    3.6075071637223607e-12, 3.6987339163348471e-12, 3.7858823662309818e-12, 
    3.8687148703191303e-12, 3.9465660480287171e-12, 4.0184730558325669e-12, 
    4.0833641535866847e-12, 4.1402500506163484e-12, 4.1884558494733567e-12, 
    4.227812285488874e-12, 4.258728652004507e-12, 4.2822578736713896e-12, 
    4.3000163301749716e-12, 4.314028373437656e-12, 4.3265003077809701e-12, 
    4.3395584044404542e-12, 4.3549591482444042e-12, 4.3738471944601521e-12, 
    4.396553659421054e-12, 4.4225036552253051e-12, 4.4502121803144484e-12, 
    4.477393512498509e-12, 4.5011637070382766e-12, 4.5183240645585108e-12, 
    4.5256601467123044e-12, 4.520285589546321e-12, 4.4999175221343069e-12, 
    4.4631164473233187e-12, 4.4094301130376401e-12, 4.3394506256141986e-12, 
    4.2547366310909046e-12, 4.1576721935096166e-12, 4.0512472330334046e-12, 
    3.9387549393135187e-12, 3.8235265143679887e-12, 3.7086286046028151e-12, 
    3.5966191532549581e-12, 3.4893668274703631e-12, 3.3879598742238214e-12, 
    3.2926800425129977e-12, 3.2030811409482829e-12, 3.1181221633446618e-12, 
    3.0363622422808982e-12, 2.9561651197850216e-12, 2.8759404391147989e-12, 
    2.7943176228397055e-12, 2.7103155041982077e-12, 2.6234203586552944e-12, 
    2.5336459206735286e-12, 2.4414883165894103e-12, 2.3478558464334384e-12, 
    2.2539389319985152e-12, 2.1610921743043674e-12, 2.0706656086725598e-12, 
    1.9838915462540488e-12, 1.9017662933652027e-12, 1.8249872175170805e-12, 
    1.7539178409851008e-12, 1.6886190732125037e-12, 1.6288842435684743e-12, 
    1.5743529355066397e-12, 1.5245816181888404e-12, 1.4791981293935324e-12, 
    1.4379966597890604e-12, 1.4010403450918595e-12, 1.3687245433487361e-12, 
    1.3418147529230291e-12, 1.3214038340715062e-12, 1.308871999241309e-12, 
    1.3057422446099622e-12, 1.3135340424400204e-12, 1.3335664804502055e-12, 
    1.3667595293895174e-12, 1.4134384717080879e-12, 1.4731682164382378e-12, 
    1.5446251773501279e-12, 1.6255605636308649e-12, 1.7128095942613142e-12, 
    1.8023947801607165e-12, 1.8897027816913224e-12, 1.9697194402473753e-12, 
    2.037316196924737e-12, 2.0875516695128587e-12, 2.1159585016972798e-12, 
    2.1188218888350206e-12, 2.0933696601891694e-12, 2.0379325517470857e-12, 
    1.951988357845144e-12, 1.8361597265220034e-12, 1.6921256398249112e-12, 
    1.5224855481770421e-12, 1.3305903905220762e-12, 1.1203674502514439e-12, 
    8.9612992518598487e-13, 6.6243535487507941e-13, 4.2393547570694273e-13, 
    1.8528339696762634e-13, -4.8958737007415924e-14, -2.7439045996248909e-13, 
    -4.8683353569987473e-13, -6.8241982587051948e-13, 
    -8.5765827963053093e-13, -1.0095329391707961e-12, 
    -1.1356044577723733e-12, -1.2340926833631496e-12, 
    -1.3039505862620302e-12, -1.3449114250845612e-12, 
    -1.3575050165513019e-12, -1.3429930317903762e-12, 
    -1.3032864939442681e-12, -1.2408242766739151e-12, 
    -1.1584063434311518e-12, -1.059007232001001e-12, -9.4560720617359732e-13, 
    -8.2100723097967791e-13, -6.876951197271589e-13, -5.4773571943102824e-13, 
    -4.0269219264183973e-13, -2.5362140271964508e-13, 
    -1.0108265207614212e-13, 5.4805980667828488e-14, 2.142907121292563e-13, 
    3.7784395108386554e-13, 5.4604176401204837e-13, 7.1942572814776034e-13, 
    8.9836017632324202e-13, 1.0828904120471728e-12, 1.2726245192646728e-12, 
    1.4666400937908376e-12, 1.6634318430418348e-12, 1.8608913523099456e-12, 
    2.0563383396859265e-12, 2.2466050738070022e-12, 2.4281642020901828e-12, 
    2.5972966104650787e-12, 2.7502996727149422e-12, 2.8837107489421661e-12, 
    2.9945301743973115e-12, 3.0804355157151202e-12, 3.1399617147419552e-12, 
    3.1726311754874496e-12, 3.1790225927410832e-12, 3.1607679348219645e-12, 
    3.1204685341660194e-12, 3.061543522783504e-12, 2.9879989779008634e-12, 
    2.9041527483198325e-12, 2.8143209203190784e-12, 2.7224887772131772e-12, 
    2.6319880891583583e-12, 2.545248183774137e-12, 2.4635805271310457e-12, 
    2.3870753136165227e-12, 2.3146027510368441e-12, 2.2439279996804617e-12, 
    2.1719458760815006e-12, 2.0950113340850837e-12, 2.0093520585359406e-12, 
    1.9115177817946318e-12, 1.7988254293424206e-12, 1.6697739312822143e-12, 
    1.5243413475874018e-12, 1.3641921829278746e-12, 1.1926937902565903e-12, 
    1.0147911221293703e-12, 8.3670661111607609e-13, 6.6551173206876608e-13, 
    5.0858313623396749e-13, 3.7302775362975682e-13, 2.650727001396569e-13, 
    1.8957103171661439e-13, 1.4960197337587117e-13, 1.4618174946577233e-13, 
    1.7820892576275387e-13, 2.4257318370821883e-13, 3.3442775603435439e-13, 
    4.4759967967776482e-13, 5.7510140912607604e-13, 7.0967376113571593e-13, 
    8.443156785956887e-13, 9.7274673578090887e-13, 1.0897635297254765e-12, 
    1.1914468173163099e-12, 1.2752334872649828e-12, 1.3398506821832988e-12, 
    1.3851078782075169e-12, 1.4116382781406532e-12, 1.420578080000235e-12, 
    1.4132484554179181e-12, 1.3909062207485974e-12, 1.3545453721094069e-12, 
    1.3048102898555242e-12, 1.2420183712150472e-12, 1.166291613086091e-12, 
    1.0777244859293142e-12, 9.7662706250671112e-13, 8.6378483387774767e-13, 
    7.406806006709625e-13, 6.0963133508899375e-13, 4.7388251325481234e-13, 
    3.3757546508883365e-13, 2.0562814029613948e-13, 8.3504157567192089e-14, 
    -2.3066929521444503e-14, -1.0845506538661507e-13, 
    -1.6747780185122607e-13, -1.957589570893613e-13, -1.90036747844483e-13, 
    -1.484122911520089e-13, -7.0487504796477218e-14, 4.2560021206832097e-14, 
    1.8804185875536487e-13, 3.6189467506106011e-13, 5.5893537159081216e-13, 
    7.731324741422155e-13, 9.9797805327308769e-13, 1.2268325784733785e-12, 
    1.4532851084533452e-12, 1.6714634310496098e-12, 1.8763053521863032e-12, 
    2.0637346876161385e-12, 2.2307809928835456e-12, 2.37559214979482e-12, 
    2.4973985112352079e-12, 2.5963651858324469e-12, 2.6734583767910085e-12, 
    2.7301823583962885e-12, 2.7683631938454636e-12, 2.7899161421105416e-12, 
    2.7966068606266883e-12, 2.7898470047404535e-12, 2.7705315976372931e-12, 
    2.7389261547749458e-12, 2.6946139271247081e-12, 2.6365158567608325e-12, 
    2.562976891054979e-12, 2.4719336560056326e-12, 2.3611505263453626e-12, 
    2.2285220899635889e-12, 2.0724115051872473e-12, 1.8920140949201793e-12, 
    1.687701392176016e-12, 1.4613324411659578e-12, 1.2164571111969391e-12, 
    9.5844203502864572e-13, 6.9442203555880445e-13, 4.3311097814374431e-13, 
    1.8443342863271432e-13, -4.0932243027520948e-14, -2.3217866616915031e-13, 
    -3.7902403400317731e-13, -4.7239402092291094e-13, 
    -5.0504305742097946e-13, -4.7207890844913268e-13, 
    -3.7133158591647591e-13, -2.0354591144261909e-13, 2.7643019516919023e-14, 
    3.1590546720458415e-13, 6.5262364678314548e-13, 1.0274003297173056e-12, 
    1.4286663049442695e-12, 1.8443231971866935e-12, 2.2623708551798238e-12, 
    2.6714540028456513e-12, 3.0613129191309638e-12, 3.4231169733735245e-12, 
    3.7496682594825383e-12, 4.0354819526556141e-12, 4.276770051866379e-12, 
    4.471348169481444e-12, 4.618509133032762e-12, 4.7188568213659106e-12, 
    4.7741781666787334e-12, 4.7873134627421637e-12, 4.7620529680512515e-12, 
    4.7030607381610768e-12, 4.6157991892496458e-12, 4.5064400190402791e-12, 
    4.381740965148432e-12, 4.2488810684896622e-12, 4.115209542964635e-12, 
    3.9879539057096913e-12, 3.8738580060372022e-12, 3.7787839113111565e-12, 
    3.707299405751076e-12, 3.6622945040819836e-12, 3.6446767364282069e-12, 
    3.6531607271711445e-12, 3.6842014716380779e-12, 3.7320779672995079e-12, 
    3.7891669494186111e-12, 3.8463754008710089e-12, 3.8936776064912165e-12, 
    3.9207853112122422e-12, 3.917853229430924e-12, 3.876158992582218e-12, 
    3.7887352827795003e-12, 3.6508631042944849e-12, 3.4603987323309715e-12, 
    3.2179240404513853e-12, 2.9266795780004175e-12, 2.5923084351268408e-12, 
    2.2224743955039959e-12, 1.8263284217322758e-12, 1.4139117001200243e-12, 
    9.9555864852732031e-13, 5.8132696045710801e-13, 1.8050557309937652e-13, 
    -1.9877587047324931e-13, -5.4981138461368487e-13, 
    -8.6747173067912959e-13, -1.1482386757609155e-12, -1.390154387735838e-12, 
    -1.592688237650132e-12, -1.756557346177347e-12, -1.8835218694438718e-12, 
    -1.976148736829324e-12, -2.0375888352828932e-12, -2.0713242539090412e-12, 
    -2.0809394977316554e-12, -2.0698896683241876e-12, 
    -2.0412949306603712e-12, -1.9977361525540802e-12, 
    -1.9411242662755893e-12, -1.8725951367259956e-12, 
    -1.7924948945803607e-12, -1.7004377924238674e-12, 
    -1.5954578520349464e-12, -1.4762331005199996e-12, -1.341395983189077e-12, 
    -1.1898429409886859e-12, -1.0211087073110016e-12, 
    -8.3562877524548286e-13, -6.3498071442105295e-13, 
    -4.2201072807366649e-13, -2.0081448672071235e-13, 2.3436951296185061e-14, 
    2.4476880473235621e-13, 4.5683569591708087e-13, 6.5338027441574305e-13, 
    8.2876548256133101e-13, 9.7842837538546008e-13, 1.0993118352702797e-12, 
    1.1900977802956841e-12, 1.2513696662882691e-12, 1.2855159966191277e-12, 
    1.2965335851159905e-12, 1.2896239103687564e-12, 1.2707542760625346e-12, 
    1.2460868677630756e-12, 1.2214966325218706e-12, 1.2020760442162435e-12, 
    1.191813642978958e-12, 1.1933586214525052e-12, 1.2080101467147049e-12, 
    1.2357936978729544e-12, 1.2757469589016088e-12, 1.3262222853624392e-12, 
    1.3853056578624547e-12, 1.4511635427412874e-12, 1.5223867336320092e-12, 
    1.5981865235598536e-12, 1.6785083775243851e-12, 1.7639617915813377e-12, 
    1.855680669768615e-12, 1.9550103577500979e-12, 2.0632080003136684e-12, 
    2.1810559454224157e-12, 2.3085375597067229e-12, 2.4445604980249065e-12, 
    2.5868145409914443e-12, 2.7317323073612413e-12, 2.8745985647176291e-12, 
    3.00979107842073e-12, 3.1311405835162047e-12, 3.232362126821672e-12, 
    3.3075302520830741e-12, 3.3515534881715052e-12, 3.3605874422889743e-12, 
    3.3323694821111691e-12, 3.2664263805066183e-12, 3.1641327847595294e-12, 
    3.0286408203735299e-12, 2.8646554954804425e-12, 2.6780936794349374e-12, 
    2.4756536790017988e-12, 2.2643465618788958e-12, 2.0510038480952121e-12, 
    1.8418252460642764e-12, 1.6419812232984593e-12, 1.4553378102877978e-12, 
    1.2842623442382054e-12, 1.1295814165160997e-12, 9.9064805476087024e-13, 
    8.6553703069561872e-13, 7.5132109384773878e-13, 6.4443987973483611e-13, 
    5.4109620690827968e-13, 4.3767325528396796e-13, 3.3112407964433731e-13, 
    2.1931570975973422e-13, 1.0128336647820412e-13, -2.2620517937370907e-14, 
    -1.5068999678666551e-13, -2.7997337927909224e-13, 
    -4.0646524249024327e-13, -5.2545327611906311e-13, -6.318880019320021e-13, 
    -7.2083215118604159e-13, -7.878906335562216e-13, -8.296085573656531e-13, 
    -8.4377155225592361e-13,
  // Sqw-total(2, 0-1999)
    0.084250805145234489, 0.084016349327142748, 0.083319196383707786, 
    0.082177664994932037, 0.080621229019015583, 0.078689018365431823, 
    0.076427884437272192, 0.073890173800329167, 0.071131368436441259, 
    0.068207750661243585, 0.065174236575843911, 0.062082496334050295, 
    0.058979446158292259, 0.055906160047665104, 0.05289721254321756, 
    0.049980431241567924, 0.047177011559403084, 0.04450192804008489, 
    0.041964566657883666, 0.039569500562539696, 0.037317336254330188, 
    0.035205566601782798, 0.033229379582959635, 0.031382385414719348, 
    0.029657238365566156, 0.028046141919893519, 0.026541236354277933, 
    0.025134875838794545, 0.023819807824195932, 0.022589270875165872, 
    0.021437028558411522, 0.020357356863593128, 0.019345001317186947, 
    0.018395117820402682, 0.017503208639349673, 0.016665062185248519, 
    0.015876702475967796, 0.015134351644078453, 0.014434406675261377, 
    0.013773429800580373, 0.013148150660191751, 0.012555477500911598, 
    0.011992514232047884, 0.011456580086967009, 0.010945228851559921, 
    0.01045626504832298, 0.0099877550302501193, 0.0095380315730818205, 
    0.0091056911994867977, 0.0086895840792796941, 0.008288796893595669, 
    0.0079026295073397756, 0.0075305666514056254, 0.0071722460685374502, 
    0.0068274247226221803, 0.0064959447116540066, 0.0061777004631209196, 
    0.0058726086340281525, 0.0055805818977372563, 0.0053015074935646419, 
    0.0050352310658657307, 0.0047815459551994993, 0.0045401877555022122, 
    0.0043108336472106618, 0.0040931057810522833, 0.0038865778363585666, 
    0.0036907838161746474, 0.0035052281630879277, 0.0033293963691348495, 
    0.0031627653887677499, 0.0030048133219702697, 0.002855027993521967, 
    0.0027129141976558867, 0.0025779994954360846, 0.0024498385425888621, 
    0.0023280159913044319, 0.0022121480568472666, 0.0021018828753682274, 
    0.0019968998081264433, 0.0018969078716127873, 0.0018016434921225306, 
    0.0017108677945020089, 0.0016243636349446838, 0.0015419325747322208, 
    0.0014633919657033557, 0.0013885722814509635, 0.0013173147852679663, 
    0.0012494695821684918, 0.0011848940631041559, 0.0011234517186086111, 
    0.0010650112783114479, 0.0010094461217433715, 0.00095663390266419396, 
    0.0009064563310819464, 0.00085879906162940778, 0.00081355164231072721, 
    0.00077060748324854055, 0.00072986381138285888, 0.00069122158501975974, 
    0.00065458535247897999, 0.00061986305187146807, 0.00058696576323158595, 
    0.00055580743780366524, 0.00052630463963603685, 0.00049837633923481431, 
    0.00047194379614971051, 0.00044693055663975675, 0.00042326257527610067, 
    0.00040086844825504791, 0.00037967972511382598, 0.00035963124850941141, 
    0.00034066146221668677, 0.0003227126276906608, 0.00030573089982461411, 
    0.00028966623145138112, 0.00027447210063250862, 0.00026010508080445786, 
    0.00024652429712233197, 0.00023369082912027091, 0.00022156712755179146, 
    0.00021011651101411627, 0.00019930279639645768, 0.00018909009845108322, 
    0.00017944281098924154, 0.00017032575886535766, 0.00016170448936270271, 
    0.00015354565646358094, 0.00014581744339382924, 0.00013848996823370677, 
    0.00013153562366598244, 0.00012492931359557458, 0.00011864856439234942, 
    0.00011267350464049093, 0.0001069867224193137, 0.00010157302155987468, 
    9.6419106847544836e-05, 9.1513232217080528e-05, 8.6844845674697381e-05, 
    8.240426055960405e-05, 7.8182375799142745e-05, 7.4170459208943226e-05, 
    7.0359998895406326e-05, 6.6742619575308016e-05, 6.3310054051778761e-05, 
    6.0054155762633306e-05, 5.6966936476715439e-05, 5.404061372375887e-05, 
    5.1267654983928506e-05, 4.8640809400038064e-05, 4.6153122088957085e-05, 
    4.3797930312456609e-05, 4.1568844242431537e-05, 3.9459717424889274e-05, 
    3.746461314581522e-05, 3.5577772775403342e-05, 3.3793591047092372e-05, 
    3.2106601456546433e-05, 3.0511472938407881e-05, 2.9003017060239113e-05, 
    2.7576203458095516e-05, 2.6226180302536094e-05, 2.4948296288039451e-05, 
    2.3738120925374598e-05, 2.2591460648398005e-05, 2.1504369232537824e-05, 
    2.0473152063211217e-05, 1.949436470699696e-05, 1.85648068980149e-05, 
    1.7681513382810177e-05, 1.6841743068557708e-05, 1.6042967640960052e-05, 
    1.5282860360227242e-05, 1.4559285221688306e-05, 1.3870286205069389e-05, 
    1.3214076027989279e-05, 1.2589023728753465e-05, 1.1993640540729997e-05, 
    1.1426563852604197e-05, 1.0886539496462895e-05, 1.037240307036492e-05, 
    9.8830613755355675e-06, 9.417475245302699e-06, 8.9746450083533426e-06, 
    8.553599560445507e-06, 8.1533895572336996e-06, 7.7730846733984078e-06, 
    7.4117743040316425e-06, 7.0685706255840021e-06, 6.7426126704421699e-06, 
    6.4330700537337719e-06, 6.139145221480104e-06, 5.8600735201146591e-06, 
    5.5951209311912556e-06, 5.3435798674441001e-06, 5.104763880246208e-06, 
    4.8780024022478958e-06, 4.6626366943077588e-06, 4.4580179823081351e-06, 
    4.2635083960605378e-06, 4.0784848346516706e-06, 3.902345369676961e-06, 
    3.7345173519961831e-06, 3.5744660808388087e-06, 3.4217027730531733e-06, 
    3.2757906435699059e-06, 3.1363481551865783e-06, 3.0030488661872213e-06, 
    2.8756177368473044e-06, 2.7538241825795391e-06, 2.6374725269465058e-06, 
    2.526390769310269e-06, 2.4204187206926937e-06, 2.319396575347589e-06, 
    2.2231548920324981e-06, 2.1315067823920832e-06, 2.0442428757741094e-06, 
    1.961129377323655e-06, 1.8819092836318242e-06, 1.8063065826730491e-06, 
    1.7340330543381066e-06, 1.6647971086720533e-06, 1.5983139573213479e-06, 
    1.5343163129646964e-06, 1.4725647589422415e-06, 1.4128569324344689e-06, 
    1.355034727169201e-06, 1.2989888471460197e-06, 1.2446602304555168e-06, 
    1.1920381006850619e-06, 1.1411546772947872e-06, 1.0920768598264046e-06, 
    1.0448954684881498e-06, 9.9971284528047383e-07, 9.5662977301264195e-07, 
    9.1573273490047736e-07, 8.7708250972539606e-07, 8.4070497706172044e-07, 
    8.0658481015018751e-07, 7.7466247892213546e-07, 7.448347019041067e-07, 
    7.1695819857803133e-07, 6.9085633245088254e-07, 6.6632801935985451e-07, 
    6.4315812397299095e-07, 6.2112848709833096e-07, 6.0002872199224391e-07, 
    5.7966598326855888e-07, 5.5987304028070763e-07, 5.4051416208707898e-07, 
    5.2148852879420086e-07, 5.0273110301910348e-07, 4.8421110799683275e-07, 
    4.6592844452738316e-07, 4.4790852330869193e-07, 4.3019607796428278e-07, 
    4.1284855312060382e-07, 3.9592962958543535e-07, 3.7950336428731766e-07, 
    3.6362929781497219e-07, 3.483587369198205e-07, 3.3373227092327633e-07, 
    3.1977845010702855e-07, 3.0651345400233749e-07, 2.9394151888985253e-07, 
    2.8205587680522281e-07, 2.7083998062831786e-07, 2.602688391351303e-07, 
    2.5031035074790253e-07, 2.4092658932084019e-07, 2.3207504907309138e-07, 
    2.2370988808858231e-07, 2.1578321903027187e-07, 2.0824648104063232e-07, 
    2.0105189585761716e-07, 1.941539703989683e-07, 1.8751096899963298e-07, 
    1.8108624811907132e-07, 1.7484933326352635e-07, 1.6877662371047695e-07, 
    1.6285163746902947e-07, 1.5706475130906817e-07, 1.5141244487862153e-07, 
    1.4589611405437162e-07, 1.4052057097237036e-07, 1.3529238669247642e-07, 
    1.3021825396273847e-07, 1.2530354617428708e-07, 1.2055122602938509e-07, 
    1.1596121424666625e-07, 1.1153027169579657e-07, 1.0725238327773447e-07, 
    1.0311956890378265e-07, 9.9122992632534947e-08, 9.5254205083404598e-08, 
    9.1506339239636723e-08, 8.7875090653264585e-08, 8.4359345637406933e-08, 
    8.0961373149902183e-08, 7.768655805697866e-08, 7.4542718111118908e-08, 
    7.1539103032896e-08, 6.8685215383156328e-08, 6.5989611792913143e-08, 
    6.3458839235215436e-08, 6.1096634017494291e-08, 5.890346770741664e-08, 
    5.687646982588223e-08, 5.5009702401568942e-08, 5.3294713077635837e-08, 
    5.1721260310979789e-08, 5.0278088570935858e-08, 4.8953636898445477e-08, 
    4.7736586303891777e-08, 4.661618790431393e-08, 4.5582355663903658e-08, 
    4.4625549974285735e-08, 4.3736512530603911e-08, 4.2905935715817912e-08, 
    4.2124156536231271e-08, 4.1380957253733465e-08, 4.0665533090413787e-08, 
    3.9966657320859657e-08, 3.9273039321536909e-08, 3.857383896176397e-08, 
    3.7859274460675746e-08, 3.7121245545622732e-08, 3.6353889729799845e-08, 
    3.5553998081551969e-08, 3.4721234868379943e-08, 3.385813084055069e-08, 
    3.2969847520518314e-08, 3.2063736944223305e-08, 3.114874314606445e-08, 
    3.0234706826663934e-08, 2.933164077876978e-08, 2.8449041985268389e-08, 
    2.759529667981101e-08, 2.6777220341164588e-08, 2.5999757007978279e-08, 
    2.5265844620399051e-08, 2.457643693386929e-08, 2.3930660064207627e-08, 
    2.3326073086354238e-08, 2.2758998361329596e-08, 2.2224887146002969e-08, 
    2.1718689587785488e-08, 2.1235203476716489e-08, 2.0769382979490426e-08, 
    2.0316594994018736e-08, 1.987281700265029e-08, 1.9434774821178066e-08, 
    1.9000022288203359e-08, 1.8566966702206244e-08, 1.8134844973987575e-08, 
    1.7703655542799078e-08, 1.7274051368440038e-08, 1.6847199361555245e-08, 
    1.64246128290034e-08, 1.6007964596051972e-08, 1.5598890979425829e-08, 
    1.5198798722496149e-08, 1.4808689260464136e-08, 1.4429015575062488e-08, 
    1.4059586775243772e-08, 1.3699533120936842e-08, 1.3347340231806869e-08, 
    1.3000955104844022e-08, 1.2657959567641575e-08, 1.2315798939038036e-08, 
    1.1972046934899883e-08, 1.1624681978023973e-08, 1.1272347325049828e-08, 
    1.0914566826482571e-08, 1.055189157116536e-08, 1.018595806142445e-08, 
    9.8194473442712958e-09, 9.4559437975386834e-09, 9.0997026892760334e-09, 
    8.7553448214125168e-09, 8.4275043148353422e-09, 8.1204605009239778e-09, 
    7.8377870038080322e-09, 7.5820495129330356e-09, 7.3545796366170221e-09, 
    7.1553447970438617e-09, 6.9829256773415972e-09, 6.8346024749414405e-09, 
    6.7065419131942923e-09, 6.5940679255141737e-09, 6.4919922968410869e-09, 
    6.3949768808616789e-09, 6.2978976988645234e-09, 6.1961819678873744e-09, 
    6.0860931702800373e-09, 5.9649447278607919e-09, 5.8312301824614268e-09, 
    5.6846651788786322e-09, 5.5261443536010487e-09, 5.3576223401169365e-09, 
    5.1819334734731706e-09, 5.0025676929695055e-09, 4.8234216486310235e-09, 
    4.6485433058206904e-09, 4.4818865508511997e-09, 4.3270891868598356e-09, 
    4.1872843794389479e-09, 4.0649519925738247e-09, 3.9618132304722719e-09, 
    3.8787692534004754e-09, 3.8158826719193166e-09, 3.7723990766835161e-09, 
    3.7468051334804855e-09, 3.73691860810283e-09, 3.7400051812869005e-09, 
    3.7529159913680041e-09, 3.7722392948368304e-09, 3.7944588065312425e-09, 
    3.8161111669344616e-09, 3.8339348510598993e-09, 3.8450037570638596e-09, 
    3.8468395229381739e-09, 3.8374985825690761e-09, 3.8156314821633622e-09, 
    3.7805140480107777e-09, 3.732051375995814e-09, 3.6707569860997742e-09, 
    3.5977098764428531e-09, 3.514492735110988e-09, 3.4231141772006845e-09, 
    3.32591796116169e-09, 3.2254818241493073e-09, 3.1245089746449663e-09, 
    3.0257155591502244e-09, 2.9317183575250169e-09, 2.8449274269077858e-09, 
    2.7674493356707686e-09, 2.7010063961226724e-09, 2.6468771465489886e-09, 
    2.6058618357977838e-09, 2.5782751349818829e-09, 2.5639657569074781e-09, 
    2.5623605238724995e-09, 2.5725279194632771e-09, 2.5932548010799697e-09, 
    2.6231286812314293e-09, 2.6606183498073577e-09, 2.7041461565576075e-09, 
    2.7521472376494964e-09, 2.8031128994582885e-09, 2.8556178259523411e-09, 
    2.9083327993400245e-09, 2.9600264450014988e-09, 3.0095602954208706e-09, 
    3.0558819701201512e-09, 3.0980204646643838e-09, 3.135086670975368e-09, 
    3.1662805991261368e-09, 3.1909053389218946e-09, 3.2083861831014631e-09, 
    3.2182924482774373e-09, 3.2203587875177385e-09, 3.2145028301552362e-09, 
    3.200836343673345e-09, 3.1796679691774941e-09, 3.1514964730392025e-09, 
    3.1169946246366421e-09, 3.0769844993530716e-09, 3.0324060182399043e-09, 
    2.984280583884104e-09, 2.9336722634724318e-09, 2.8816485509935318e-09, 
    2.8292428357582214e-09, 2.7774201974707623e-09, 2.7270479185347693e-09, 
    2.678871695572237e-09, 2.6334982192589396e-09, 2.5913843938923671e-09, 
    2.552833252059269e-09, 2.5179961846905683e-09, 2.4868809832651844e-09, 
    2.459364807227582e-09, 2.4352111601444399e-09, 2.4140897275664563e-09, 
    2.3955980293457262e-09, 2.3792837676923097e-09, 2.364666997677351e-09, 
    2.3512612800578368e-09, 2.3385932056259855e-09, 2.3262198226393665e-09, 
    2.3137435887904841e-09, 2.300824536511048e-09, 2.2871894953447471e-09, 
    2.2726381063269787e-09, 2.2570454998858251e-09, 2.2403615128040271e-09, 
    2.2226064348009514e-09, 2.203863343608804e-09, 2.1842673372160046e-09, 
    2.1639921094947004e-09, 2.1432345519700572e-09, 2.1221982630258139e-09, 
    2.1010770363832735e-09, 2.0800394351385327e-09, 2.0592156540723559e-09, 
    2.038687650406442e-09, 2.0184834072219655e-09, 1.9985758101913944e-09, 
    1.9788862585896395e-09, 1.9592926541167598e-09, 1.9396410898084769e-09, 
    1.9197600984379766e-09, 1.8994762101096858e-09, 1.8786293356472645e-09, 
    1.8570866539568648e-09, 1.8347538423924874e-09, 1.8115827918329502e-09, 
    1.7875753430020017e-09, 1.7627830638417965e-09, 1.7373033460709492e-09, 
    1.7112725857399038e-09, 1.6848572290906321e-09, 1.658243764724451e-09, 
    1.6316284921090651e-09, 1.6052079648589682e-09, 1.5791706238287528e-09, 
    1.5536900559672202e-09, 1.5289199518777136e-09, 1.5049907284062086e-09, 
    1.4820075275302615e-09, 1.4600493974804463e-09, 1.4391692485647385e-09, 
    1.419394405004576e-09, 1.400727474186503e-09, 1.3831475311808108e-09, 
    1.366611527565829e-09, 1.3510560587218537e-09, 1.3363994838254184e-09, 
    1.322544569159253e-09, 1.3093816239282725e-09, 1.296792181472896e-09, 
    1.2846530825443358e-09, 1.2728408683015665e-09, 1.2612362294887793e-09, 
    1.2497283371256531e-09, 1.2382187399328611e-09, 1.2266246919465515e-09, 
    1.21488159013841e-09, 1.2029445322429396e-09, 1.1907888335859056e-09, 
    1.1784095439897436e-09, 1.1658199977846588e-09, 1.1530496325663953e-09, 
    1.1401411254648347e-09, 1.1271471956509839e-09, 1.114127210971889e-09, 
    1.1011438804654327e-09, 1.0882601646225574e-09, 1.0755366213042025e-09, 
    1.0630291985294889e-09, 1.05078759742627e-09, 1.0388540888362688e-09, 
    1.0272628161141393e-09, 1.0160394336106226e-09, 1.0052010510482363e-09, 
    9.947563027438361e-10, 9.8470562486216033e-10, 9.7504160626200091e-10, 
    9.6574948420883667e-10, 9.5680777445850114e-10, 9.4818918026595602e-10, 
    9.3986168625142362e-10, 9.3179004156287083e-10, 9.2393748768085481e-10, 
    9.1626778666873725e-10, 9.0874740544072174e-10, 9.0134775619475075e-10, 
    8.9404726720867537e-10, 8.8683315499551908e-10, 8.7970261702602344e-10, 
    8.7266337783405789e-10, 8.6573336690499102e-10, 8.5893958864972305e-10, 
    8.5231614803326717e-10, 8.459016346843916e-10, 8.397360140516163e-10, 
    8.3385739247443471e-10, 8.2829883298304209e-10, 8.2308564079196724e-10, 
    8.1823321138329177e-10, 8.1374572025251308e-10, 8.0961559563530073e-10, 
    8.0582381100378432e-10, 8.0234076379985858e-10, 7.9912763867326665e-10, 
    7.9613791086990625e-10, 7.9331889915778142e-10, 7.9061312259288279e-10, 
    7.8795945415834919e-10, 7.8529401312717632e-10, 7.8255100056539662e-10, 
    7.796635143855077e-10, 7.7656464899753432e-10, 7.7318894044420884e-10, 
    7.6947438706598007e-10, 7.6536495916507687e-10, 7.608136665222496e-10, 
    7.5578587234369905e-10, 7.5026273176415737e-10, 7.4424430998491933e-10, 
    7.3775214229179548e-10, 7.308307741748865e-10, 7.2354814305529761e-10, 
    7.1599445110315412e-10, 7.0827961008711668e-10, 7.0052916389163005e-10, 
    6.9287899998779286e-10, 6.854690203915722e-10, 6.7843630388631801e-10, 
    6.7190805325071704e-10, 6.6599495835941222e-10, 6.6078528160026611e-10, 
    6.5634018181147457e-10, 6.5269045375428979e-10, 6.4983500887846882e-10, 
    6.4774102161170442e-10, 6.4634582105485198e-10, 6.4556023019654864e-10, 
    6.4527323684222741e-10, 6.4535752160453946e-10, 6.4567566198883283e-10, 
    6.4608649552688788e-10, 6.4645144494227179e-10, 6.4664037078760369e-10, 
    6.4653679677216779e-10, 6.460422361670288e-10, 6.4507952070962206e-10, 
    6.4359493978091825e-10, 6.415592950455953e-10, 6.3896767332841998e-10, 
    6.3583819738579048e-10, 6.3220966540116242e-10, 6.2813836422658553e-10, 
    6.2369413212433272e-10, 6.1895598124798174e-10, 6.1400746911717684e-10, 
    6.089321387751003e-10, 6.0380925375822312e-10, 5.9871015725338439e-10, 
    5.9369538634069976e-10, 5.888127877133331e-10, 5.8409667342357837e-10, 
    5.7956807625787484e-10, 5.7523589714046444e-10, 5.7109895823184834e-10, 
    5.671485348091671e-10, 5.6337120459056222e-10, 5.5975159959672531e-10, 
    5.5627486072134567e-10, 5.529284567718548e-10, 5.4970326583854291e-10, 
    5.4659377862790698e-10, 5.4359752621467482e-10, 5.4071377687843944e-10, 
    5.3794181961541824e-10, 5.3527898605584556e-10, 5.3271881303706576e-10, 
    5.3024955578442632e-10, 5.2785328395479603e-10, 5.2550573478013746e-10, 
    5.2317694817396985e-10, 5.2083265986158819e-10, 5.1843631959594809e-10, 
    5.1595150357691521e-10, 5.1334452100505534e-10, 5.1058690093868429e-10, 
    5.0765756961199192e-10, 5.0454446717463439e-10, 5.0124551885796922e-10, 
    4.9776885088491686e-10, 4.9413229796459021e-10, 4.9036226166786525e-10, 
    4.8649204553632938e-10, 4.8255983725164573e-10, 4.7860650894994791e-10, 
    4.7467340365502619e-10, 4.7080024468894289e-10, 4.6702329409087588e-10, 
    4.6337382265305632e-10, 4.5987692185316809e-10, 4.5655069175547378e-10, 
    4.5340574874696088e-10, 4.5044506495957203e-10, 4.4766404948217546e-10, 
    4.4505089962094154e-10, 4.4258715359321431e-10, 4.4024845914516423e-10, 
    4.3800550685520616e-10, 4.3582519183927601e-10, 4.3367190497415352e-10, 
    4.3150901057103191e-10, 4.2930041346803394e-10, 4.2701218606637221e-10, 
    4.2461417030633544e-10, 4.2208148161814439e-10, 4.1939577759425183e-10, 
    4.1654626955172705e-10, 4.1353031148373941e-10, 4.1035359101815128e-10, 
    4.0702984688353138e-10, 4.035801590864408e-10, 4.0003181715466563e-10, 
    3.9641689263313361e-10, 3.9277057750652384e-10, 3.8912944147407366e-10, 
    3.8552967468640731e-10, 3.8200548137100485e-10, 3.785876715456093e-10, 
    3.7530254501857119e-10, 3.7217106632399941e-10, 3.6920839218142e-10, 
    3.6642368877156959e-10, 3.6382025589706956e-10, 3.6139585508873307e-10, 
    3.5914325061574732e-10, 3.5705088119072651e-10, 3.5510364625013755e-10, 
    3.532837184466803e-10, 3.5157143663812888e-10, 3.4994617397325972e-10, 
    3.4838722731630105e-10, 3.4687466023772198e-10, 3.4539012456436851e-10, 
    3.4391758622887594e-10, 3.4244397399315166e-10, 3.4095964554130978e-10, 
    3.3945872840402259e-10, 3.3793920346632525e-10, 3.3640279854897467e-10, 
    3.3485460059574396e-10, 3.3330247390527768e-10, 3.3175626415019492e-10, 
    3.3022687450507643e-10, 3.2872525277375295e-10, 3.2726143226122846e-10, 
    3.2584360304054765e-10, 3.2447741994283632e-10, 3.2316549478817173e-10, 
    3.2190719294276402e-10, 3.2069868994161966e-10, 3.1953336509616898e-10, 
    3.1840235583988063e-10, 3.1729538862465922e-10, 3.1620168353701007e-10, 
    3.151109414518637e-10, 3.140142536172239e-10, 3.1290494465796679e-10, 
    3.1177917216010447e-10, 3.1063632830684991e-10, 3.0947910589227036e-10, 
    3.0831330009454396e-10, 3.0714724369409347e-10, 3.0599102646654683e-10, 
    3.0485545158906526e-10, 3.0375088483068918e-10, 3.0268603787349086e-10, 
    3.0166686368910805e-10, 3.0069555657366852e-10, 2.9976988909339383e-10, 
    2.9888286044918087e-10, 2.9802275817485551e-10, 2.9717357406352036e-10, 
    2.9631587374066151e-10, 2.9542791855136182e-10, 2.9448706054864803e-10, 
    2.9347124888634907e-10, 2.9236055020242809e-10, 2.9113852167709056e-10, 
    2.8979341194681132e-10, 2.8831897065692033e-10, 2.8671493891706995e-10, 
    2.8498707204380147e-10, 2.8314678459064036e-10, 2.8121036306441482e-10, 
    2.7919790550591649e-10, 2.7713197047765466e-10, 2.7503614444870506e-10, 
    2.7293352670081909e-10, 2.7084536179880698e-10, 2.6878978128727322e-10, 
    2.6678088614831539e-10, 2.6482809041197955e-10, 2.6293587482355571e-10, 
    2.6110388693826336e-10, 2.593274040578769e-10, 2.5759808487046617e-10, 
    2.5590499921212273e-10, 2.5423578164496447e-10, 2.5257790979880829e-10, 
    2.5091991479938759e-10, 2.492525467278264e-10, 2.4756969160040978e-10, 
    2.4586908198839111e-10, 2.4415265116737259e-10, 2.4242657883786653e-10, 
    2.4070094502283647e-10, 2.3898907939179897e-10, 2.3730657458462942e-10, 
    2.3567011246372938e-10, 2.3409610324329799e-10, 2.3259932059970023e-10, 
    2.3119161217044556e-10, 2.2988078927213603e-10, 2.2866980012134337e-10, 
    2.2755630256789972e-10, 2.2653257837489073e-10, 2.2558593210274503e-10, 
    2.2469942131417512e-10, 2.2385294210252649e-10, 2.230245064642438e-10, 
    2.2219166495848226e-10, 2.2133290227486923e-10, 2.2042894309958916e-10, 
    2.1946381884002097e-10, 2.1842571222919693e-10, 2.1730743253154183e-10, 
    2.1610662866892843e-10, 2.1482567362571909e-10, 2.1347130867174494e-10, 
    2.1205408006635734e-10, 2.1058765332265648e-10, 2.0908802851376102e-10, 
    2.0757275739881836e-10, 2.0606014648319117e-10, 2.0456853308589304e-10, 
    2.0311561262539576e-10, 2.0171786588025808e-10, 2.0039004454518594e-10, 
    1.9914478020848321e-10, 1.9799226227830973e-10, 1.9694003248924087e-10, 
    1.9599286147900536e-10, 1.9515274813337582e-10, 1.9441898916804615e-10, 
    1.9378836581938624e-10, 1.9325537234179171e-10, 1.9281250476364084e-10, 
    1.9245057567290527e-10, 1.921590074131188e-10, 1.919260869082355e-10, 
    1.9173917988469469e-10, 1.9158487532999993e-10, 1.9144907565336317e-10, 
    1.9131705782553338e-10, 1.9117353588373454e-10, 1.9100275876292963e-10, 
    1.9078870228891564e-10, 1.9051536028761759e-10, 1.9016718779960762e-10, 
    1.8972966392789693e-10, 1.8918996184679872e-10, 1.8853770652433897e-10, 
    1.8776571870349776e-10, 1.8687067988109374e-10, 1.858536699114697e-10, 
    1.8472047639394399e-10, 1.8348165379909536e-10, 1.8215226488125512e-10, 
    1.8075135260550624e-10, 1.7930112814088594e-10, 1.7782594980664803e-10, 
    1.7635115368115049e-10, 1.7490182536611911e-10, 1.7350157155790272e-10, 
    1.721714363630692e-10, 1.7092892070675097e-10, 1.6978728395306365e-10, 
    1.6875506827930569e-10, 1.6783590644340677e-10, 1.6702857615297348e-10, 
    1.6632731129458798e-10, 1.6572230744085032e-10, 1.6520040771546826e-10, 
    1.647458661877326e-10, 1.6434120684354918e-10, 1.6396807241559462e-10, 
    1.6360806203832302e-10, 1.6324346336251111e-10, 1.6285793013452674e-10, 
    1.6243700537527094e-10, 1.6196855285091891e-10, 1.6144301795304053e-10, 
    1.6085359373242678e-10, 1.6019624291813803e-10, 1.5946965180162304e-10, 
    1.5867504053899553e-10, 1.5781596227323909e-10, 1.5689798999870635e-10, 
    1.5592842618135204e-10, 1.5491593643315313e-10, 1.5387022375632614e-10, 
    1.5280168680077802e-10, 1.5172111385667605e-10, 1.5063937868106006e-10, 
    1.4956718678715562e-10, 1.4851482682410892e-10, 1.4749196421209505e-10, 
    1.4650743003685363e-10, 1.4556905369769271e-10, 1.4468346653958305e-10, 
    1.438559655225462e-10, 1.4309035132985589e-10, 1.4238882109683857e-10, 
    1.4175187819694926e-10, 1.4117830975027034e-10, 1.406651956437762e-10, 
    1.4020802772610129e-10, 1.3980085367353041e-10, 1.3943654952258836e-10, 
    1.3910711250395577e-10, 1.3880403171535286e-10, 1.3851867170299324e-10, 
    1.3824267383059859e-10, 1.3796830317871855e-10, 1.3768878579125462e-10, 
    1.3739850589589771e-10, 1.370931602659373e-10, 1.367697569226676e-10, 
    1.3642655300207259e-10, 1.3606284351250352e-10, 1.3567873366340555e-10, 
    1.3527481636855984e-10, 1.3485188117384384e-10, 1.3441062096683752e-10, 
    1.3395143516179869e-10, 1.3347424790017507e-10, 1.3297849313355239e-10, 
    1.3246312762557132e-10, 1.3192678856140387e-10, 1.3136795005715678e-10, 
    1.3078517209439372e-10, 1.3017732827541546e-10, 1.295438580329413e-10, 
    1.2888492250696492e-10, 1.2820157800038826e-10, 1.2749584221976621e-10, 
    1.26770741823199e-10, 1.2603026009699938e-10, 1.2527927842736016e-10, 
    1.2452342369472446e-10, 1.2376892657173953e-10, 1.2302239414795496e-10, 
    1.2229062570768209e-10, 1.2158030390387926e-10, 1.2089777455795347e-10, 
    1.202487453274689e-10, 1.1963804765317844e-10, 1.1906936507061455e-10, 
    1.1854505707873382e-10, 1.1806599286538901e-10, 1.1763150804067043e-10, 
    1.172394036773371e-10, 1.1688608557888796e-10, 1.1656676407631063e-10, 
    1.1627577290965317e-10, 1.1600693621512182e-10, 1.1575400432625624e-10, 
    1.1551106787671665e-10, 1.1527299238439025e-10, 1.150357408031438e-10, 
    1.1479662036741408e-10, 1.1455438820869536e-10, 1.1430920741112661e-10, 
    1.1406242110353122e-10, 1.1381618993430489e-10, 1.1357301272265847e-10, 
    1.1333515784793011e-10, 1.131040469759853e-10, 1.1287971393182461e-10, 
    1.1266032765347812e-10, 1.1244189778376188e-10, 1.1221814780389593e-10, 
    1.1198065839269825e-10, 1.1171917335596157e-10, 1.1142215985669601e-10, 
    1.1107751122250296e-10, 1.1067335539837294e-10, 1.1019889930481729e-10, 
    1.096452488197201e-10, 1.0900612490882257e-10, 1.0827841680060533e-10, 
    1.0746257203780259e-10, 1.065627484403875e-10, 1.0558673674046213e-10, 
    1.0454570622684133e-10, 1.0345374557121099e-10, 1.0232727988351728e-10, 
    1.0118437172806639e-10, 1.0004397882513035e-10, 9.8925204895985068e-11, 
    9.7846580532719391e-11, 9.6825412171902728e-11, 9.5877225345314214e-11, 
    9.5015302728335025e-11, 9.4250363194292997e-11, 9.3590325347086236e-11, 
    9.304020562988743e-11, 9.2602078495733755e-11, 9.2275143469866025e-11, 
    9.2055840709576486e-11, 9.1938010606256733e-11, 9.1913131898661438e-11, 
    9.1970569787015442e-11, 9.209787347147606e-11, 9.2281132138957565e-11, 
    9.2505366055893847e-11, 9.27549719325244e-11, 9.3014205299029631e-11, 
    9.326771505616971e-11, 9.350105808544904e-11, 9.3701221091789697e-11, 
    9.3857096189903443e-11, 9.3959873270738944e-11, 9.4003318094408968e-11, 
    9.3983936284939492e-11, 9.390097279382825e-11, 9.3756291576153688e-11, 
    9.3554081592844675e-11, 9.3300490660123037e-11, 9.3003148048077867e-11, 
    9.2670670425074508e-11, 9.2312133474307831e-11, 9.1936610122916366e-11, 
    9.1552738908067154e-11, 9.1168403177842496e-11, 9.079047805264778e-11, 
    9.0424707473770985e-11, 9.007561740359592e-11, 8.974655051997054e-11, 
    8.9439710147340698e-11, 8.9156266333248226e-11, 8.8896444575793394e-11, 
    8.8659643446264343e-11, 8.8444509002357031e-11, 8.8249024104337303e-11, 
    8.807056253009509e-11, 8.7905951636921451e-11, 8.7751531949142738e-11, 
    8.7603243324801338e-11, 8.7456716961858352e-11, 8.7307412438469714e-11, 
    8.7150773886344025e-11, 8.6982437573052554e-11, 8.6798399524770877e-11, 
    8.6595245994397414e-11, 8.6370325365115941e-11, 8.6121907261835045e-11, 
    8.584926672934082e-11, 8.5552726710493825e-11, 8.523360548270491e-11, 
    8.489410088127147e-11, 8.4537088903568169e-11, 8.416589868740454e-11, 
    8.3784011602609182e-11, 8.3394784167541948e-11, 8.3001170870326794e-11, 
    8.2605504418060987e-11, 8.2209312476954561e-11, 8.1813249540425937e-11, 
    8.1417077057679757e-11, 8.1019757488663607e-11, 8.0619599896176636e-11, 
    8.021446717371253e-11, 7.9802015238009271e-11, 7.9379933033833892e-11, 
    7.8946161245293079e-11, 7.8499090266169924e-11, 7.8037662153463191e-11, 
    7.7561453978283214e-11, 7.7070681367528648e-11, 7.6566155330652858e-11, 
    7.6049199770940559e-11, 7.5521564239478248e-11, 7.4985318805767068e-11, 
    7.4442788159211935e-11, 7.3896503110413272e-11, 7.3349182238353131e-11, 
    7.2803751529660972e-11, 7.2263395557072519e-11, 7.1731560385291685e-11, 
    7.12120013398568e-11, 7.0708737569387508e-11, 7.0225987116695736e-11, 
    6.9768008089641236e-11, 6.9338894641926727e-11, 6.8942305890752172e-11, 
    6.8581177820403804e-11, 6.8257420005869728e-11, 6.7971687157851791e-11, 
    6.772318817965385e-11, 6.7509657629163704e-11, 6.7327432446859335e-11, 
    6.7171697160580472e-11, 6.7036865587836822e-11, 6.6917062817714523e-11, 
    6.6806678379990729e-11, 6.6700924913059683e-11, 6.6596322252965768e-11, 
    6.6491074843299397e-11, 6.6385262529308203e-11, 6.628084100429625e-11, 
    6.6181405018919509e-11, 6.6091777082394969e-11, 6.6017426413672232e-11, 
    6.5963791150305511e-11, 6.5935594985524563e-11, 6.5936218360271648e-11, 
    6.5967180622974593e-11, 6.6027820497559025e-11, 6.6115200035900887e-11, 
    6.6224205430118521e-11, 6.6347868785823255e-11, 6.6477824645994374e-11, 
    6.6604885598729009e-11, 6.6719642156124205e-11, 6.6813007261508844e-11, 
    6.6876691877605829e-11, 6.6903547901056535e-11, 6.6887748423612175e-11, 
    6.6824837466936362e-11, 6.6711632547776948e-11, 6.6546067208554919e-11, 
    6.6326954939163385e-11, 6.6053783670510446e-11, 6.5726524659552693e-11, 
    6.5345539742579761e-11, 6.4911559152089111e-11, 6.4425757922596999e-11, 
    6.388991557592257e-11, 6.3306605144896488e-11, 6.2679409691172305e-11, 
    6.2013115920723362e-11, 6.1313828964491902e-11, 6.0588999365051017e-11, 
    5.9847331474863538e-11, 5.9098561207234578e-11, 5.8353116068438533e-11, 
    5.7621708204273882e-11, 5.6914845069306496e-11, 5.624234448101058e-11, 
    5.5612871054996142e-11, 5.5033573605158606e-11, 5.4509803948190955e-11, 
    5.4044993653119402e-11, 5.3640649775195195e-11, 5.3296485750236595e-11, 
    5.3010632440141437e-11, 5.2779941918844828e-11, 5.2600276872905847e-11, 
    5.246680151993416e-11, 5.2374198840238915e-11, 5.2316829484300372e-11, 
    5.2288799781647738e-11, 5.2283956571796846e-11, 5.2295834759513518e-11, 
    5.2317610715625597e-11, 5.2342070700136924e-11, 5.2361644915869502e-11, 
    5.236853961761136e-11, 5.2354975348287235e-11, 5.2313515046124849e-11, 
    5.2237475702892701e-11, 5.2121370093094098e-11, 5.1961330335147786e-11, 
    5.1755469379418486e-11, 5.1504124984292253e-11, 5.12099600748465e-11, 
    5.0877893457093765e-11, 5.0514866653545644e-11, 5.0129472803814581e-11, 
    4.9731503181990366e-11, 4.9331409819830756e-11, 4.8939808004750149e-11, 
    4.8567019118972746e-11, 4.8222700669808419e-11, 4.7915580145402036e-11, 
    4.765330257769782e-11, 4.7442358049224514e-11, 4.7288074896975468e-11, 
    4.719461478205218e-11, 4.7164950962453164e-11, 4.7200811652894832e-11, 
    4.7302544867787525e-11, 4.7468914368443485e-11, 4.7696886736052412e-11, 
    4.7981381699783871e-11, 4.8315099344127778e-11, 4.8688423221465812e-11, 
    4.9089483739789318e-11, 4.9504377505861777e-11, 4.9917590949344538e-11, 
    5.0312585809406167e-11, 5.067255023462906e-11, 5.0981220353061276e-11, 
    5.1223754709997348e-11, 5.1387539716364413e-11, 5.1462895410730762e-11, 
    5.1443583031237299e-11, 5.132709676012951e-11, 5.1114689541202882e-11, 
    5.0811155023987215e-11, 5.042436059892859e-11, 4.9964604382169078e-11, 
    4.9443836949003085e-11, 4.8874832479642131e-11, 4.827035872384705e-11, 
    4.7642443839824868e-11, 4.7001785512156077e-11, 4.6357334533951439e-11, 
    4.5716100537081989e-11, 4.508315162774951e-11, 4.4461819882021004e-11, 
    4.3854061860003308e-11, 4.3260919478986606e-11, 4.2683048295993292e-11, 
    4.2121229174066774e-11, 4.1576822842980519e-11, 4.1052114003132044e-11, 
    4.0550512225020989e-11, 4.0076588617296993e-11, 3.963595219502546e-11, 
    3.9234962490077053e-11, 3.8880341299897519e-11, 3.8578680309079537e-11, 
    3.8335918938269802e-11, 3.8156850345350928e-11, 3.8044684849553995e-11, 
    3.8000680624951454e-11, 3.8023977282922546e-11, 3.811149780499083e-11, 
    3.8258089322271674e-11, 3.8456731025093347e-11, 3.8698950925843957e-11, 
    3.8975260098554649e-11, 3.9275719957245319e-11, 3.9590449754833299e-11, 
    3.9910190576553916e-11, 4.0226700817938143e-11, 4.053315234042225e-11, 
    4.0824300476691826e-11, 4.1096591725248356e-11, 4.1348054263276272e-11, 
    4.1578132612274787e-11, 4.1787339159138636e-11, 4.1976919715026953e-11, 
    4.2148410883616242e-11, 4.2303306079952145e-11, 4.2442707122174418e-11, 
    4.2567134982575449e-11, 4.2676417994620122e-11, 4.2769755829653507e-11, 
    4.284582153484881e-11, 4.2903050568211189e-11, 4.2939889309335618e-11, 
    4.2955140081077496e-11, 4.2948208756694585e-11, 4.2919330991819591e-11, 
    4.2869658941023373e-11, 4.2801300278246799e-11, 4.2717157933408493e-11, 
    4.2620759663317409e-11, 4.2515950248558889e-11, 4.2406590761859376e-11, 
    4.2296208065093383e-11, 4.2187735060434956e-11, 4.208323494927844e-11, 
    4.198378000442913e-11, 4.1889376131986921e-11, 4.1799023986120923e-11, 
    4.1710823363800051e-11, 4.1622212769396604e-11, 4.1530200840642121e-11, 
    4.1431693487050673e-11, 4.1323767013212377e-11, 4.1203984972040905e-11, 
    4.1070609831473508e-11, 4.092281335618586e-11, 4.0760778457726434e-11, 
    4.0585753749243025e-11, 4.0399989135796313e-11, 4.0206642102682605e-11, 
    4.0009571970183749e-11, 3.981311262388622e-11, 3.962177080590107e-11, 
    3.9439944015270467e-11, 3.9271570539442216e-11, 3.9119854426179636e-11, 
    3.8986959280911733e-11, 3.8873799204226014e-11, 3.8779844709305806e-11, 
    3.8703057236649323e-11, 3.8639844911054648e-11, 3.8585182801696933e-11, 
    3.853279602782843e-11, 3.8475475137989415e-11, 3.8405457934610631e-11, 
    3.8314941930921647e-11, 3.8196589219019891e-11, 3.804413301316244e-11, 
    3.7852887969358048e-11, 3.7620253546220412e-11, 3.7346065040851215e-11, 
    3.7032813075281755e-11, 3.6685630974371188e-11, 3.6312110722039124e-11, 
    3.5921855346535532e-11, 3.5525899465449661e-11, 3.5135907181436171e-11, 
    3.4763353839548871e-11, 3.4418651039688009e-11, 3.4110393028736707e-11, 
    3.384471149253775e-11, 3.3624903312550061e-11, 3.3451277634350516e-11, 
    3.3321328301950707e-11, 3.3230141292549266e-11, 3.3171061798016045e-11, 
    3.3136462002168016e-11, 3.3118634497149647e-11, 3.3110609163643375e-11, 
    3.3106899294623571e-11, 3.3103998956585667e-11, 3.3100695296792605e-11, 
    3.3098061254525309e-11, 3.3099224501638233e-11, 3.3108881663256715e-11, 
    3.3132646544622613e-11, 3.3176306521297864e-11, 3.324506374810238e-11, 
    3.3342812478633178e-11, 3.3471564406168674e-11, 3.3631031766428738e-11, 
    3.3818438176065338e-11, 3.4028514164239974e-11, 3.4253740943398498e-11, 
    3.4484728533147744e-11, 3.4710768041759599e-11, 3.4920443410459141e-11, 
    3.5102312170435748e-11, 3.5245524979012511e-11, 3.5340429784531509e-11, 
    3.5379031533163504e-11, 3.5355373429013237e-11, 3.5265718741341044e-11, 
    3.5108631155659578e-11, 3.4884899320400091e-11, 3.4597357715126011e-11, 
    3.4250585998835912e-11, 3.3850586873623567e-11, 3.3404418225997434e-11, 
    3.2919843808796214e-11, 3.2404996768708295e-11, 3.1868125414533433e-11, 
    3.1317369345915592e-11, 3.0760622490114752e-11, 3.0205432553889629e-11, 
    2.9658968235930338e-11, 2.9127970691905187e-11, 2.8618760065625546e-11, 
    2.813719568958543e-11, 2.7688643170038674e-11, 2.7277910795800886e-11, 
    2.6909170424280711e-11, 2.6585858770510539e-11, 2.6310597352726347e-11, 
    2.6085102073501163e-11, 2.5910147490737576e-11, 2.578554660461349e-11, 
    2.5710203995174764e-11, 2.5682195233556717e-11, 2.5698917704908297e-11, 
    2.5757248713051958e-11, 2.5853757757413299e-11, 2.598490106166391e-11, 
    2.6147207410411527e-11, 2.63374504899386e-11, 2.6552762662909422e-11, 
    2.6790687159552533e-11, 2.7049197051689271e-11, 2.7326633641215828e-11, 
    2.7621617187601539e-11, 2.7932906805147111e-11, 2.8259251779753487e-11, 
    2.8599246716893456e-11, 2.8951190708111508e-11, 2.9312991262708467e-11, 
    2.9682111284011053e-11, 3.0055543558250001e-11, 3.0429852907581505e-11, 
    3.0801242473059958e-11, 3.1165661071883627e-11, 3.1518899981034322e-11, 
    3.1856712284353955e-11, 3.2174915180768766e-11, 3.2469467033764525e-11, 
    3.2736510328220462e-11, 3.297241303281105e-11, 3.3173749241247522e-11, 
    3.3337303491950669e-11, 3.3460045071165153e-11, 3.3539135131149182e-11, 
    3.357191960795518e-11, 3.355598252606394e-11, 3.348922167690909e-11, 
    3.3369954263608428e-11, 3.3197067492728827e-11, 3.2970197363967296e-11, 
    3.2689899844034707e-11, 3.2357847532779242e-11, 3.1976981733403933e-11, 
    3.1551645082049657e-11, 3.1087617300114659e-11, 3.0592133249219416e-11, 
    3.0073726411176068e-11, 2.9542038853371951e-11, 2.9007514059801444e-11, 
    2.8481010548917309e-11, 2.7973319696858654e-11, 2.7494679519102977e-11, 
    2.7054271438397107e-11, 2.6659752027471822e-11, 2.6316833642287961e-11, 
    2.6029012457262196e-11, 2.5797373256190786e-11, 2.5620577863698328e-11, 
    2.5495002367537141e-11, 2.5415023016153206e-11, 2.5373403678895471e-11, 
    2.5361820814970083e-11, 2.5371422712445894e-11, 2.5393431257891184e-11, 
    2.5419683814017467e-11, 2.5443135384146659e-11, 2.5458241028951671e-11, 
    2.5461216978096073e-11, 2.5450127775861932e-11, 2.5424856141796893e-11, 
    2.5386893837514705e-11, 2.5339054964664056e-11, 2.5285057553925194e-11, 
    2.5229093659089456e-11, 2.517536060808458e-11, 2.5127652412658678e-11, 
    2.5088999014387703e-11, 2.506142079086783e-11, 2.5045767010073818e-11, 
    2.5041718116045693e-11, 2.5047847277215945e-11, 2.5061833990962435e-11, 
    2.5080711892874165e-11, 2.5101175360303808e-11, 2.5119889638872093e-11, 
    2.5133792544733672e-11, 2.5140315448242373e-11, 2.5137564947978417e-11, 
    2.5124399132311584e-11, 2.5100454288624053e-11, 2.5066042473736686e-11, 
    2.5022040734879043e-11, 2.4969710644306466e-11, 2.4910528817519585e-11, 
    2.4846003246539892e-11, 2.477753489212925e-11, 2.4706315437615699e-11, 
    2.4633288134719153e-11, 2.4559104272206263e-11, 2.448416702136195e-11, 
    2.4408644598720228e-11, 2.4332509661584029e-11, 2.4255527366342281e-11, 
    2.4177244494153911e-11, 2.409692097425789e-11, 2.4013462328956118e-11, 
    2.3925317796906432e-11, 2.3830429448053251e-11, 2.3726182961961833e-11, 
    2.3609454071499522e-11, 2.347670255481236e-11, 2.3324175347628733e-11, 
    2.31481394781701e-11, 2.2945207998465327e-11, 2.2712640707467345e-11, 
    2.2448662749762634e-11, 2.2152690606554073e-11, 2.1825518764966702e-11, 
    2.1469349783865665e-11, 2.1087758280973557e-11, 2.0685528839481834e-11, 
    2.0268445105054841e-11, 1.9842969811276137e-11, 1.9415970347712369e-11, 
    1.8994423016968749e-11, 1.8585165215514223e-11, 1.8194694571154254e-11, 
    1.7829034203337121e-11, 1.749363027092447e-11, 1.7193302637604989e-11, 
    1.6932176581079274e-11, 1.6713656985485307e-11, 1.6540326003458341e-11, 
    1.6413878546210666e-11, 1.6334982363172091e-11, 1.6303190398431576e-11, 
    1.6316819198711082e-11, 1.6372936769655448e-11, 1.6467344811287721e-11, 
    1.6594731986694385e-11, 1.6748845974152977e-11, 1.692283283871704e-11, 
    1.7109594836480114e-11, 1.7302253990526617e-11, 1.7494564566164023e-11, 
    1.7681358176176073e-11, 1.7858862524146943e-11, 1.8024963824394864e-11, 
    1.8179278448351666e-11, 1.8323131305439726e-11, 1.8459361605398455e-11, 
    1.8592031848613864e-11, 1.8726016610295275e-11, 1.8866568518399297e-11, 
    1.9018857958600114e-11, 1.9187553757027234e-11, 1.9376458926767942e-11, 
    1.9588240307051045e-11, 1.982425177171731e-11, 2.0084463571826475e-11, 
    2.0367455380599194e-11, 2.0670504108316828e-11, 2.0989703974686791e-11, 
    2.1320122877426351e-11, 2.1655966425401325e-11, 2.1990765111403601e-11, 
    2.2317549332018783e-11, 2.2629046545956955e-11, 2.2917886342080973e-11, 
    2.317681509747341e-11, 2.3398952920715147e-11, 2.3578048573889975e-11, 
    2.3708734327817578e-11, 2.3786787112489435e-11, 2.3809325411498477e-11, 
    2.3774976441389684e-11, 2.3683958514537056e-11, 2.3538081710222354e-11, 
    2.3340661125825494e-11, 2.3096356444185129e-11, 2.2810951089079222e-11, 
    2.2491085498550306e-11, 2.2144001835917569e-11, 2.1777277222626537e-11, 
    2.1398597875045929e-11, 2.1015587762408846e-11, 2.0635658366160507e-11, 
    2.0265919435515974e-11, 1.991310602812411e-11, 1.958351463711618e-11, 
    1.9282934221002311e-11, 1.9016558283467803e-11, 1.8788874069374103e-11, 
    1.8603521096238909e-11, 1.8463154430623101e-11, 1.8369298776728552e-11, 
    1.8322243654859452e-11, 1.8320972213042948e-11, 1.8363189787534386e-11, 
    1.8445423512045575e-11, 1.8563190826176097e-11, 1.8711273152143344e-11, 
    1.8884044058806388e-11, 1.9075817676084531e-11, 1.9281212615688148e-11, 
    1.9495454646102427e-11, 1.9714623535166381e-11, 1.9935782493498344e-11, 
    2.0156999508025931e-11, 2.0377242317762394e-11, 2.0596168667605346e-11, 
    2.0813839072004218e-11, 2.1030379574629269e-11, 2.1245642278336145e-11, 
    2.1458932471283595e-11, 2.1668807033831678e-11, 2.1872984390056538e-11, 
    2.2068400182548901e-11, 2.2251397225044521e-11, 2.2417994326550977e-11, 
    2.2564286383103809e-11, 2.2686837472229836e-11, 2.278303757520077e-11, 
    2.2851431369009811e-11, 2.2891894233172404e-11, 2.2905670408899904e-11, 
    2.2895271621300609e-11, 2.2864206598370494e-11, 2.281660710909398e-11, 
    2.2756779869951911e-11, 2.268874253051191e-11, 2.2615803309010051e-11, 
    2.2540254449715935e-11, 2.2463182231857696e-11, 2.238446494603612e-11, 
    2.2302917455426449e-11, 2.2216578311604327e-11, 2.2123095913613733e-11, 
    2.2020141363264476e-11, 2.1905802940394628e-11, 2.1778905341113225e-11, 
    2.1639198605934234e-11, 2.1487379361823987e-11, 2.1324973639843153e-11, 
    2.115409921078156e-11, 2.0977096967003697e-11, 2.0796184062665564e-11, 
    2.0613095486381412e-11, 2.0428815295847765e-11, 2.0243434622272822e-11, 
    2.0056169376777426e-11, 1.9865501641193946e-11, 1.9669464684741784e-11, 
    1.9466003365759141e-11, 1.9253352577046111e-11, 1.9030392273772799e-11, 
    1.8796925908453855e-11, 1.8553826638816383e-11, 1.8303031176076595e-11, 
    1.804740427688383e-11, 1.7790472799278407e-11, 1.7536082743293614e-11, 
    1.7288009561734742e-11, 1.7049599907295591e-11, 1.6823482430449769e-11, 
    1.6611383350521718e-11, 1.6414061116685632e-11, 1.6231396302684692e-11, 
    1.606256442111315e-11, 1.5906317403621516e-11, 1.5761294650913678e-11, 
    1.5626336367819217e-11, 1.5500736651181348e-11, 1.5384416872641993e-11, 
    1.5277996398181435e-11, 1.5182738306036784e-11, 1.510037887635387e-11, 
    1.5032884579366674e-11, 1.4982129758263376e-11, 1.4949562913726384e-11, 
    1.4935895111397742e-11, 1.4940844184170669e-11, 1.4962946271166174e-11, 
    1.4999508788590249e-11, 1.5046647171605619e-11, 1.5099461483851791e-11, 
    1.5152306730158263e-11, 1.5199132069736114e-11, 1.5233899706647221e-11, 
    1.5250996070042923e-11, 1.5245628874489843e-11, 1.521417617903078e-11, 
    1.5154451521314834e-11, 1.506586224134708e-11, 1.4949449537433832e-11, 
    1.4807784634195814e-11, 1.4644774711783424e-11, 1.4465321885888053e-11, 
    1.4274937490899275e-11, 1.4079284535690065e-11, 1.3883725916421873e-11, 
    1.3692903954888046e-11, 1.3510404577748576e-11, 1.3338527993257886e-11, 
    1.3178221529838664e-11, 1.3029141487124604e-11, 1.2889891795335282e-11, 
    1.2758370176140075e-11, 1.2632215238760015e-11, 1.2509284718987339e-11, 
    1.2388119078225858e-11, 1.2268325524445405e-11, 1.2150844279885052e-11, 
    1.2038040532402532e-11, 1.1933645636062469e-11, 1.1842515357351181e-11, 
    1.1770260168178766e-11, 1.1722783986946914e-11, 1.1705782908836203e-11, 
    1.1724256800638733e-11, 1.178212678182887e-11, 1.1881932866454789e-11, 
    1.2024682287921296e-11, 1.2209841582151201e-11, 1.2435451240133744e-11, 
    1.2698334935683853e-11, 1.2994377240406263e-11, 1.3318808022281851e-11, 
    1.3666477157353668e-11, 1.4032080738265234e-11, 1.4410318407770967e-11, 
    1.4795982506629979e-11, 1.5184007323856147e-11, 1.5569476133085627e-11, 
    1.594757917757964e-11, 1.6313608333238329e-11, 1.6662971839986835e-11, 
    1.6991228074403774e-11, 1.7294158780135748e-11, 1.756786916442761e-11, 
    1.780890457507411e-11, 1.8014360916103806e-11, 1.8181970605102909e-11, 
    1.8310152257411152e-11, 1.8398011985930009e-11, 1.8445301435224818e-11, 
    1.8452320528055627e-11, 1.8419813508071498e-11, 1.8348838741849906e-11, 
    1.8240670366442361e-11, 1.8096718245445186e-11, 1.7918526369014545e-11, 
    1.7707793358115133e-11, 1.7466478406650143e-11, 1.719692377061207e-11, 
    1.6902008268611776e-11, 1.6585271077511122e-11, 1.6251007049367062e-11, 
    1.5904267400265276e-11, 1.5550796329238817e-11, 1.5196827156408752e-11, 
    1.4848817565227458e-11, 1.4513095609673905e-11, 1.4195480849245857e-11, 
    1.3900885918281266e-11, 1.3633000792260198e-11, 1.3394050133590845e-11, 
    1.31847019255666e-11, 1.3004114898522063e-11, 1.2850153684241724e-11, 
    1.271973037669269e-11, 1.2609258713407779e-11, 1.2515154023758889e-11, 
    1.2434330950589567e-11, 1.2364627678266837e-11, 1.2305118071324396e-11, 
    1.2256246322923729e-11, 1.2219789558950222e-11, 1.2198620986263694e-11, 
    1.2196320510540704e-11, 1.221664243368816e-11, 1.2262925909671038e-11, 
    1.2337504411674822e-11, 1.244120866789396e-11, 1.2572929066103202e-11, 
    1.2729448596580519e-11, 1.2905420826981137e-11, 1.309360727013666e-11, 
    1.3285294635117324e-11, 1.3470888385249322e-11, 1.3640594542533079e-11, 
    1.3785161070496321e-11, 1.3896544640762642e-11, 1.3968504376214248e-11, 
    1.3996983623368782e-11, 1.3980324157427511e-11, 1.3919225911824727e-11, 
    1.3816516072781668e-11, 1.3676725356117362e-11, 1.3505563015223262e-11, 
    1.3309299176119633e-11, 1.3094210258005665e-11, 1.286605587054017e-11, 
    1.2629735758660344e-11, 1.2389080152685944e-11, 1.2146863567433538e-11, 
    1.1904948086506331e-11, 1.1664593866140574e-11, 1.1426870852873467e-11, 
    1.1193103615163835e-11, 1.0965261678870481e-11, 1.0746320714640317e-11, 
    1.0540459708995593e-11, 1.035312813853258e-11, 1.0190913743572908e-11, 
    1.0061278656799861e-11, 9.9721114067574691e-12, 9.9312006238685873e-12, 
    9.9456204120461574e-12, 1.0021124024858851e-11, 1.0161552371033416e-11, 
    1.0368362448550032e-11, 1.0640267482549403e-11, 1.0973060381289836e-11, 
    1.1359623549164686e-11, 1.17901523619074e-11, 1.2252524958853556e-11, 
    1.2732895256504278e-11, 1.3216366483322186e-11, 1.3687784413979757e-11, 
    1.4132538513565779e-11, 1.4537350744466331e-11, 1.489097704366823e-11, 
    1.5184789411165434e-11, 1.5413178322964289e-11, 1.5573777761358885e-11, 
    1.5667458700155222e-11, 1.5698171804455624e-11, 1.5672526756938962e-11, 
    1.5599285115312138e-11, 1.5488711788464251e-11, 1.5351855396985859e-11, 
    1.5199809157781441e-11, 1.504300542530435e-11, 1.4890583325132019e-11, 
    1.4749872461837662e-11, 1.4626024207782711e-11, 1.452181897077591e-11, 
    1.4437645911805428e-11, 1.4371677339146062e-11, 1.4320211567992409e-11, 
    1.4278164594520108e-11, 1.4239670754277598e-11, 1.4198746179462674e-11, 
    1.4149968324812289e-11, 1.4089103219980733e-11, 1.4013635520428038e-11, 
    1.3923148035044303e-11, 1.3819506564883915e-11, 1.3706829435016381e-11, 
    1.3591274093580111e-11, 1.3480605529985091e-11, 1.3383619302990499e-11, 
    1.3309474063447993e-11, 1.3266973851943478e-11, 1.3263889403788265e-11, 
    1.3306353250908209e-11, 1.3398401322155916e-11, 1.3541680294478952e-11, 
    1.3735326014601608e-11, 1.3976037180198842e-11, 1.4258283984055256e-11, 
    1.457465020944291e-11, 1.4916242415522352e-11, 1.5273158735121869e-11, 
    1.5634940302182772e-11, 1.5991005285831873e-11, 1.6331047452591934e-11, 
    1.6645381594878778e-11, 1.6925239322626315e-11, 1.7163042182765789e-11, 
    1.7352631529363474e-11, 1.748948552254283e-11, 1.7570897548942824e-11, 
    1.759615213596026e-11, 1.7566631110163475e-11, 1.7485856462100311e-11, 
    1.7359458200752433e-11, 1.7195009620204372e-11, 1.7001765753288863e-11, 
    1.6790244320212514e-11, 1.6571719624170122e-11, 1.6357589111199363e-11, 
    1.6158710885216167e-11, 1.598470761327809e-11, 1.5843325268159347e-11, 
    1.5739876646345238e-11, 1.5676818312816666e-11, 1.5653536028061842e-11, 
    1.5666312600006711e-11, 1.5708515225013417e-11, 1.5770982801147402e-11, 
    1.58426082223613e-11, 1.5911056947109189e-11, 1.5963532647985975e-11, 
    1.5987618239847694e-11, 1.597205467532247e-11, 1.5907422304196295e-11, 
    1.5786698098969438e-11, 1.5605625090612834e-11, 1.5362880293158762e-11, 
    1.5060062854181744e-11, 1.4701473106781655e-11, 1.4293740482006216e-11, 
    1.384535506868443e-11, 1.336610832363241e-11, 1.2866506838074131e-11, 
    1.2357218818137333e-11, 1.1848578241943017e-11, 1.1350166644813742e-11, 
    1.0870508478730227e-11, 1.0416849873265951e-11, 9.9950676075356901e-12, 
    9.6096338667933319e-12, 9.2636646375683232e-12, 8.9590110945738148e-12, 
    8.6963931189311286e-12, 8.4755375831408267e-12, 8.295347202702537e-12, 
    8.1540626765112049e-12, 8.0494448911417552e-12, 7.9789461200627619e-12, 
    7.9399090378648481e-12, 7.9297319088056372e-12, 7.9460463540561362e-12, 
    7.9868436399243214e-12, 8.0505786346893055e-12, 8.1361890268340082e-12, 
    8.2430608815814229e-12, 8.3709107886586138e-12, 8.5195986636259469e-12, 
    8.6888718672701977e-12, 8.8781311058460437e-12, 9.0861332010458827e-12, 
    9.3108192886857179e-12, 9.5491733086563155e-12, 9.7972110559636283e-12, 
    1.0050095234137846e-11, 1.0302390284058352e-11, 1.0548405993286067e-11, 
    1.0782630540559785e-11, 1.1000175433518352e-11, 1.1197208398520369e-11, 
    1.1371278552875176e-11, 1.1521543603718673e-11, 1.1648799729973142e-11, 
    1.1755382251446319e-11, 1.1844874519670168e-11, 1.1921690876195651e-11, 
    1.1990582785523796e-11, 1.2056105664403296e-11, 1.2122128210400677e-11, 
    1.2191428180568851e-11, 1.2265427136164115e-11, 1.2344090229297416e-11, 
    1.2426006631111403e-11, 1.2508636022031245e-11, 1.2588694410172605e-11, 
    1.266264348322508e-11, 1.272721297503173e-11, 1.2779901430518534e-11, 
    1.2819422904518623e-11, 1.2845997683970336e-11, 1.2861514181747702e-11, 
    1.2869484949631282e-11, 1.2874830090907994e-11, 1.2883489936558677e-11, 
    1.2901887527233936e-11, 1.2936324118716883e-11, 1.2992332415362364e-11, 
    1.307403978082818e-11, 1.3183650481688582e-11, 1.3321060446361916e-11, 
    1.3483664063902772e-11, 1.3666368312884161e-11, 1.3861838127296321e-11, 
    1.4060940439753183e-11, 1.425335973905694e-11, 1.4428337186267776e-11, 
    1.4575463002436626e-11, 1.4685436629107544e-11, 1.4750767410573676e-11, 
    1.4766305392022332e-11, 1.4729591604460669e-11, 1.4640979535471654e-11, 
    1.4503542878840253e-11, 1.4322750909194778e-11, 1.4105988832185011e-11, 
    1.3861931964521359e-11, 1.3599873304376414e-11, 1.332901960676884e-11, 
    1.305786388574433e-11, 1.2793646700467903e-11, 1.2541973062900046e-11, 
    1.2306581155407486e-11, 1.2089301714621178e-11, 1.1890171707378814e-11, 
    1.1707708237929801e-11, 1.1539284283192005e-11, 1.1381585505311297e-11, 
    1.1231101835988527e-11, 1.1084589804061984e-11, 1.093950460443052e-11, 
    1.0794320695789048e-11, 1.0648737979522008e-11, 1.0503764170755116e-11, 
    1.0361650970573798e-11, 1.0225707471134605e-11, 1.0099999263899658e-11, 
    9.9889752998917628e-12, 9.8970522500256125e-12, 9.8281904328199117e-12, 
    9.7855269773721453e-12, 9.7710733514645748e-12,
  // Sqw-total(3, 0-1999)
    0.059404233212714076, 0.059308920163845293, 0.059025018429395303, 
    0.05855854092259806, 0.057919185734532058, 0.0571198769451556, 
    0.056176170882820654, 0.055105570821353062, 0.053926797531044762, 
    0.052659063069613432, 0.051321391031465505, 0.049932018940058394, 
    0.048507908654617266, 0.047064379799071542, 0.045614870509003057, 
    0.044170820254442675, 0.042741661871904861, 0.041334904634005215, 
    0.039956287276913117, 0.038609979195154846, 0.037298809104756935, 
    0.036024502872447565, 0.034787915399888417, 0.033589244982434971, 
    0.032428222074240343, 0.031304267640491552, 0.030216619121268554, 
    0.029164424406925956, 0.028146806117866831, 0.027162899900196422, 
    0.026211871405986072, 0.025292917135094375, 0.024405254391132492, 
    0.023548105278522882, 0.022720678997621639, 0.021922155768908096, 
    0.021151674651854864, 0.020408326451793708, 0.019691151957836907, 
    0.018999145030380946, 0.018331259617697989, 0.017686419633198926, 
    0.017063530720387302, 0.01646149318265298, 0.015879215651419403, 
    0.015315629305571534, 0.014769702562660997, 0.014240456107240293, 
    0.013726977921818487, 0.013228437701476038, 0.012744099749866301, 
    0.012273333261668998, 0.011815618865715643, 0.011370550469861811, 
    0.010937831805450235, 0.010517267566446093, 0.010108749596016903, 
    0.009712239098445246, 0.0093277462601691463, 0.0089553088874251459, 
    0.0085949716811740094, 0.0082467675826596483, 0.0079107022785336392, 
    0.0075867425190193211, 0.0072748084503011946, 0.0069747697610487765, 
    0.0066864451425034683, 0.0064096043869198037, 0.0061439723997021309, 
    0.0058892344542828597, 0.0056450421401491166, 0.0054110196039208712, 
    0.0051867698260823509, 0.0049718807876911585, 0.0047659314513338593, 
    0.0045684975105115258, 0.0043791568622236678, 0.0041974947434976215, 
    0.0040231084577903725, 0.0038556116109113529, 0.0036946377816380739, 
    0.0035398435672594542, 0.0033909109632009743, 0.0032475490524540734, 
    0.0031094949906090622, 0.002976514275436003, 0.0028484002895707919, 
    0.0027249731070003703, 0.0026060775652659079, 0.002491580630361884, 
    0.0023813681212554094, 0.002275340912344295, 0.0021734107874866195, 
    0.0020754961684289613, 0.0019815179731864424, 0.0018913958679083324, 
    0.0018050451546392562, 0.0017223744877365985, 0.0016432845389432738, 
    0.0015676676444541554, 0.0014954083780006581, 0.0014263849133087558, 
    0.0013604709767448754, 0.0012975381529082297, 0.0012374582949171511, 
    0.0011801058060223774, 0.00112535959573681, 0.0010731045656370926, 
    0.0010232325401935472, 0.00097564261940185487, 0.00093024098653858881, 
    0.0008869402514009154, 0.00084565844388226493, 0.00080631779321687627, 
    0.00076884343458274865, 0.0007331621779828292, 0.0006992014562573522, 
    0.00066688854217901645, 0.00063615009172996676, 0.00060691203501179515, 
    0.00057909980101956277, 0.00055263883081976318, 0.0005274553082363733, 
    0.00050347702009255816, 0.00048063425066757043, 0.00045886061762765709, 
    0.00043809376855879931, 0.00041827587669765676, 0.00039935389907781472, 
    0.00038127958716243656, 0.00036400926606652454, 0.00034750342087210695, 
    0.0003317261450541697, 0.00031664451522933499, 0.00030222795781485821, 
    0.00028844766720344402, 0.0002752761230112863, 0.00026268673776290501, 
    0.00025065364829039439, 0.00023915164643864708, 0.00022815622940960208, 
    0.00021764373878860273, 0.00020759155086621579, 0.00019797827950415929, 
    0.00018878395604490997, 0.00017999015767515612, 0.0001715800649322563, 
    0.00016353843929200692, 0.00015585152167597006, 0.00014850686120204259, 
    0.00014149308985140572, 0.00013479966260777841, 0.00012841658406041975, 
    0.00012233414175958032, 0.0001165426642506575, 0.00011103231824900318, 
    0.00010579295537614878, 0.00010081401470293622, 9.6084483348339526e-05, 
    9.159291375960322e-05, 8.7327493139384158e-05, 8.3276157821157002e-05, 
    7.9426743228425047e-05, 7.576715840257267e-05, 7.2285572981666986e-05, 
    6.8970604021417896e-05, 6.5811490234476979e-05, 6.2798242142489332e-05, 
    5.9921758295891415e-05, 5.7173900075067717e-05, 5.4547520518377293e-05, 
    5.2036445939818913e-05, 4.9635412549023746e-05, 4.7339963590097642e-05, 
    4.5146315384529478e-05, 4.305120284270872e-05, 4.1051716294909905e-05, 
    3.9145141768034478e-05, 3.7328816069163457e-05, 3.5600006306438049e-05, 
    3.3955820945611e-05, 3.2393156417046788e-05, 3.0908679954405812e-05, 
    2.9498846098108423e-05, 2.8159941456280806e-05, 2.6888150167678443e-05, 
    2.5679631256442463e-05, 2.4530598810960782e-05, 2.3437396636797817e-05, 
    2.2396560593632998e-05, 2.1404863987666266e-05, 2.0459343851737839e-05, 
    1.9557308372034589e-05, 1.8696327809077675e-05, 1.7874212769348962e-05, 
    1.7088984477901957e-05, 1.6338841756797042e-05, 1.5622128824593836e-05, 
    1.4937306976156776e-05, 1.4282931916364789e-05, 1.3657637244037523e-05, 
    1.3060123522332701e-05, 1.2489151664599633e-05, 1.1943539066006438e-05, 
    1.1422156987762771e-05, 1.0923928057103316e-05, 1.0447823243856542e-05, 
    9.9928581758955451e-06, 9.5580890431729652e-06, 9.1426085493691013e-06, 
    8.7455423857583701e-06, 8.3660465646906622e-06, 8.003305727953634e-06, 
    7.6565323235483606e-06, 7.3249663905251693e-06, 7.0078756497272383e-06, 
    6.7045556706365957e-06, 6.4143300417808921e-06, 6.1365506573342357e-06, 
    5.8705983838240037e-06, 5.6158844327676814e-06, 5.3718527094369653e-06, 
    5.13798323419282e-06, 4.9137964749831232e-06, 4.6988581408858019e-06, 
    4.4927837336641464e-06, 4.2952419953246609e-06, 4.1059563680315065e-06, 
    3.9247037119402653e-06, 3.7513097941135877e-06, 3.5856414267262305e-06, 
    3.4275955406505615e-06, 3.2770858678975301e-06, 3.1340282187663154e-06, 
    2.9983255337184003e-06, 2.8698539468551406e-06, 2.7484510150467735e-06, 
    2.6339070655754365e-06, 2.5259603250642843e-06, 2.4242961546232799e-06, 
    2.3285503672694176e-06, 2.2383162801874632e-06, 2.1531548805508363e-06, 
    2.0726072787954361e-06, 1.9962084945516693e-06, 1.9235015713648664e-06, 
    1.8540510423710384e-06, 1.7874548643237282e-06, 1.7233540910453335e-06, 
    1.6614397580041383e-06, 1.6014566812621196e-06, 1.5432041202733833e-06, 
    1.4865334938913003e-06, 1.4313435539491913e-06, 1.3775735901298009e-06, 
    1.3251953499637344e-06, 1.2742043978243642e-06, 1.2246116069012747e-06, 
    1.1764353835997235e-06, 1.1296950815744758e-06, 1.0844058908933861e-06, 
    1.0405753120260658e-06, 9.9820116417906278e-07, 9.5727095257406452e-07, 
    9.1776233792911932e-07, 8.7964441792141609e-07, 8.4287953748699482e-07, 
    8.074253825635873e-07, 7.7323716426031365e-07, 7.4026975431052207e-07, 
    7.0847967492154001e-07, 6.7782687187194139e-07, 6.482762067398174e-07, 
    6.1979859892068402e-07, 5.9237173794987376e-07, 5.6598028316702718e-07, 
    5.4061547857611993e-07, 5.1627414269046393e-07, 4.9295704512153093e-07, 
    4.7066674993685172e-07, 4.4940507904225169e-07, 4.2917041587989332e-07, 
    4.0995511592377579e-07, 3.9174330692117714e-07, 3.7450934071611757e-07, 
    3.5821710163229957e-07, 3.4282028826944534e-07, 3.2826367936147359e-07, 
    3.1448528315181461e-07, 3.0141917057344968e-07, 2.8899871743163731e-07, 
    2.7715994042632923e-07, 2.6584460880359698e-07, 2.5500284747024283e-07, 
    2.4459500999058132e-07, 2.3459268289417242e-07, 2.2497877278821126e-07, 
    2.1574671556158213e-07, 2.0689892197849877e-07, 1.9844463153956111e-07, 
    1.9039738210409118e-07, 1.8277231794947118e-07, 1.7558355352246584e-07, 
    1.6884178930270573e-07, 1.6255234138054374e-07, 1.5671370343478184e-07, 
    1.5131671043521298e-07, 1.4634432312524013e-07, 1.4177200290577949e-07, 
    1.375686038003938e-07, 1.336976729790864e-07, 1.3011902887079839e-07, 
    1.267904759258781e-07, 1.23669519877699e-07, 1.2071496372436903e-07, 
    1.178882914130037e-07, 1.1515477747204172e-07, 1.124842936438732e-07, 
    1.0985181176709424e-07, 1.0723762434373348e-07, 1.0462731683205782e-07, 
    1.0201153110147032e-07, 9.938555750496492e-08, 9.6748788525914988e-08, 
    9.4104061619627355e-08, 9.1456916781009491e-08, 8.8814795437300455e-08, 
    8.6186212918354818e-08, 8.357994377264424e-08, 8.1004266584102989e-08, 
    7.8466317936764555e-08, 7.5971603402217012e-08, 7.3523703495676797e-08, 
    7.1124196927269075e-08, 6.8772802036627504e-08, 6.6467714895074186e-08, 
    6.4206101167342339e-08, 6.1984683415419193e-08, 5.9800356879896939e-08, 
    5.7650767667543191e-08, 5.5534795531603196e-08, 5.3452898840688289e-08, 
    5.1407297551159697e-08, 4.9401989491709701e-08, 4.7442611843373131e-08, 
    4.5536172773438907e-08, 4.3690685402067415e-08, 4.1914739192400021e-08, 
    4.0217041936187624e-08, 3.8605961485030255e-08, 3.7089090513183829e-08, 
    3.5672852292766513e-08, 3.436216036020019e-08, 3.3160141684616129e-08, 
    3.206793002029267e-08, 3.1084534720546874e-08, 3.0206788514027072e-08, 
    2.9429376668476955e-08, 2.874494789004216e-08, 2.8144305621917575e-08, 
    2.7616675630603993e-08, 2.7150043242212091e-08, 2.6731550293461172e-08, 
    2.6347938902281835e-08, 2.59860254844677e-08, 2.563318567522921e-08, 
    2.5277827600407606e-08, 2.4909829407694313e-08, 2.4520915848741579e-08, 
    2.4104950040851804e-08, 2.3658119154798875e-08, 2.3178998095782901e-08, 
    2.2668481949415692e-08, 2.2129586777748885e-08, 2.1567127368563704e-08, 
    2.0987290238237239e-08, 2.0397128385880399e-08, 1.9804011323713235e-08, 
    1.9215067972325533e-08, 1.8636661696564748e-08, 1.8073934728538923e-08, 
    1.7530454763600259e-08, 1.7007988675325209e-08, 1.6506419003547526e-08, 
    1.602380753363834e-08, 1.5556599252521578e-08, 1.5099948720543032e-08, 
    1.464814192148744e-08, 1.4195079253563238e-08, 1.3734781628609666e-08, 
    1.3261880536196998e-08, 1.277205593022469e-08, 1.2262391080720635e-08, 
    1.1731621880360779e-08, 1.1180267322410552e-08, 1.0610638178670994e-08, 
    1.0026730008435238e-08, 9.434014910409231e-09, 8.8391519625882201e-09, 
    8.2496399426593838e-09, 7.6734366074505519e-09, 7.1185680735611838e-09, 
    6.5927488418004581e-09, 6.1030301024955814e-09, 5.6554899873921188e-09, 
    5.2549766247156179e-09, 4.904911867916196e-09, 4.6071617277552536e-09, 
    4.361977446590478e-09, 4.1680094947242654e-09, 4.0223941533980384e-09, 
    3.9209096917511475e-09, 3.8581951441561856e-09, 3.8280209719752206e-09, 
    3.8235966519663006e-09, 3.837897132021014e-09, 3.8639879054506415e-09, 
    3.895328367380848e-09, 3.9260346745584814e-09, 3.9510872552592373e-09, 
    3.9664729614434622e-09, 3.9692581806351198e-09, 3.9575950355218897e-09, 
    3.9306683218717803e-09, 3.8885946065785988e-09, 3.8322872898945807e-09, 
    3.7633015906090836e-09, 3.6836724593270759e-09, 3.5957557595742548e-09, 
    3.5020804888237581e-09, 3.4052166439732829e-09, 3.3076612367506524e-09, 
    3.2117431383166281e-09, 3.1195467978141784e-09, 3.0328545001965093e-09, 
    2.9531072505428657e-09, 2.8813842088244475e-09, 2.8184007867067604e-09, 
    2.7645246574481999e-09, 2.7198081060957348e-09, 2.6840336302413388e-09, 
    2.6567685512794955e-09, 2.6374230926087156e-09, 2.6253061805743469e-09, 
    2.6196732655603812e-09, 2.6197617598690441e-09, 2.6248113124066212e-09, 
    2.6340685216228872e-09, 2.646777830854391e-09, 2.6621625448805496e-09, 
    2.6794012319038269e-09, 2.6976055648541703e-09, 2.7158052844185118e-09, 
    2.7329451121210417e-09, 2.7478965243054765e-09, 2.7594854316557849e-09, 
    2.7665343779477418e-09, 2.7679161389419486e-09, 2.7626137706684156e-09, 
    2.749781496721875e-09, 2.7288003239944321e-09, 2.6993229618944435e-09, 
    2.6613035114241602e-09, 2.6150090603340325e-09, 2.5610119704267507e-09, 
    2.5001636792334977e-09, 2.4335522912759582e-09, 2.3624478436191449e-09, 
    2.2882397819084333e-09, 2.2123718023758712e-09, 2.1362787614042841e-09, 
    2.0613300050942476e-09, 1.9887822185208027e-09, 1.9197438744777473e-09, 
    1.8551519093780096e-09, 1.7957602718161515e-09, 1.7421387960020332e-09, 
    1.6946804380965373e-09, 1.6536143220541552e-09, 1.6190223029853146e-09, 
    1.5908568025452501e-09, 1.5689583441301498e-09, 1.5530716568302948e-09, 
    1.542859931910876e-09, 1.5379172304177044e-09, 1.5377795640534432e-09, 
    1.5419352334606189e-09, 1.5498351728796739e-09, 1.5609038069446931e-09, 
    1.5745507718408179e-09, 1.5901834060173318e-09, 1.6072198058807356e-09, 
    1.6251017166410513e-09, 1.6433066658741416e-09, 1.6613583872093904e-09, 
    1.6788349892956741e-09, 1.6953741576163999e-09, 1.7106752301473676e-09, 
    1.724497990461557e-09, 1.7366584925696365e-09, 1.7470222617473754e-09, 
    1.7554955348470779e-09, 1.7620151559664076e-09, 1.7665379503250526e-09, 
    1.7690301478553187e-09, 1.7694577029251601e-09, 1.7677779791255514e-09, 
    1.7639335115652992e-09, 1.7578481777260994e-09, 1.7494263399684863e-09, 
    1.7385550985780754e-09, 1.7251099130202458e-09, 1.7089633848987911e-09, 
    1.6899970504880602e-09, 1.6681154644466112e-09, 1.6432618418948037e-09, 
    1.6154340632139987e-09, 1.5846998417732325e-09, 1.5512095693897572e-09, 
    1.5152055526334507e-09, 1.4770263008579913e-09, 1.437105017315802e-09, 
    1.3959616494251092e-09, 1.3541885175334645e-09, 1.3124299051797942e-09, 
    1.2713567152578911e-09, 1.2316375841724914e-09, 1.1939084258293697e-09, 
    1.1587423532051834e-09, 1.1266222641229686e-09, 1.097917981267153e-09, 
    1.0728697326839218e-09, 1.0515790940018039e-09, 1.0340081521768518e-09, 
    1.0199868122629341e-09, 1.0092276867487592e-09, 1.0013472995246909e-09, 
    9.9589202545839143e-10, 9.9236667938153345e-10, 9.9026376548057598e-10, 
    9.8909119702871752e-10, 9.8839676594909812e-10, 9.877877515542501e-10, 
    9.8694475883038214e-10, 9.8562919567760968e-10, 9.8368446486853887e-10, 
    9.8103130959220649e-10, 9.7765828530486571e-10, 9.7360849017409361e-10, 
    9.6896400907373122e-10, 9.6382942540193202e-10, 9.5831586074655617e-10, 
    9.5252668017024299e-10, 9.4654590921163606e-10, 9.4042996580754601e-10, 
    9.3420314665834947e-10, 9.278568098279973e-10, 9.2135208584262512e-10, 
    9.146255131489358e-10, 9.0759696286210329e-10, 9.0017891793936864e-10, 
    8.9228632837728713e-10, 8.8384606146962546e-10, 8.7480527475146288e-10, 
    8.651379243226361e-10, 8.5484911154561113e-10, 8.4397684777799316e-10, 
    8.3259127846788814e-10, 8.2079140182166393e-10, 8.086996502620015e-10, 
    7.9645469419486169e-10, 7.8420307277293189e-10, 7.7209018458966441e-10, 
    7.6025134591373476e-10, 7.4880347483465777e-10, 7.3783807411121792e-10, 
    7.2741593221877212e-10, 7.1756403521697882e-10, 7.0827484101295248e-10, 
    6.9950812835787788e-10, 6.9119516887498881e-10, 6.8324508916472526e-10, 
    6.7555281233399051e-10, 6.6800811636825872e-10, 6.6050494781685237e-10, 
    6.5295038225048976e-10, 6.4527237167133114e-10, 6.3742573169998152e-10, 
    6.2939576343217693e-10, 6.2119928516290237e-10, 6.1288288071948476e-10, 
    6.0451859279007992e-10, 5.961973066620857e-10, 5.8802048712869615e-10, 
    5.8009083679862608e-10, 5.7250276657564108e-10, 5.6533340468246813e-10, 
    5.5863498712526102e-10, 5.5242920371959772e-10, 5.4670414237473692e-10, 
    5.4141400263050489e-10, 5.3648180455587574e-10, 5.3180479712475487e-10, 
    5.2726230231116714e-10, 5.2272525716596434e-10, 5.1806681281081329e-10, 
    5.1317298006155634e-10, 5.0795254803882846e-10, 5.0234529938549929e-10, 
    4.9632793721701474e-10, 4.8991707282716962e-10, 4.8316916461258769e-10, 
    4.7617726565819498e-10, 4.6906504014204381e-10, 4.6197843415400423e-10, 
    4.5507583640091314e-10, 4.4851744293957251e-10, 4.4245477342413101e-10, 
    4.3702103760119493e-10, 4.3232310111080158e-10, 4.2843545347557772e-10, 
    4.253965748950865e-10, 4.2320765674245723e-10, 4.2183372343249649e-10, 
    4.2120676073368049e-10, 4.212305926234609e-10, 4.2178695837883762e-10, 
    4.2274241644781178e-10, 4.2395550963229662e-10, 4.2528384455817664e-10, 
    4.2659061790439886e-10, 4.277503593613323e-10, 4.2865357375845124e-10, 
    4.2921019159551501e-10, 4.2935169902555859e-10, 4.2903199134442414e-10, 
    4.2822693808299187e-10, 4.2693291935168585e-10, 4.2516435519232934e-10, 
    4.2295060649137028e-10, 4.2033238116063236e-10, 4.1735797529559549e-10, 
    4.1407954779115339e-10, 4.1054973240137918e-10, 4.068187001978176e-10, 
    4.0293193479585401e-10, 3.9892872449857934e-10, 3.9484154742047188e-10, 
    3.9069621168262488e-10, 3.865128010478008e-10, 3.8230722407964503e-10, 
    3.7809324630160821e-10, 3.73884708600284e-10, 3.6969778826293473e-10, 
    3.6555294607342482e-10, 3.6147641951307734e-10, 3.5750094966323368e-10, 
    3.5366571361768288e-10, 3.5001532076307451e-10, 3.4659796066700508e-10, 
    3.434627476113106e-10, 3.4065658269357041e-10, 3.3822066269773106e-10, 
    3.3618708642528932e-10, 3.3457575908775764e-10, 3.3339199231441082e-10, 
    3.3262495565014094e-10, 3.3224723026647875e-10, 3.3221545014184551e-10, 
    3.3247208674994119e-10, 3.3294816656756223e-10, 3.3356678584852783e-10, 
    3.3424708385345788e-10, 3.3490843815815189e-10, 3.3547450153732868e-10, 
    3.358768865449971e-10, 3.3605817561131125e-10, 3.3597419844246448e-10, 
    3.3559540222980559e-10, 3.3490738781670505e-10, 3.3391060121804881e-10, 
    3.3261936297727746e-10, 3.3106026740643186e-10, 3.292702092940791e-10, 
    3.2729407653896112e-10, 3.2518228765431149e-10, 3.2298821983304892e-10, 
    3.2076565329943428e-10, 3.1856623624839654e-10, 3.1643710074604107e-10, 
    3.1441862730767526e-10, 3.1254251708188216e-10, 3.1083018477086125e-10, 
    3.0929164251602264e-10, 3.0792490770530752e-10, 3.067160661591635e-10, 
    3.056399587732404e-10, 3.0466158405464675e-10, 3.0373805031117048e-10, 
    3.0282109966516094e-10, 3.0185994649843803e-10, 3.0080433057538708e-10, 
    2.9960753172914199e-10, 2.9822920191773095e-10, 2.9663775421946746e-10, 
    2.9481223883940479e-10, 2.927435080225445e-10, 2.9043466983623341e-10, 
    2.8790077005330691e-10, 2.8516778876071779e-10, 2.822709750706846e-10, 
    2.7925273878180475e-10, 2.7616016465591909e-10, 2.7304241547461532e-10, 
    2.6994812665930451e-10, 2.6692302238272313e-10, 2.6400786776389974e-10, 
    2.6123687750180777e-10, 2.5863661578537797e-10, 2.5622547110292824e-10, 
    2.540136001303406e-10, 2.5200336287854778e-10, 2.5019007020404141e-10, 
    2.4856302599647714e-10, 2.4710669837916846e-10, 2.4580196077315658e-10, 
    2.4462729047824609e-10, 2.435599226879497e-10, 2.4257687657239728e-10, 
    2.4165588425188384e-10, 2.4077619808441307e-10, 2.3991929870599108e-10, 
    2.3906948761687972e-10, 2.3821438580582176e-10, 2.3734526605666948e-10, 
    2.3645726395068272e-10, 2.3554936614015685e-10, 2.3462420106604815e-10, 
    2.3368757718094652e-10, 2.327478130258383e-10, 2.3181485215062918e-10, 
    2.308992614487016e-10, 2.3001115799979967e-10, 2.2915919826767839e-10, 
    2.2834967388787494e-10, 2.2758587115425813e-10, 2.2686769732268636e-10, 
    2.261916628042937e-10, 2.255511690855249e-10, 2.2493713218404637e-10, 
    2.24338786530918e-10, 2.237446740712836e-10, 2.2314364151680747e-10, 
    2.2252580144747085e-10, 2.2188330966735508e-10, 2.2121095227850911e-10, 
    2.2050642455413672e-10, 2.197703704437899e-10, 2.1900609975578276e-10, 
    2.1821909906507329e-10, 2.1741631681966501e-10, 2.1660533903843564e-10, 
    2.1579348775024482e-10, 2.1498693703270828e-10, 2.1418988488974506e-10, 
    2.1340388491727289e-10, 2.1262732019415914e-10, 2.1185513285748338e-10, 
    2.1107878314902272e-10, 2.1028649557539428e-10, 2.0946371585337453e-10, 
    2.0859387543185933e-10, 2.0765930932155361e-10, 2.0664238488577713e-10, 
    2.055266959774602e-10, 2.0429830504047429e-10, 2.0294689234138555e-10, 
    2.0146679693545686e-10, 1.998577594995732e-10, 1.9812541122937456e-10, 
    1.962813496022454e-10, 1.9434284234174264e-10, 1.9233210549873706e-10, 
    1.9027523685313075e-10, 1.8820082961880982e-10, 1.8613839390117969e-10, 
    1.8411667229147699e-10, 1.8216201253565072e-10, 1.8029685728769282e-10, 
    1.7853854507921132e-10, 1.7689844384446798e-10, 1.7538149924962619e-10, 
    1.7398623081650059e-10, 1.7270514769169405e-10, 1.7152552605032987e-10, 
    1.7043051978530477e-10, 1.6940044847571638e-10, 1.6841424243255101e-10, 
    1.6745084871850818e-10, 1.6649059828277816e-10, 1.6551636464957802e-10, 
    1.6451451525398313e-10, 1.6347554220600203e-10, 1.623944127121839e-10, 
    1.6127054524649708e-10, 1.6010750388805657e-10, 1.589123724044741e-10, 
    1.5769492513865074e-10, 1.5646657613795857e-10, 1.55239289837043e-10, 
    1.5402446709282461e-10, 1.5283194142202127e-10, 1.5166915259474693e-10, 
    1.5054060661201347e-10, 1.494476077710886e-10, 1.4838836136525953e-10, 
    1.4735835603798359e-10, 1.463510535110928e-10, 1.4535872007640788e-10, 
    1.4437340013720467e-10, 1.4338785408482848e-10, 1.4239640947895692e-10, 
    1.4139561005844079e-10, 1.4038465302921251e-10, 1.3936552539313488e-10, 
    1.383429257963235e-10, 1.3732393534993982e-10, 1.363175404409895e-10, 
    1.3533404607965075e-10, 1.3438445077006677e-10, 1.3347984156824162e-10, 
    1.3263085464498907e-10, 1.3184718423629939e-10, 1.3113722449772851e-10, 
    1.3050774616063938e-10, 1.2996368390126037e-10, 1.2950794358795099e-10, 
    1.2914129299894909e-10, 1.2886227144028886e-10, 1.2866718359959315e-10, 
    1.2855012637770185e-10, 1.2850313038379387e-10, 1.2851635706989813e-10, 
    1.2857840944104052e-10, 1.2867668675859424e-10, 1.2879781726779826e-10, 
    1.289280938363779e-10, 1.2905390673238923e-10, 1.2916210393688423e-10, 
    1.2924029933546985e-10, 1.2927707362481062e-10, 1.2926211374978432e-10, 
    1.2918625727114078e-10, 1.2904153072769327e-10, 1.2882117056765232e-10, 
    1.2851969763262743e-10, 1.281330371089565e-10, 1.2765872766953224e-10, 
    1.2709616770403242e-10, 1.2644690523791622e-10, 1.2571489713256117e-10, 
    1.249067025577483e-10, 1.2403152524487369e-10, 1.231010889327741e-10, 
    1.2212931257304171e-10, 1.2113179584956116e-10, 1.201251013501224e-10, 
    1.1912598928520413e-10, 1.1815055461622531e-10, 1.1721348335934949e-10, 
    1.1632738526691638e-10, 1.1550236686152723e-10, 1.1474580417207883e-10, 
    1.1406238474632677e-10, 1.1345430291869294e-10, 1.1292163789966304e-10, 
    1.1246277980127624e-10, 1.1207484386129934e-10, 1.1175396691950042e-10, 
    1.1149550399675099e-10, 1.1129400829605095e-10, 1.1114310279465891e-10, 
    1.1103520551128652e-10, 1.1096123689204893e-10, 1.1091035922443896e-10, 
    1.1086986217052872e-10, 1.1082519481069676e-10, 1.1076028488979379e-10, 
    1.10658063216052e-10, 1.1050124788359022e-10, 1.1027323914108672e-10, 
    1.0995914618528547e-10, 1.0954676151141032e-10, 1.0902745074717701e-10, 
    1.0839681030730952e-10, 1.0765511205448458e-10, 1.068073803624378e-10, 
    1.0586323351473381e-10, 1.0483638829753075e-10, 1.037439781350574e-10, 
    1.0260566857363887e-10, 1.0144273496979118e-10, 1.0027707057922355e-10, 
    9.9130306974702905e-11, 9.8022991592049795e-11, 9.6973941164565718e-11, 
    9.5999708686067908e-11, 9.5114229551755706e-11, 9.4328554899078768e-11, 
    9.3650731611502686e-11, 9.3085722412015611e-11, 9.2635410343308934e-11, 
    9.2298629584633302e-11, 9.2071271141811084e-11, 9.194638564974545e-11, 
    9.191441201035485e-11, 9.1963433187120982e-11, 9.2079566917841716e-11, 
    9.2247412068342616e-11, 9.2450636077904988e-11, 9.2672580251383489e-11, 
    9.2896958849086538e-11, 9.3108511733964158e-11, 9.3293646110021012e-11, 
    9.3440928298277085e-11, 9.3541480448697372e-11, 9.3589156237392087e-11, 
    9.358056324953932e-11, 9.3514849925633972e-11, 9.3393373825307451e-11, 
    9.3219185280372239e-11, 9.2996471571314999e-11, 9.2729945754342383e-11, 
    9.2424294982504516e-11, 9.2083660750086462e-11, 9.1711286357631026e-11, 
    9.1309267160588278e-11, 9.0878487305975504e-11, 9.0418677345628141e-11, 
    8.9928620701784786e-11, 8.9406457440681022e-11, 8.8850083458861744e-11, 
    8.8257535051107825e-11, 8.7627419956978759e-11, 8.695928195766261e-11, 
    8.6253919204908244e-11, 8.551358260749289e-11, 8.4742089050668076e-11, 
    8.3944799827654026e-11, 8.3128500610037858e-11, 8.23011408694741e-11, 
    8.1471536913979555e-11, 8.0648933166311123e-11, 7.984260523293652e-11, 
    7.9061408711145947e-11, 7.8313400085640707e-11, 7.7605486349961786e-11, 
    7.6943204927249895e-11, 7.6330572887545789e-11, 7.5770107128584881e-11, 
    7.5262910146200561e-11, 7.4808906120776654e-11, 7.4407141818156876e-11, 
    7.4056166379565767e-11, 7.3754408316008458e-11, 7.3500580915465551e-11, 
    7.3293987311161081e-11, 7.3134779268587364e-11, 7.3024049079426466e-11, 
    7.2963803734069548e-11, 7.2956738159987216e-11, 7.3005884433049721e-11, 
    7.3114058942858936e-11, 7.3283235242697588e-11, 7.3513847802827967e-11, 
    7.3804094215530831e-11, 7.414930230714923e-11, 7.4541480344774279e-11, 
    7.4969043097744092e-11, 7.5416842303277276e-11, 7.5866453286910846e-11, 
    7.6296795121751825e-11, 7.6684965704587357e-11, 7.7007324417881326e-11, 
    7.7240686969658342e-11, 7.7363576244564609e-11, 7.7357400444346991e-11, 
    7.7207520666553137e-11, 7.6904068698218331e-11, 7.6442520640224938e-11, 
    7.5823949345383734e-11, 7.5054993922804406e-11, 7.4147483120652162e-11, 
    7.3117866129728517e-11, 7.198639701229252e-11, 7.0776203121787791e-11, 
    6.9512258085581695e-11, 6.8220372362063267e-11, 6.6926196844871185e-11, 
    6.5654349807412803e-11, 6.4427653121770563e-11, 6.3266536538650653e-11, 
    6.2188588298595896e-11, 6.1208290901059922e-11, 6.0336883227044456e-11, 
    5.9582390046465164e-11, 5.8949714004792869e-11, 5.844085423402693e-11, 
    5.8055140190372545e-11, 5.7789511100051227e-11, 5.7638795615199984e-11, 
    5.7595979595063805e-11, 5.7652437845537334e-11, 5.7798173464326388e-11, 
    5.8022006645148208e-11, 5.8311786288694474e-11, 5.8654582460303129e-11, 
    5.9036916357687451e-11, 5.9444990289966938e-11, 5.9864972180398981e-11, 
    6.0283288236643922e-11, 6.068695381645348e-11, 6.1063906254268728e-11, 
    6.1403350285477152e-11, 6.1696075656242337e-11, 6.1934777437132562e-11, 
    6.2114297985096343e-11, 6.2231848671916416e-11, 6.2287131456282122e-11, 
    6.2282418890343352e-11, 6.2222478494562695e-11, 6.2114443849162219e-11, 
    6.1967518203018449e-11, 6.1792592377354287e-11, 6.1601719212307643e-11, 
    6.1407517021765622e-11, 6.1222472095291493e-11, 6.1058253735968725e-11, 
    6.0925006787460177e-11, 6.0830756581776502e-11, 6.0780895839048356e-11, 
    6.0777859833846041e-11, 6.0820962651638297e-11, 6.0906453913256627e-11, 
    6.1027734093147289e-11, 6.1175753521952892e-11, 6.1339519330192424e-11, 
    6.150669905052912e-11, 6.1664233350594355e-11, 6.1798962096818122e-11, 
    6.1898188144068576e-11, 6.1950195491724074e-11, 6.1944651207294031e-11, 
    6.1872966197194981e-11, 6.1728540949260348e-11, 6.1506968368386757e-11, 
    6.1206139614356491e-11, 6.0826319747442198e-11, 6.0370135086799888e-11, 
    5.984252651642206e-11, 5.9250600727902589e-11, 5.8603458687052626e-11, 
    5.7911899101033282e-11, 5.7188098335652805e-11, 5.6445196539140195e-11, 
    5.5696865935060983e-11, 5.4956803262612699e-11, 5.423825247588335e-11, 
    5.3553503914772472e-11, 5.2913434405210585e-11, 5.2327089819111047e-11, 
    5.180133813554256e-11, 5.1340594320978255e-11, 5.0946659698212718e-11, 
    5.061864268054056e-11, 5.0353037643983657e-11, 5.0143878635204468e-11, 
    4.9983057270344117e-11, 4.9860739210812649e-11, 4.9765886542141899e-11, 
    4.9686856901987175e-11, 4.9612062016495473e-11, 4.953062697415983e-11, 
    4.9433034380671747e-11, 4.931168634668651e-11, 4.916136315267332e-11, 
    4.8979538885942192e-11, 4.8766524880866877e-11, 4.8525404524047413e-11, 
    4.826180583287447e-11, 4.7983463595954313e-11, 4.7699645437052305e-11, 
    4.7420436036427311e-11, 4.7155964020878548e-11, 4.6915605944481551e-11, 
    4.6707239192737311e-11, 4.653661193089762e-11, 4.6406882240669628e-11, 
    4.6318360538681791e-11, 4.6268514967449397e-11, 4.6252213923685907e-11, 
    4.6262214595008129e-11, 4.628983970068487e-11, 4.6325787586851132e-11, 
    4.6360995657601583e-11, 4.6387478393986196e-11, 4.6399028929620977e-11, 
    4.639175031347695e-11, 4.6364330351366104e-11, 4.6318049165778097e-11, 
    4.6256505520437739e-11, 4.6185131493976337e-11, 4.6110490909326227e-11, 
    4.6039505110360669e-11, 4.5978642751793656e-11, 4.5933192697828969e-11, 
    4.5906646221306029e-11, 4.5900311092084579e-11, 4.5913125404395425e-11, 
    4.5941718104229269e-11, 4.5980662591970855e-11, 4.6022914424045755e-11, 
    4.6060349421601688e-11, 4.6084364702036738e-11, 4.6086439980277861e-11, 
    4.6058669994727229e-11, 4.5994158760690617e-11, 4.5887310565161092e-11, 
    4.5733970369526231e-11, 4.553145585090656e-11, 4.527847951424033e-11, 
    4.4975013960534418e-11, 4.4622115848578647e-11, 4.4221745263110788e-11, 
    4.3776622827314614e-11, 4.3290108267577481e-11, 4.2766126103780727e-11, 
    4.2209141670699622e-11, 4.162412587567724e-11, 4.1016552351778205e-11, 
    4.0392361022321664e-11, 3.9757883019084743e-11, 3.9119717824713115e-11, 
    3.8484570775044679e-11, 3.785902861146464e-11, 3.724932717912991e-11, 
    3.6661133192765944e-11, 3.6099348901586415e-11, 3.5567978713528034e-11, 
    3.5070087067702129e-11, 3.4607850001663735e-11, 3.4182697951113185e-11, 
    3.3795524305670847e-11, 3.344695426021527e-11, 3.3137604753438457e-11, 
    3.2868313298566513e-11, 3.2640286179023049e-11, 3.2455134523691444e-11, 
    3.231477542104606e-11, 3.222119737032251e-11, 3.2176108929270612e-11, 
    3.2180505838421919e-11, 3.2234192617721955e-11, 3.2335335397075216e-11, 
    3.2480102878431044e-11, 3.2662455899940791e-11, 3.2874106081477346e-11, 
    3.3104709051028777e-11, 3.3342270309923414e-11, 3.3573737609566156e-11, 
    3.3785754608193216e-11, 3.3965497150171013e-11, 3.4101512147961212e-11, 
    3.4184499771723152e-11, 3.4207950591041469e-11, 3.4168587338975508e-11, 
    3.4066565059047712e-11, 3.3905428034227493e-11, 3.3691827750018817e-11, 
    3.3435048461624065e-11, 3.3146360984581052e-11, 3.2838309841054234e-11, 
    3.2523959372731622e-11, 3.2216185870423975e-11, 3.1927024079807789e-11, 
    3.1667156078354398e-11, 3.1445488830426306e-11, 3.12688891571057e-11, 
    3.114200511150749e-11, 3.1067197140304191e-11, 3.1044538996437798e-11, 
    3.1071877540038828e-11, 3.1144925270429287e-11, 3.1257410914187807e-11, 
    3.1401248349399559e-11, 3.1566772253431775e-11, 3.1743019586414033e-11, 
    3.19180943175405e-11, 3.2079578406628033e-11, 3.2215037900647567e-11, 
    3.2312558164672085e-11, 3.236132584345883e-11, 3.2352190145235378e-11, 
    3.2278191056341663e-11, 3.2134995840260947e-11, 3.1921211581986423e-11, 
    3.1638522770221821e-11, 3.1291669077344777e-11, 3.0888197487165045e-11, 
    3.0438064883787491e-11, 2.9953037826507791e-11, 2.9446013856754243e-11, 
    2.893023835545969e-11, 2.8418543692098066e-11, 2.7922609908420837e-11, 
    2.7452368977824581e-11, 2.7015536454877294e-11, 2.6617363450007441e-11, 
    2.6260560800236117e-11, 2.59454589926013e-11, 2.5670299005533281e-11, 
    2.5431709445900696e-11, 2.5225203837862138e-11, 2.5045774946664584e-11, 
    2.4888404242247126e-11, 2.4748562404991831e-11, 2.4622542886499116e-11, 
    2.4507737272483647e-11, 2.4402730636664145e-11, 2.4307320772337448e-11, 
    2.4222385474529159e-11, 2.4149728736982935e-11, 2.409180422668323e-11, 
    2.4051468058560482e-11, 2.4031675513090244e-11, 2.4035237260997525e-11, 
    2.4064532920836403e-11, 2.4121340532144114e-11, 2.4206632828558282e-11, 
    2.4320508637920695e-11, 2.4462114964646832e-11, 2.4629709565494219e-11, 
    2.4820726181565308e-11, 2.5031983511350192e-11, 2.5259876050689203e-11, 
    2.5500693487003334e-11, 2.5750860237382338e-11, 2.6007266421831824e-11, 
    2.6267462627531155e-11, 2.6529870775370191e-11, 2.6793819844840838e-11, 
    2.7059565543135908e-11, 2.7328114367314757e-11, 2.7601055660179347e-11, 
    2.7880230593007043e-11, 2.8167468073892497e-11, 2.8464226722861183e-11, 
    2.877135993413285e-11, 2.9088870673004086e-11, 2.9415816007252896e-11, 
    2.9750213646767785e-11, 3.0089111826154676e-11, 3.0428640653474838e-11, 
    3.0764178700457183e-11, 3.1090474580998209e-11, 3.1401842979112779e-11, 
    3.1692275739839986e-11, 3.1955635230053481e-11, 3.2185740024548889e-11, 
    3.2376539713456185e-11, 3.2522242747933359e-11, 3.2617504266442714e-11, 
    3.2657596676405344e-11, 3.2638677923804474e-11, 3.2557976184643725e-11, 
    3.2414084327023929e-11, 3.2207151237927473e-11, 3.1939104691882332e-11, 
    3.1613736382893666e-11, 3.1236768605373109e-11, 3.0815754164036579e-11, 
    3.0359912384803122e-11, 2.9879796491966564e-11, 2.9386919409875671e-11, 
    2.8893210688896999e-11, 2.8410489409427252e-11, 2.7949854418789751e-11, 
    2.7521136652464182e-11, 2.713236070290785e-11, 2.6789354502925616e-11, 
    2.6495439535579342e-11, 2.6251323469071977e-11, 2.6055115387502037e-11, 
    2.5902569554571156e-11, 2.5787400581610364e-11, 2.5701806878097051e-11, 
    2.5636998828138869e-11, 2.5583827182568377e-11, 2.5533341407235343e-11, 
    2.5477343640851055e-11, 2.5408777959096263e-11, 2.5322062511071982e-11, 
    2.5213240025823011e-11, 2.5080040034817799e-11, 2.4921802698264352e-11, 
    2.4739356216292821e-11, 2.4534815496922516e-11, 2.4311419257439606e-11, 
    2.4073310639314055e-11, 2.3825412218614567e-11, 2.3573262470454745e-11, 
    2.3322913832689899e-11, 2.3080772330834889e-11, 2.285342951487134e-11, 
    2.264742291372628e-11, 2.2468937897973099e-11, 2.2323403858598803e-11, 
    2.221509300020675e-11, 2.2146657849642965e-11, 2.211875192144016e-11, 
    2.2129704380063922e-11, 2.2175394371517837e-11, 2.2249275583333518e-11, 
    2.2342672286400581e-11, 2.2445265835682185e-11, 2.2545821621798724e-11, 
    2.2633026051106038e-11, 2.2696438360768134e-11, 2.2727398012618022e-11, 
    2.2719862909239667e-11, 2.2671016737771396e-11, 2.2581652710085492e-11, 
    2.2456224585363741e-11, 2.2302601751299515e-11, 2.213150166596735e-11, 
    2.195567634646099e-11, 2.1788912817459627e-11, 2.1644946155534284e-11, 
    2.1536354400915802e-11, 2.1473569792215358e-11, 2.1464043728564825e-11, 
    2.1511682349141763e-11, 2.1616526471471339e-11, 2.1774771993007553e-11, 
    2.1979031545747564e-11, 2.2218873371297441e-11, 2.2481538048714849e-11, 
    2.2752798882174076e-11, 2.3017849289265827e-11, 2.3262193829085437e-11, 
    2.3472440050198545e-11, 2.3636979915809922e-11, 2.3746456534652885e-11, 
    2.379408039464448e-11, 2.3775742765150621e-11, 2.3689967706783154e-11, 
    2.3537681317005353e-11, 2.3321926526780118e-11, 2.3047476840173643e-11, 
    2.2720460080601174e-11, 2.2347957501059327e-11, 2.1937695825489104e-11, 
    2.1497761165732883e-11, 2.1036413233544222e-11, 2.0561951330460913e-11, 
    2.008264436881642e-11, 1.9606680823333182e-11, 1.9142149184166e-11, 
    1.8696990850589732e-11, 1.8278943149418e-11, 1.7895431589430173e-11, 
    1.7553434490623309e-11, 1.7259305888405445e-11, 1.7018584293205461e-11, 
    1.6835782938235353e-11, 1.6714216263404823e-11, 1.6655823779230358e-11, 
    1.6661070774696146e-11, 1.6728867579443359e-11, 1.6856581134850649e-11, 
    1.7040067060087178e-11, 1.7273800890455527e-11, 1.7551022823156765e-11, 
    1.7863962214770909e-11, 1.8204095677083738e-11, 1.8562463021826817e-11, 
    1.8929989952246721e-11, 1.9297871489374374e-11, 1.9657935111157797e-11, 
    2.0003028115588867e-11, 2.0327339969714577e-11, 2.0626695543296436e-11, 
    2.0898741918030283e-11, 2.1143038915563982e-11, 2.1361016728627561e-11, 
    2.1555805743090333e-11, 2.1731923358731181e-11, 2.1894863749113155e-11, 
    2.2050591816331524e-11, 2.2205007218692285e-11, 2.2363380386715312e-11, 
    2.2529860698303167e-11, 2.2707056352314959e-11, 2.2895745203741938e-11, 
    2.30947093268459e-11, 2.3300746464796083e-11, 2.3508808463631633e-11, 
    2.371228283892292e-11, 2.3903366836624363e-11, 2.4073531443349153e-11, 
    2.4213984486434121e-11, 2.4316166449895651e-11, 2.4372197666440825e-11, 
    2.4375286363200376e-11, 2.4320058162973571e-11, 2.4202835459141307e-11, 
    2.4021815491438386e-11, 2.3777212396091912e-11, 2.3471293500233201e-11, 
    2.3108390233530858e-11, 2.269480242014457e-11, 2.2238670766975031e-11, 
    2.1749732258278832e-11, 2.1239022845394154e-11, 2.0718488039350358e-11, 
    2.0200533060803364e-11, 1.9697470185016852e-11, 1.9220977619914097e-11, 
    1.8781525225451346e-11, 1.8387856483801442e-11, 1.8046535162578221e-11, 
    1.7761651458818744e-11, 1.7534659217076137e-11, 1.7364420856861069e-11, 
    1.7247449441737407e-11, 1.71783398444473e-11, 1.7150311293027755e-11, 
    1.7155888896917612e-11, 1.7187589114596935e-11, 1.7238587435705731e-11, 
    1.7303244145063067e-11, 1.7377498499146562e-11, 1.7459035924461478e-11, 
    1.7547261151902116e-11, 1.7643026513994573e-11, 1.774823374744691e-11, 
    1.7865278726140795e-11, 1.7996489770232644e-11, 1.814355442343029e-11, 
    1.8307067414402468e-11, 1.848620258808986e-11, 1.8678574347512403e-11, 
    1.8880270490627664e-11, 1.9086084364944416e-11, 1.9289837999500214e-11, 
    1.948485360317694e-11, 1.9664407963595069e-11, 1.9822221693791356e-11, 
    1.9952841799929414e-11, 2.005196324205531e-11, 2.0116603335362793e-11, 
    2.0145183259057385e-11, 2.013744700134877e-11, 2.009433136188442e-11, 
    2.0017726098695373e-11, 1.9910241573088072e-11, 1.9774909831992516e-11, 
    1.9614965267349612e-11, 1.9433635958695873e-11, 1.9234031038433873e-11, 
    1.9019048992094137e-11, 1.8791396846842106e-11, 1.8553617460172014e-11, 
    1.8308188082490923e-11, 1.8057565132262975e-11, 1.7804260407200691e-11, 
    1.7550828368195817e-11, 1.7299829963248016e-11, 1.705368957831133e-11, 
    1.6814537703851269e-11, 1.6583979569765818e-11, 1.6362880538138895e-11, 
    1.6151151887247085e-11, 1.5947626781947058e-11, 1.5749983616611461e-11, 
    1.5554825618508503e-11, 1.5357836356947767e-11, 1.5154086574854101e-11, 
    1.4938382218487256e-11, 1.4705706944681418e-11, 1.4451640047947625e-11, 
    1.4172772554016286e-11, 1.3867002133119414e-11, 1.3533768378963861e-11, 
    1.3174116065667445e-11, 1.2790660546460528e-11, 1.2387416180911869e-11, 
    1.1969568786669823e-11, 1.1543140151920506e-11, 1.1114685276130003e-11, 
    1.0690993632954419e-11, 1.0278835854883686e-11, 9.8847625978802207e-12, 
    9.5149928790228238e-12, 9.1753170250889215e-12, 8.8710714297037768e-12, 
    8.6070752387769166e-12, 8.3875972433611134e-12, 8.2162265128260312e-12, 
    8.0957499122759359e-12, 8.0279507501464239e-12, 8.0134037004456018e-12, 
    8.0512628005118626e-12, 8.1391166857708337e-12, 8.2728874907024726e-12, 
    8.4468963591416049e-12, 8.6540293278692093e-12, 8.886083086819748e-12, 
    9.1342400984861449e-12, 9.3896624836787136e-12, 9.6441338428885427e-12, 
    9.8907285343084094e-12, 1.012439333283373e-11, 1.0342420316224154e-11, 
    1.054470769183954e-11, 1.0733818458025628e-11, 1.091477625752266e-11, 
    1.1094644169170986e-11, 1.1281865571131878e-11, 1.1485499102621893e-11, 
    1.1714338069904443e-11, 1.1976055244182979e-11, 1.2276411687347969e-11, 
    1.2618615421452669e-11, 1.300289548394829e-11, 1.3426290748910544e-11, 
    1.3882694120098667e-11, 1.4363130096818985e-11, 1.4856227819561989e-11, 
    1.5348855071215115e-11, 1.5826854961377217e-11, 1.6275823861410235e-11, 
    1.6681880666623654e-11, 1.7032383711012693e-11, 1.7316542350096128e-11, 
    1.7525896203081596e-11, 1.7654677417060126e-11, 1.7699981927676917e-11, 
    1.7661822955719105e-11, 1.7543018564715169e-11, 1.7348955059691067e-11, 
    1.7087241003632786e-11, 1.6767285295484082e-11, 1.6399800175749488e-11, 
    1.5996286463421642e-11, 1.5568510368755705e-11, 1.5128026967730468e-11, 
    1.4685731244344252e-11, 1.4251533776400124e-11, 1.383408878233356e-11, 
    1.34406630562103e-11, 1.3077085977458284e-11, 1.2747813559412983e-11, 
    1.2456059166174823e-11, 1.2203992897369798e-11, 1.1992952848933089e-11, 
    1.1823664154426337e-11, 1.1696416339321307e-11, 1.1611198362951486e-11, 
    1.1567752420353493e-11, 1.1565577511044638e-11, 1.1603847518702194e-11, 
    1.168130217301665e-11, 1.1796097352321878e-11, 1.1945694964383875e-11, 
    1.2126766359073516e-11, 1.2335165767538443e-11, 1.2565986484941141e-11, 
    1.2813721641192467e-11, 1.3072472565279325e-11, 1.3336267907690604e-11, 
    1.3599375360485198e-11, 1.3856649176709708e-11, 1.4103823291073489e-11, 
    1.4337744734762946e-11, 1.4556501847183658e-11, 1.4759451327410303e-11, 
    1.494712664273362e-11, 1.5121036230464767e-11, 1.528338319041064e-11, 
    1.5436750238420651e-11, 1.5583762347865317e-11, 1.5726773847527609e-11, 
    1.5867627645306275e-11, 1.6007497283395575e-11, 1.6146801225987448e-11, 
    1.6285255117537658e-11, 1.6421965581896174e-11, 1.6555571005225725e-11, 
    1.6684431387592129e-11, 1.6806790329117963e-11, 1.6920894117213354e-11, 
    1.7025065946766268e-11, 1.7117709897542273e-11, 1.7197259945312751e-11, 
    1.7262092445975477e-11, 1.7310435126485524e-11, 1.7340293115690617e-11, 
    1.7349443187867912e-11, 1.7335489244781971e-11, 1.7296027828515836e-11, 
    1.7228872995623756e-11, 1.7132352165621224e-11, 1.7005623252085238e-11, 
    1.6848954950245154e-11, 1.6663950414520832e-11, 1.6453641811138967e-11, 
    1.6222463619699601e-11, 1.5976033822450254e-11, 1.5720824672860947e-11, 
    1.5463709168497075e-11, 1.5211436632284133e-11, 1.4970118486552649e-11, 
    1.4744778246543984e-11, 1.4538985040584078e-11, 1.4354686214143166e-11, 
    1.4192190603492618e-11, 1.4050334174425787e-11, 1.3926790921220998e-11, 
    1.3818494790253831e-11, 1.372208520937999e-11, 1.3634344710186176e-11, 
    1.3552560136710494e-11, 1.3474774691396795e-11, 1.339986116425431e-11, 
    1.3327486044789643e-11, 1.3257921786800112e-11, 1.3191782042803603e-11, 
    1.3129692585306407e-11, 1.3071980134293107e-11, 1.3018413564891683e-11, 
    1.2968026896587681e-11, 1.2919050760736039e-11, 1.2868976063394881e-11, 
    1.281470049482761e-11, 1.2752776460967974e-11, 1.2679703385434096e-11, 
    1.259223773072041e-11, 1.248768298775305e-11, 1.2364140925748117e-11, 
    1.2220690661171527e-11, 1.2057502665803918e-11, 1.1875858351497656e-11, 
    1.1678113992887317e-11, 1.1467579964980902e-11, 1.1248359410994175e-11, 
    1.1025145936335541e-11, 1.080299274634163e-11, 1.0587058708388766e-11, 
    1.0382368014579658e-11, 1.0193553694348966e-11, 1.0024644588276722e-11, 
    9.8788520978506056e-12, 9.7584000215592066e-12, 9.6644115929079725e-12, 
    9.5968262610782727e-12, 9.5543670463466641e-12, 9.5345836269512371e-12, 
    9.5339267873431819e-12, 9.5478998311818249e-12, 9.5712168742840957e-12, 
    9.598032468434986e-12, 9.6221645774875903e-12, 9.637333109272165e-12, 
    9.637404624131115e-12, 9.6166167694157336e-12, 9.5697772764664495e-12, 
    9.4924635377589836e-12, 9.381172717288339e-12, 9.2334814393842096e-12, 
    9.048172082115176e-12, 8.8253594537111232e-12, 8.5665883046462064e-12, 
    8.2749216810885415e-12, 7.9549738875782104e-12, 7.6129104917316997e-12, 
    7.2563454901665234e-12, 6.8941868957363855e-12, 6.5363329571724713e-12, 
    6.1933087082890974e-12, 5.8757912337324498e-12, 5.5940855263997284e-12, 
    5.3575674037319928e-12, 5.1741698681815485e-12, 5.049930105623012e-12, 
    4.9886693067215796e-12, 4.9918341119545048e-12, 5.0585175354682658e-12, 
    5.1856348653608344e-12, 5.3682831815244639e-12, 5.6001786972271106e-12, 
    5.8741791371043231e-12, 6.182785182060574e-12, 6.5185947929633477e-12, 
    6.8746520578162703e-12, 7.2446746602867651e-12, 7.623127235533612e-12, 
    8.0051844772087497e-12, 8.3865942200061286e-12, 8.7634984204348482e-12, 
    9.1321978161904277e-12, 9.4889956812966188e-12, 9.8300715828779454e-12, 
    1.0151451270163664e-11, 1.0449041385218384e-11, 1.0718760793373143e-11, 
    1.0956703055344154e-11, 1.1159343599154063e-11, 1.1323720505315471e-11, 
    1.1447603874032306e-11, 1.1529591217863034e-11, 1.1569161905735851e-11, 
    1.1566645652353997e-11, 1.152315335322225e-11, 1.1440454714828156e-11, 
    1.1320840406747508e-11, 1.1166983047889494e-11, 1.0981814877042094e-11, 
    1.0768426470287779e-11, 1.053001956337748e-11, 1.0269873448611939e-11, 
    9.9913592306711982e-12, 9.6979628826768973e-12, 9.3933129930772501e-12, 
    9.081201665451829e-12, 8.7655895574406618e-12, 8.4505629210057904e-12, 
    8.1402826205402537e-12, 7.8388943164714024e-12, 7.550427006442577e-12, 
    7.2786752516149546e-12, 7.0271113471719845e-12, 6.798793596857137e-12, 
    6.596333106230871e-12, 6.4218788211383907e-12, 6.2771524892398254e-12, 
    6.1635023743185335e-12, 6.0819789913175465e-12, 6.0334101306542503e-12, 
    6.0184558734569715e-12, 6.0376361724233654e-12, 6.0913130466039724e-12, 
    6.1796173125873135e-12, 6.3023400464139285e-12, 6.4587753397008415e-12, 
    6.6475526212834228e-12, 6.8664587769236343e-12, 7.1122855763798831e-12, 
    7.3807458872033419e-12, 7.6664575099832733e-12, 7.962992919360448e-12, 
    8.2630724434320426e-12, 8.5588167114586287e-12, 8.8421129596720244e-12, 
    9.1050168810586389e-12, 9.3401893821781688e-12, 9.5413079180357563e-12, 
    9.7034183862049928e-12, 9.8231759613908452e-12, 9.8989716204679932e-12, 
    9.9308775151882679e-12, 9.9204674784332477e-12, 9.8704874176859705e-12, 
    9.7844369449675298e-12, 9.6660946287866655e-12, 9.5190639597407213e-12, 
    9.3463597665218188e-12, 9.1501393568790877e-12, 8.9315668457011325e-12, 
    8.6908697844910105e-12, 8.4275573334078803e-12, 8.1408142892140951e-12, 
    7.8299866765899929e-12, 7.4951359960556054e-12, 7.1376045625718068e-12, 
    6.7605133015811034e-12, 6.3691103050220048e-12, 5.9709824680900344e-12, 
    5.5760458951171774e-12, 5.1963265524347637e-12, 4.8455246830211805e-12, 
    4.5383892739217834e-12, 4.2899371811192533e-12, 4.1145682647873686e-12, 
    4.0251378823550565e-12, 4.032048996085601e-12, 4.1424106779644226e-12, 
    4.3593655615894996e-12, 4.6815977978708631e-12, 5.103093819942833e-12, 
    5.6131823409407816e-12, 6.1968779901822008e-12, 6.835475001475457e-12, 
    7.5074438732553585e-12, 8.1895155292268496e-12, 8.8579215735445099e-12, 
    9.4896947458706845e-12, 1.006393946280371e-11, 1.0562988294385266e-11, 
    1.097334522835233e-11, 1.1286350505448014e-11, 1.149852520223307e-11, 
    1.1611550461667627e-11, 1.1631938169191109e-11, 1.1570348243127531e-11, 
    1.1440704986852093e-11, 1.1259141924615645e-11, 1.1042865540822736e-11, 
    1.080904235271446e-11, 1.0573788367406565e-11, 1.0351314677725299e-11, 
    1.0153306616218219e-11, 9.988516682631011e-12, 9.8626165967464162e-12, 
    9.7782489149476848e-12, 9.7352737333708801e-12, 9.7311636000721775e-12, 
    9.7614895620804502e-12, 9.8204552576485458e-12, 9.901454801984903e-12, 
    9.9976003567365706e-12, 1.010221595057535e-11, 1.0209268068885941e-11, 
    1.0313738743556964e-11, 1.0411896039463312e-11, 1.0501505927345022e-11, 
    1.0581947085845226e-11, 1.0654223061112396e-11, 1.072087505389684e-11, 
    1.0785790101753917e-11, 1.0853899525292715e-11, 1.0930789028537193e-11, 
    1.1022224098158701e-11, 1.1133635756972153e-11, 1.126959247717429e-11, 
    1.1433307123660449e-11, 1.1626224431656781e-11, 1.1847724897509162e-11, 
    1.2094981605817576e-11, 1.2362986692004451e-11, 1.2644756768184009e-11, 
    1.2931695722730263e-11, 1.3214084587569013e-11, 1.3481677134087774e-11, 
    1.3724323576675103e-11, 1.3932596464059902e-11, 1.4098361554568206e-11, 
    1.4215261996561167e-11, 1.427906477672261e-11, 1.4287879614727725e-11, 
    1.4242238848923465e-11, 1.4145021932568115e-11, 1.400125935284311e-11, 
    1.3817831124749963e-11, 1.3603059657050268e-11, 1.3366257696325169e-11, 
    1.3117214392866398e-11, 1.2865675139261508e-11, 1.2620820937200238e-11, 
    1.2390770481912416e-11, 1.2182146936721588e-11, 1.1999716586114927e-11, 
    1.1846117070367173e-11, 1.1721702577375156e-11, 1.1624543749063885e-11, 
    1.1550530124944443e-11, 1.1493627138382816e-11, 1.1446233085431144e-11, 
    1.1399659654178367e-11, 1.1344666250995724e-11, 1.127200335656925e-11, 
    1.1172965149273788e-11, 1.1039899224946426e-11, 1.0866593689950746e-11, 
    1.0648595522622947e-11, 1.0383374728132893e-11, 1.0070372035231775e-11, 
    9.7109375434910705e-12, 9.3081617451828798e-12, 8.8666350654319028e-12, 
    8.3921969528077414e-12, 7.8916489719582299e-12, 7.3724901419653305e-12, 
    6.8426803977783531e-12, 6.3104616520545336e-12, 5.7841856465371644e-12, 
    5.2721962480261616e-12, 4.7826972786494714e-12, 4.3236512054826375e-12, 
    3.9026316943723313e-12, 3.5266766242758374e-12, 3.2020957098948042e-12, 
    2.9342828350231001e-12, 2.7274822929633653e-12, 2.5846095191448848e-12, 
    2.507053944341922e-12, 2.4945536758702334e-12, 2.5451112259964741e-12, 
    2.655005586719828e-12, 2.8188497047916675e-12, 3.029766575069391e-12, 
    3.2795978548740194e-12, 3.5592134852732816e-12, 3.8588396103185578e-12, 
    4.1684431171159652e-12, 4.478111600243229e-12, 4.7784400227982468e-12, 
    5.0608738755315462e-12, 5.3180548633644154e-12, 5.5440572519425147e-12, 
    5.7346168972993218e-12, 5.8872560934621804e-12, 6.0013313077475067e-12, 
    6.0780183280075599e-12, 6.1202164548950557e-12, 6.1323642590595127e-12, 
    6.1202117997725157e-12, 6.0905102200984619e-12, 6.0506851108761204e-12, 
    6.0084507370237281e-12, 5.9714446631731769e-12, 5.9468417634305692e-12, 
    5.9410281634335044e-12, 5.9592996643539578e-12, 6.0056320580282128e-12, 
    6.0825294064919263e-12, 6.1909495639642948e-12, 6.3303175133883825e-12, 
    6.4986205908768994e-12, 6.6925719092511976e-12, 6.9078307067030113e-12, 
    7.1392773068336899e-12, 7.3813088343445801e-12, 7.6281474099130493e-12, 
    7.8741612901134864e-12, 8.1141513135296751e-12, 8.3436168637426859e-12, 
    8.5589849240814292e-12, 8.7577604114732555e-12, 8.9386349125142514e-12, 
    9.1014887424009239e-12, 9.2473275239253273e-12, 9.3781187009737762e-12, 
    9.4965396705466757e-12, 9.605672164371183e-12, 9.7086453798772899e-12, 
    9.8082461051012262e-12, 9.9065694526341211e-12, 1.0004723225184164e-11, 
    1.0102620749746272e-11, 1.0198888815639123e-11, 1.0290922464884878e-11, 
    1.0375064432529073e-11, 1.0446902905500933e-11, 1.0501659544831154e-11, 
    1.0534636528307818e-11, 1.0541637569856926e-11, 1.0519372120242776e-11, 
    1.0465754393223399e-11, 1.0380096652383608e-11, 1.026316276501102e-11, 
    1.011709297157662e-11, 9.9451920527264135e-12, 9.7516277574980478e-12, 
    9.5410536466529067e-12, 9.3181998762334607e-12, 9.0874567446412557e-12, 
    8.852505403559947e-12, 8.6160107196651844e-12, 8.3794101294466344e-12, 
    8.1428099356327295e-12, 7.9050214732466657e-12, 7.6637200512831086e-12, 
    7.4157441632166345e-12, 7.157494977487745e-12, 6.8854444221522695e-12, 
    6.5966745937352489e-12, 6.2894347707258117e-12, 5.9636408593464619e-12, 
    5.6212815857864479e-12, 5.2666374762950127e-12, 4.9063283564149343e-12, 
    4.5491195933592217e-12, 4.205508703489503e-12, 3.8871027711598538e-12, 
    3.6058438599063923e-12, 3.3731385757023639e-12, 3.1989885293486479e-12, 
    3.0911847149145891e-12, 3.0546837048940664e-12,
  // Sqw-total(4, 0-1999)
    0.043018282567298415, 0.04298695458052211, 0.042893399044599205, 
    0.042738881910236351, 0.042525450081051561, 0.042255841647339525, 
    0.041933369288812243, 0.041561784953714556, 0.041145134968361786, 
    0.040687615008227027, 0.040193433873168941, 0.039666693830002729, 
    0.039111293549970567, 0.038530857554774187, 0.037928693794510533, 
    0.037307778719231278, 0.036670767162011057, 0.036020022682264827, 
    0.035357662836255771, 0.034685613209191779, 0.034005663969732515, 
    0.033319523154562741, 0.032628861778871622, 0.031935347089238356, 
    0.031240661701626607, 0.030546507865485188, 0.029854597535792626, 
    0.029166630201227523, 0.028484261411224222, 0.027809065595987954, 
    0.027142497041118763, 0.026485852757173425, 0.025840240507008401, 
    0.025206554490213938, 0.024585460236948624, 0.023977389257621259, 
    0.023382543061103475, 0.022800905410564679, 0.022232261218085032, 
    0.021676220323862148, 0.02113224454328904, 0.020599676721364438, 
    0.020077770994304689, 0.01956572389121412, 0.019062706193609662, 
    0.018567895524982524, 0.018080509441570435, 0.017599838379292937, 
    0.017125277278227886, 0.016656354190050383, 0.01619275381786478, 
    0.015734333859572448, 0.015281132291174645, 0.014833364333072885, 
    0.014391408718838063, 0.013955783904446356, 0.013527115858252732, 
    0.013106099900337611, 0.012693459587882629, 0.012289905799041666, 
    0.011896098945397228, 0.011512616700172769, 0.011139928872386448, 
    0.010778380218044519, 0.010428181189155276, 0.010089405985516407, 
    0.0097619968565480844, 0.0094457734157009331, 0.0091404457476640753, 
    0.0088456302453994804, 0.0085608673313678375, 0.008285640420264551, 
    0.0080193956136418582, 0.0077615616538167474, 0.0075115696110782931, 
    0.0072688716670574341, 0.0070329582375430657, 0.0068033726029945374, 
    0.0065797222282338455, 0.0063616860788762537, 0.0061490174812351747, 
    0.0059415424009883911, 0.0057391533913240707, 0.0055417998310927476, 
    0.0053494753852951328, 0.0051622038312950837, 0.0049800244783537503, 
    0.0048029783594309783, 0.0046310962063431521, 0.0044643889617999007, 
    0.0043028412737397244, 0.0041464081005114176, 0.0039950142674859456, 
    0.0038485565851394646, 0.0037069079819837549, 0.0035699230269318981, 
    0.0034374442079676904, 0.0033093083829245115, 0.0031853529055667295, 
    0.0030654210377299446, 0.0029493663705490482, 0.0028370560838656775, 
    0.0027283729667839512, 0.0026232162023340673, 0.0025215009864096275, 
    0.0024231571077799607, 0.0023281266637921257, 0.0022363611256633487, 
    0.002147817996532863, 0.0020624573218432415, 0.0019802383118637059, 
    0.0019011163177325536, 0.0018250403646216109, 0.0017519513904723056, 
    0.0016817812709403607, 0.0016144526377523893, 0.001549879426941811, 
    0.0014879680336644097, 0.0014286189082890715, 0.001371728408384891, 
    0.001317190723916543, 0.0012648997158708291, 0.001214750546288569, 
    0.0011666410231383104, 0.0011204726290966202, 0.00107615124249294, 
    0.0010335875868395202, 0.00099269746052702956, 0.00095340180108779515, 
    0.0009156266317365653, 0.0008793029257743993, 0.00084436641119935022, 
    0.0008107573270788106, 0.00077842013707583521, 0.00074730320448073968, 
    0.0007173584361785801, 0.00068854090816652155, 0.00066080849018569762, 
    0.00063412148973966567, 0.00060844233506519841, 0.00058373531236187892, 
    0.0005599663656055446, 0.00053710295902442988, 0.00051511399446096181, 
    0.00049396976977378467, 0.00047364196099718847, 0.00045410361032581698, 
    0.0004353291036969759, 0.00041729412499718867, 0.00039997557785736282, 
    0.00038335146994329184, 0.00036740075827218412, 0.00035210315741751033, 
    0.00033743891576881008, 0.00032338856857155987, 0.00030993268038419106, 
    0.00029705159360735983, 0.00028472520325703289, 0.00027293278028821369, 
    0.00026165286560596329, 0.00025086325370621265, 0.00024054107841787388, 
    0.00023066300382542878, 0.00022120551213694202, 0.00021214526853199092, 
    0.00020345953265012848, 0.00019512657906833612, 0.00018712608618957986, 
    0.00017943945509292126, 0.00017205002696730215, 0.0001649431788660799, 
    0.0001581062911540872, 0.00015152859427182639, 0.00014520091536364619, 
    0.00013911535521209808, 0.00013326493161152424, 0.00012764322627980429, 
    0.00012224406883208207, 0.00011706128401757076, 0.00011208851859788511, 
    0.00010731915339066503, 0.00010274629558678038, 9.8362837734412647e-05, 
    9.4161563684469336e-05, 9.013527878960447e-05, 8.627694178914744e-05, 
    8.257977874158639e-05, 7.903736443272767e-05, 7.5643663041648855e-05, 
    7.2393026570462732e-05, 6.9280155754422259e-05, 6.630003312488612e-05, 
    6.3447841064785123e-05, 6.0718878805019353e-05, 5.8108491364124715e-05, 
    5.5612020706282543e-05, 5.3224785372349807e-05, 5.0942090167560424e-05, 
    4.8759262863335562e-05, 4.6671710949792216e-05, 4.4674988783931265e-05, 
    4.2764864341246734e-05, 4.0937375273313914e-05, 3.9188865938108462e-05, 
    3.7516000128433551e-05, 3.5915747867048181e-05, 3.4385348297284857e-05, 
    3.2922253850749063e-05, 3.1524063105343466e-05, 3.0188450819395564e-05, 
    2.8913103488778547e-05, 2.7695667557442109e-05, 2.6533715386506234e-05, 
    2.5424731610968638e-05, 2.4366119957735775e-05, 2.335522830200752e-05, 
    2.238938795130371e-05, 2.1465962016101903e-05, 2.0582397288674341e-05, 
    1.9736274252848366e-05, 1.8925350561904266e-05, 1.8147594392505282e-05, 
    1.7401205342255594e-05, 1.6684621839701864e-05, 1.5996515256333792e-05, 
    1.5335771966168975e-05, 1.4701465432531221e-05, 1.409282098661986e-05, 
    1.3509176285742994e-05, 1.2949940507433572e-05, 1.2414555163666633e-05, 
    1.1902459039162483e-05, 1.141305921007101e-05, 1.0945709442233807e-05, 
    1.0499696565797412e-05, 1.0074234747048991e-05, 9.6684669926064328e-06, 
    9.2814727798575281e-06, 8.9122804392316348e-06, 8.5598828254570935e-06, 
    8.2232548823246026e-06, 7.9013718884846214e-06, 7.5932274129795753e-06, 
    7.2978502558680619e-06, 7.0143198539627061e-06, 6.7417797710941866e-06, 
    6.4794489612647582e-06, 6.2266305119784696e-06, 5.9827175747887629e-06, 
    5.7471962100853676e-06, 5.5196449423964947e-06, 5.2997309587164333e-06, 
    5.087203079167732e-06, 4.8818818639948831e-06, 4.6836474530602279e-06, 
    4.4924259217868105e-06, 4.3081750413522362e-06, 4.1308703303821375e-06, 
    3.9604921773957621e-06, 3.7970146201796721e-06, 3.6403961260738888e-06, 
    3.4905724736764838e-06, 3.3474516339143728e-06, 3.2109104204212161e-06, 
    3.080792636706637e-06, 2.9569084849930444e-06, 2.8390350908606633e-06, 
    2.7269181043830327e-06, 2.6202744224242431e-06, 2.5187961098833089e-06, 
    2.4221555629903817e-06, 2.330011860122763e-06, 2.2420181031236592e-06, 
    2.1578293982948281e-06, 2.0771109945811398e-06, 1.9995460207920772e-06, 
    1.9248422614479772e-06, 1.8527374893771795e-06, 1.7830030187848157e-06, 
    1.7154453333555122e-06, 1.6499058462245269e-06, 1.5862590320092733e-06, 
    1.5244093069149163e-06, 1.4642871067455683e-06, 1.4058446182696858e-06, 
    1.3490515669868603e-06, 1.2938913680619658e-06, 1.2403578308641029e-06, 
    1.1884524899254674e-06, 1.1381825357917982e-06, 1.089559246902187e-06, 
    1.0425967840535085e-06, 9.9731119783681501e-07, 9.5371951212898504e-07, 
    9.1183877308990719e-07, 8.7168498765651429e-07, 8.3327191062856503e-07, 
    7.9660967400642492e-07, 7.6170328326012265e-07, 7.2855103462152921e-07, 
    6.971429328688693e-07, 6.6745921149268351e-07, 6.3946907177307523e-07, 
    6.1312976317161277e-07, 5.8838611913801046e-07, 5.6517064052871999e-07, 
    5.4340418133215231e-07, 5.2299724396846271e-07, 5.0385183751506384e-07, 
    4.8586380125191613e-07, 4.6892545332957716e-07, 4.5292839837107426e-07, 
    4.3776631976873886e-07, 4.2333759463346003e-07, 4.0954759648779402e-07, 
    3.963105892335876e-07, 3.8355115654675376e-07, 3.712051491391559e-07, 
    3.5922016114530571e-07, 3.4755556585266077e-07, 3.3618214861704216e-07, 
    3.2508137605761742e-07, 3.142443378264286e-07, 3.0367039709134644e-07, 
    2.9336558993183405e-07, 2.833408255106908e-07, 2.7360995535262963e-07, 
    2.6418780009434348e-07, 2.5508823904864363e-07, 2.4632247887105468e-07, 
    2.3789761619548762e-07, 2.2981559514573767e-07, 2.2207263215748441e-07, 
    2.1465914219414159e-07, 2.0756015510347957e-07, 2.0075616638814495e-07, 
    1.942243271885917e-07, 1.879398509592009e-07, 1.8187750041315217e-07, 
    1.7601302080357666e-07, 1.7032440132999475e-07, 1.6479287402884836e-07, 
    1.5940359285755783e-07, 1.5414597153043515e-07, 1.4901369137430844e-07, 
    1.4400441786851288e-07, 1.3911928325223099e-07, 1.343622034273873e-07, 
    1.2973909925567741e-07, 1.252570881542114e-07, 1.2092370194848119e-07, 
    1.1674617480824727e-07, 1.1273083090119209e-07, 1.088825886487133e-07, 
    1.0520458658989057e-07, 1.0169792747998389e-07, 9.8361531295143916e-08, 
    9.5192085981551441e-08, 9.2184084963430587e-08, 8.9329943672168777e-08, 
    8.6620190609986679e-08, 8.4043732054670738e-08, 8.1588190562294249e-08, 
    7.9240316189184116e-08, 7.6986464037364861e-08, 7.481312405246658e-08, 
    7.2707478557370421e-08, 7.0657953213123599e-08, 6.8654718603468211e-08, 
    6.6690096279023321e-08, 6.4758824889399088e-08, 6.2858151400239755e-08, 
    6.0987727355706251e-08, 5.9149310508282464e-08, 5.7346293830126507e-08, 
    5.5583105183456959e-08, 5.3864536907752018e-08, 5.2195074200040187e-08, 
    5.0578291355012447e-08, 4.9016376798471438e-08, 4.7509831251290895e-08, 
    4.6057362161886369e-08, 4.4655973462990652e-08, 4.3301227646900418e-08, 
    4.1987638764080029e-08, 4.0709143877377327e-08, 3.945959641352993e-08, 
    3.8233228919180655e-08, 3.7025042413912036e-08, 3.5831093796524523e-08, 
    3.464866809414422e-08, 3.3476337444642474e-08, 3.2313920333632423e-08, 
    3.1162362788721784e-08, 3.0023566432131128e-08, 2.8900187852257292e-08, 
    2.7795429641262244e-08, 2.671283812552043e-08, 2.5656116337182252e-08, 
    2.4628955712647002e-08, 2.3634885822971344e-08, 2.2677139894905999e-08, 
    2.1758533449784623e-08, 2.0881355237902803e-08, 2.0047271540246578e-08, 
    1.9257247711928321e-08, 1.851149241639702e-08, 1.7809431261713083e-08, 
    1.7149715893780748e-08, 1.6530273250707314e-08, 1.594839653519548e-08, 
    1.5400876132451872e-08, 1.4884164379797613e-08, 1.4394564465928528e-08, 
    1.3928430331029813e-08, 1.3482362554938925e-08, 1.3053384514362783e-08, 
    1.2639084389480569e-08, 1.2237711201150435e-08, 1.1848217598083803e-08, 
    1.1470247007928292e-08, 1.1104068586185098e-08, 1.0750468322291105e-08, 
    1.0410608923225373e-08, 1.0085873315112429e-08, 9.7777073202537747e-09, 
    9.4874752500841682e-09, 9.2163393721069572e-09, 8.9651696216106765e-09, 
    8.7344857146258453e-09, 8.5244294039892525e-09, 8.3347618993641265e-09, 
    8.1648797010137449e-09, 8.013842427064386e-09, 7.880407425262785e-09, 
    7.7630684562701755e-09, 7.660097989206807e-09, 7.5695947840971938e-09, 
    7.4895391727308446e-09, 7.4178581851388112e-09, 7.352500853898816e-09, 
    7.2915215490533221e-09, 7.2331660712796077e-09, 7.175952864968092e-09, 
    7.1187398486684201e-09, 7.0607675715474634e-09, 7.0016706969755676e-09, 
    6.9414531960410661e-09, 6.880426672523409e-09, 6.8191161091598179e-09, 
    6.758141604474586e-09, 6.6980882762351265e-09, 6.6393782857901097e-09, 
    6.5821592960630762e-09, 6.5262218750538983e-09, 6.4709553812764388e-09, 
    6.4153475375847161e-09, 6.3580283315860626e-09, 6.2973541285518028e-09, 
    6.2315240845716014e-09, 6.1587177304981584e-09, 6.0772411183554682e-09, 
    5.9856682587802293e-09, 5.8829656921049857e-09, 5.7685897615592338e-09, 
    5.6425491907240734e-09, 5.5054286216140363e-09, 5.3583725104908186e-09, 
    5.2030318534987909e-09, 5.0414793281948607e-09, 4.8761003667363948e-09, 
    4.7094692595130552e-09, 4.544219494954576e-09, 4.3829173949659297e-09, 
    4.2279466049830678e-09, 4.0814095566262595e-09, 3.9450498379756378e-09, 
    3.8201976439718665e-09, 3.7077385225763676e-09, 3.6081045226962017e-09, 
    3.5212855974693884e-09, 3.4468588920018996e-09, 3.3840330690095887e-09, 
    3.3317049610472356e-09, 3.288525720677731e-09, 3.252973750303161e-09, 
    3.2234313983607633e-09, 3.1982623507646276e-09, 3.1758862703735242e-09, 
    3.1548472372756813e-09, 3.1338724034905872e-09, 3.1119178362532491e-09, 
    3.0881989244114356e-09, 3.0622038792648031e-09, 3.0336898924262976e-09, 
    3.0026629309168189e-09, 2.9693432242204635e-09, 2.9341197810668372e-09, 
    2.8974978051578819e-09, 2.8600434302633104e-09, 2.8223299903667138e-09, 
    2.784889804782646e-09, 2.7481744755984344e-09, 2.7125260308548889e-09, 
    2.6781598613535892e-09, 2.6451596666652399e-09, 2.6134833998513997e-09, 
    2.5829786306958996e-09, 2.5534049858644344e-09, 2.5244611897088753e-09, 
    2.4958139528551184e-09, 2.4671262828019576e-09, 2.4380829277831108e-09, 
    2.4084113771820458e-09, 2.377897222254462e-09, 2.3463934942463675e-09, 
    2.3138240440354573e-09, 2.2801817083050919e-09, 2.2455221972814939e-09, 
    2.2099550237794728e-09, 2.173632629682672e-09, 2.1367389269111738e-09, 
    2.0994779724741114e-09, 2.062063477553433e-09, 2.024709265268495e-09, 
    1.9876208695662936e-09, 1.9509881303189793e-09, 1.9149788671450267e-09, 
    1.8797336272506294e-09, 1.8453619052109127e-09, 1.8119401440031177e-09, 
    1.7795120924263962e-09, 1.7480918278926862e-09, 1.7176697698201283e-09, 
    1.6882214120435806e-09, 1.659718321905956e-09, 1.6321402945721874e-09, 
    1.6054874568195417e-09, 1.5797906546781253e-09, 1.5551187743951748e-09, 
    1.5315816281498863e-09, 1.5093277582917816e-09, 1.4885368656335692e-09, 
    1.469407469739876e-09, 1.4521408027856256e-09, 1.436922625709685e-09, 
    1.4239046846645703e-09, 1.4131878660379424e-09, 1.4048085830516921e-09, 
    1.3987298339051698e-09, 1.3948375575859226e-09, 1.3929426388508657e-09, 
    1.3927880630681785e-09, 1.3940605521849664e-09, 1.3964054397772251e-09, 
    1.3994436023379623e-09, 1.4027890503808728e-09, 1.4060660876091244e-09, 
    1.4089249095145418e-09, 1.4110550421551162e-09, 1.4121959083295866e-09, 
    1.412144431866845e-09, 1.4107594276792999e-09, 1.4079629806622712e-09, 
    1.4037388496206453e-09, 1.3981283303244988e-09, 1.391223801297792e-09, 
    1.3831604440010564e-09, 1.3741064947648062e-09, 1.3642526450563744e-09, 
    1.3538009328708474e-09, 1.3429538034048576e-09, 1.3319036628879767e-09, 
    1.3208235301134325e-09, 1.3098590461043621e-09, 1.2991222905573556e-09, 
    1.2886875551411315e-09, 1.2785893632126017e-09, 1.2688227002112667e-09, 
    1.2593456417866599e-09, 1.250084102668466e-09, 1.2409386692364642e-09, 
    1.2317930465006605e-09, 1.2225237566154971e-09, 1.213010345837421e-09, 
    1.2031454910959906e-09, 1.1928440860217983e-09, 1.1820506291466666e-09, 
    1.1707440798343581e-09, 1.1589398154112525e-09, 1.146688290562285e-09, 
    1.1340705849215473e-09, 1.1211911269859518e-09, 1.1081683851370171e-09, 
    1.0951243305074169e-09, 1.0821738334775381e-09, 1.0694149123059369e-09, 
    1.05692089230919e-09, 1.0447350408799343e-09, 1.032868251380046e-09, 
    1.0212997367824848e-09, 1.0099806668162157e-09, 9.9884016039141869e-10, 
    9.8779310085988787e-10, 9.7674887301911917e-10, 9.656203644043128e-10, 
    9.5433234125702505e-10, 9.4282867052551737e-10, 9.3107776834730404e-10, 
    9.1907602805939509e-10, 9.0684895896384621e-10, 8.9445012903865608e-10, 
    8.8195793065027315e-10, 8.6947059364843657e-10, 8.5709969559681624e-10, 
    8.4496278298470694e-10, 8.3317551196844674e-10, 8.2184400328365108e-10, 
    8.1105785128770838e-10, 8.0088439572956809e-10, 7.9136459238512072e-10, 
    7.8251086880875618e-10, 7.7430702774865311e-10, 7.6671026449232625e-10, 
    7.5965505734839651e-10, 7.5305863054468125e-10, 7.4682744713221228e-10, 
    7.4086428137619342e-10, 7.3507515343559656e-10, 7.2937567470284703e-10, 
    7.2369619314807279e-10, 7.1798547940979655e-10, 7.1221260749637731e-10, 
    7.0636707934676516e-10, 7.0045719884153781e-10, 6.9450699486564195e-10, 
    6.8855197571364105e-10, 6.8263421994810272e-10, 6.7679711194092505e-10, 
    6.7108032155844974e-10, 6.6551527163561061e-10, 6.601215545558891e-10, 
    6.5490443238593131e-10, 6.4985369467894205e-10, 6.4494379696916311e-10, 
    6.4013538517012028e-10, 6.3537792799796713e-10, 6.3061338994550282e-10, 
    6.2578052964769134e-10, 6.208196201145034e-10, 6.1567715902600894e-10, 
    6.1031028753674049e-10, 6.046905083376111e-10, 5.9880653009154529e-10, 
    5.9266592948802074e-10, 5.8629558678547484e-10, 5.797407486177557e-10, 
    5.7306290595607107e-10, 5.6633650068945851e-10, 5.5964481637433772e-10, 
    5.5307521028476363e-10, 5.4671416215417073e-10, 5.4064235272616709e-10, 
    5.349302319883012e-10, 5.2963425167270475e-10, 5.2479410690194619e-10, 
    5.2043101932871194e-10, 5.1654722434841348e-10, 5.1312653385545111e-10, 
    5.101359439039348e-10, 5.0752803985064671e-10, 5.0524406129359012e-10, 
    5.0321733484492831e-10, 5.0137691499075583e-10, 4.9965117075645002e-10, 
    4.9797122730036216e-10, 4.9627402716060613e-10, 4.9450500480760819e-10, 
    4.9262018850934477e-10, 4.9058774741582766e-10, 4.8838886455357105e-10, 
    4.8601797329868792e-10, 4.8348225250021788e-10, 4.8080052020475933e-10, 
    4.7800146529700294e-10, 4.7512139922854349e-10, 4.7220157625878688e-10, 
    4.6928532470425191e-10, 4.6641506785267634e-10, 4.6362952018122898e-10, 
    4.6096113996708901e-10, 4.5843407736639198e-10, 4.5606264294245701e-10, 
    4.5385046555581641e-10, 4.5179029687815542e-10, 4.498645114785212e-10, 
    4.4804619308553382e-10, 4.4630078988068246e-10, 4.4458816741598613e-10, 
    4.4286500456592366e-10, 4.4108731803602055e-10, 4.392130538637862e-10, 
    4.372045221569123e-10, 4.3503062652744358e-10, 4.3266867277804378e-10, 
    4.3010574406562453e-10, 4.2733948472965595e-10, 4.2437831046705136e-10, 
    4.2124099250138544e-10, 4.1795568351000321e-10, 4.1455841273408144e-10, 
    4.1109120829613071e-10, 4.0759991386846366e-10, 4.0413191480306694e-10, 
    4.0073383556728873e-10, 3.9744943393613667e-10, 3.9431773206058322e-10, 
    3.9137152549778513e-10, 3.8863625733515148e-10, 3.8612935289466384e-10, 
    3.8385992869189178e-10, 3.8182890334373558e-10, 3.8002939373427762e-10, 
    3.784474260353317e-10, 3.770628254567982e-10, 3.7585032530346822e-10, 
    3.7478074935868388e-10, 3.7382235224305588e-10, 3.7294217630575808e-10, 
    3.7210746106366181e-10, 3.7128700638416104e-10, 3.7045247395951992e-10, 
    3.6957952187299717e-10, 3.6864875303925712e-10, 3.6764635013341993e-10, 
    3.6656441433563696e-10, 3.6540090453510847e-10, 3.6415923249398196e-10, 
    3.6284747686572476e-10, 3.6147732585614569e-10, 3.600627721063224e-10, 
    3.586187195016553e-10, 3.5715956906005092e-10, 3.5569794624151633e-10, 
    3.5424362034945595e-10, 3.5280277905459262e-10, 3.513776515477179e-10, 
    3.4996656043026431e-10, 3.4856434005183494e-10, 3.4716314538221754e-10, 
    3.4575348140667979e-10, 3.4432543490386204e-10, 3.4286992105383847e-10, 
    3.4137985963517505e-10, 3.3985112561026828e-10, 3.382832099765586e-10, 
    3.366794736902612e-10, 3.3504701238297884e-10, 3.3339607363996147e-10, 
    3.3173915090307151e-10, 3.3008973872854944e-10, 3.2846097047639327e-10, 
    3.2686417185511601e-10, 3.2530754376848648e-10, 3.2379504456532213e-10, 
    3.2232564562449748e-10, 3.2089296090810816e-10, 3.1948538076845626e-10, 
    3.1808663331069033e-10, 3.1667679937488193e-10, 3.1523361616906452e-10, 
    3.1373406993611291e-10, 3.1215604127484277e-10, 3.1047996245494191e-10, 
    3.0869028588508318e-10, 3.0677672435773772e-10, 3.0473509053222085e-10, 
    3.0256778493290141e-10, 3.0028379315039579e-10, 2.9789830877764258e-10, 
    2.9543192178603944e-10, 2.929095199305568e-10, 2.9035888758556581e-10, 
    2.8780919490333443e-10, 2.8528937882516653e-10, 2.828266018399165e-10, 
    2.8044481473802343e-10, 2.7816358674586409e-10, 2.7599716728011246e-10, 
    2.7395396192848669e-10, 2.720363266551869e-10, 2.702407762557531e-10, 
    2.6855849617600145e-10, 2.66976197576984e-10, 2.6547713949252058e-10, 
    2.6404235433587333e-10, 2.6265186710101679e-10, 2.6128593500112876e-10, 
    2.5992613381517006e-10, 2.5855630760504354e-10, 2.5716326547254351e-10, 
    2.557372734044599e-10, 2.5427224394457778e-10, 2.5276572935066069e-10, 
    2.5121864306480274e-10, 2.4963483610190154e-10, 2.4802047715437255e-10, 
    2.4638338873421859e-10, 2.4473228043541388e-10, 2.4307603759682985e-10, 
    2.4142305002636547e-10, 2.3978066617890534e-10, 2.3815477833002434e-10, 
    2.3654962441946687e-10, 2.3496772383244492e-10, 2.3341005611618243e-10, 
    2.3187633154111513e-10, 2.3036543831395435e-10, 2.2887589008122346e-10, 
    2.2740632954530389e-10, 2.2595594269690084e-10, 2.245248040607187e-10, 
    2.2311406336694209e-10, 2.2172602890524728e-10, 2.2036406573507102e-10, 
    2.1903242694647907e-10, 2.1773595384557975e-10, 2.1647977198661424e-10, 
    2.1526893879326793e-10, 2.1410814121732822e-10, 2.1300140261108201e-10, 
    2.1195186933041005e-10, 2.1096159248842146e-10, 2.1003139397703678e-10, 
    2.0916070877512394e-10, 2.0834748405736958e-10, 2.0758804985015939e-10, 
    2.0687705900366958e-10, 2.0620743032498048e-10, 2.0557040558015689e-10, 
    2.049556585234341e-10, 2.0435156544394762e-10, 2.0374557984627112e-10, 
    2.0312475991389034e-10, 2.0247637683064411e-10, 2.0178861371086863e-10, 
    2.0105125490945066e-10, 2.0025634287563604e-10, 1.9939868253337323e-10, 
    1.984762027821408e-10, 1.9749006423500371e-10, 1.9644456611825271e-10, 
    1.9534677198472707e-10, 1.94205988793768e-10, 1.9303305665539966e-10, 
    1.9183959716055855e-10, 1.906372422143256e-10, 1.8943695709475211e-10, 
    1.8824847286570902e-10, 1.8707990902941106e-10, 1.8593756370162835e-10, 
    1.8482589396079861e-10, 1.8374760193173238e-10, 1.827038454611879e-10, 
    1.8169445807342629e-10, 1.8071820688811082e-10, 1.7977296043602383e-10, 
    1.7885587806965665e-10, 1.7796350838262083e-10, 1.7709192455708945e-10, 
    1.7623684577315268e-10, 1.7539385501121477e-10, 1.7455865653211783e-10, 
    1.7372746246260859e-10, 1.7289738192300894e-10, 1.7206686880467691e-10, 
    1.712360926097417e-10, 1.7040719652677541e-10, 1.6958433628297186e-10, 
    1.6877351493149636e-10, 1.6798209549776061e-10, 1.6721813045135861e-10, 
    1.6648942840998462e-10, 1.6580256813796741e-10, 1.6516188594737401e-10, 
    1.6456862982315241e-10, 1.6402029912821891e-10, 1.6351038767923329e-10, 
    1.6302846603571498e-10, 1.6256070949002487e-10, 1.6209074196284908e-10, 
    1.6160081806577901e-10, 1.6107313695371223e-10, 1.6049123643044767e-10, 
    1.5984126186684991e-10, 1.5911306873885144e-10, 1.5830096742441206e-10, 
    1.5740416607333363e-10, 1.5642678287380828e-10, 1.5537754776476391e-10, 
    1.5426915536122485e-10, 1.5311744712877885e-10, 1.5194040840090957e-10, 
    1.5075718359369773e-10, 1.4958707690588717e-10, 1.4844870535396365e-10, 
    1.4735924647671842e-10, 1.4633388428593146e-10, 1.4538535402821652e-10, 
    1.4452365715731858e-10, 1.4375583817078024e-10, 1.4308585279517152e-10, 
    1.4251447240595065e-10, 1.4203926266646625e-10, 1.4165458031173026e-10, 
    1.4135169619546772e-10, 1.4111898947799154e-10, 1.4094231999019747e-10, 
    1.4080551971093005e-10, 1.4069108807456957e-10, 1.4058098716457366e-10, 
    1.4045757059270562e-10, 1.4030451205519778e-10, 1.4010771641733976e-10, 
    1.3985604983817879e-10, 1.3954189916502132e-10, 1.3916141040982383e-10, 
    1.3871445510422925e-10, 1.3820424591334007e-10, 1.3763673112325899e-10, 
    1.3701973949568193e-10, 1.3636206588345056e-10, 1.3567252953500089e-10, 
    1.3495916308312677e-10, 1.3422855624759445e-10, 1.3348549184836836e-10, 
    1.3273281704722972e-10, 1.3197160801711169e-10, 1.3120151541563373e-10, 
    1.3042128813747077e-10, 1.2962932808583785e-10, 1.2882426652770917e-10, 
    1.2800537691273146e-10, 1.2717290138801732e-10, 1.2632816356447632e-10, 
    1.2547352187257915e-10, 1.2461215508760226e-10, 1.237477684161559e-10, 
    1.2288423471979421e-10, 1.2202527371884425e-10, 1.2117416316423988e-10, 
    1.2033361875491521e-10, 1.1950572507636311e-10, 1.186920599868338e-10, 
    1.1789389083256515e-10, 1.171124644129671e-10, 1.1634930911554238e-10, 
    1.15606546697722e-10, 1.1488712785966568e-10, 1.1419500304358891e-10, 
    1.1353516739349655e-10, 1.1291360985840539e-10, 1.1233714273057468e-10, 
    1.1181315958135619e-10, 1.1134930416572182e-10, 1.109531201510403e-10, 
    1.1063165914798033e-10, 1.1039111844157471e-10, 1.1023645898026802e-10, 
    1.1017108482298259e-10, 1.101965124770396e-10, 1.1031211474125026e-10, 
    1.1051485405339002e-10, 1.1079909490220852e-10, 1.1115646103767315e-10, 
    1.1157578248716196e-10, 1.120431088919275e-10, 1.1254189327076639e-10, 
    1.1305327158177355e-10, 1.1355653637653123e-10, 1.1402974188854868e-10, 
    1.144504738770139e-10, 1.1479670789062835e-10, 1.1504776775771151e-10, 
    1.1518526394133816e-10, 1.1519401408112731e-10, 1.1506280749905542e-10, 
    1.1478502703808314e-10, 1.1435900261573811e-10, 1.1378812135113951e-10, 
    1.130806423097785e-10, 1.1224925292550912e-10, 1.1131034215507065e-10, 
    1.1028311551709714e-10, 1.0918854245893381e-10, 1.0804827715249961e-10, 
    1.0688356467202894e-10, 1.0571429354222129e-10, 1.0455817699839921e-10, 
    1.0343019898048852e-10, 1.0234229223115117e-10, 1.0130331611552168e-10, 
    1.0031925466317368e-10, 9.9393671757797205e-11, 9.8528271874693413e-11, 
    9.772358950577745e-11, 9.697961843180968e-11, 9.6296413237487092e-11, 
    9.567448697592707e-11, 9.5115043807618972e-11, 9.4619977838437673e-11, 
    9.419166268251757e-11, 9.3832540837819131e-11, 9.3544611149722909e-11, 
    9.3328833334503575e-11, 9.3184587169397736e-11, 9.3109191138174777e-11, 
    9.3097623798832175e-11, 9.314240941386784e-11, 9.3233759927366495e-11, 
    9.3359902752556962e-11, 9.3507618687810699e-11, 9.3662902417193025e-11, 
    9.3811712726256335e-11, 9.3940725909472559e-11, 9.4038074039626325e-11, 
    9.4093949099747985e-11, 9.4101126361464945e-11, 9.4055291811985071e-11, 
    9.3955240210306376e-11, 9.3802871261855964e-11, 9.3603056562428803e-11, 
    9.3363324916222335e-11, 9.3093434668210913e-11, 9.2804802355133425e-11, 
    9.2509866298107426e-11, 9.2221337157435395e-11, 9.1951473677052159e-11, 
    9.171131036389935e-11, 9.1510005679574496e-11, 9.1354248534866639e-11, 
    9.1247863122573726e-11, 9.1191569381838363e-11, 9.1182983695465178e-11, 
    9.121679852836085e-11, 9.1285182622879189e-11, 9.1378291536676993e-11, 
    9.1484906438755692e-11, 9.1593069804090743e-11, 9.1690713519457327e-11, 
    9.176617135355588e-11, 9.1808603910046564e-11, 9.1808228609413118e-11, 
    9.175644796663061e-11, 9.1645828592194521e-11, 9.1470012090181637e-11, 
    9.1223565549394033e-11, 9.0901865180384854e-11, 9.0501008899189862e-11, 
    9.0017843576306599e-11, 8.9450061271710997e-11, 8.8796447996965253e-11, 
    8.8057172483061833e-11, 8.7234177615202287e-11, 8.6331538410292825e-11, 
    8.5355820036021784e-11, 8.4316281870825988e-11, 8.3224976950449085e-11, 
    8.2096615236995075e-11, 8.0948239272511538e-11, 7.9798647566365576e-11, 
    7.8667648114474569e-11, 7.7575126274835433e-11, 7.6540048910568668e-11, 
    7.5579428620455865e-11, 7.4707402724068303e-11, 7.3934418195548367e-11, 
    7.3266700894137617e-11, 7.2705967882083645e-11, 7.2249478450564018e-11, 
    7.189036395247819e-11, 7.161826261789823e-11, 7.1420145893317073e-11, 
    7.1281324786278367e-11, 7.1186487076027407e-11, 7.1120741287712665e-11, 
    7.1070546162422935e-11, 7.1024484175840369e-11, 7.0973792850482025e-11, 
    7.0912675131309497e-11, 7.0838327921257849e-11, 7.0750727909570491e-11, 
    7.0652187204809634e-11, 7.0546728754125458e-11, 7.0439327373837464e-11, 
    7.0335103532115669e-11, 7.0238514128178011e-11, 7.0152648079654755e-11, 
    7.0078650373986231e-11, 7.0015390141339274e-11, 6.9959343027679698e-11, 
    6.9904773308137517e-11, 6.9844146768673059e-11, 6.9768771683761585e-11, 
    6.9669591365519422e-11, 6.9538058900979886e-11, 6.9366972802977746e-11, 
    6.915122559042643e-11, 6.8888358302358091e-11, 6.8578875196679627e-11, 
    6.8226280083793581e-11, 6.7836858761467838e-11, 6.741920138380822e-11, 
    6.6983564551147883e-11, 6.6541111444139197e-11, 6.6103145286482731e-11, 
    6.5680357891188371e-11, 6.5282219576022149e-11, 6.491651137110449e-11, 
    6.4589038068350807e-11, 6.4303504932628738e-11, 6.4061556310849824e-11, 
    6.3862923104753584e-11, 6.3705650452802533e-11, 6.3586339482545746e-11, 
    6.3500406994592445e-11, 6.3442296318066e-11, 6.3405675340256372e-11, 
    6.3383585299249466e-11, 6.3368594683381725e-11, 6.3352951554462949e-11, 
    6.3328783272232731e-11, 6.328833626189919e-11, 6.3224281539877998e-11, 
    6.3130070968995385e-11, 6.3000324450399438e-11, 6.2831200848803113e-11, 
    6.2620737356661557e-11, 6.2369060381529523e-11, 6.2078490073575132e-11, 
    6.1753459072196046e-11, 6.1400259974788515e-11, 6.1026614888490417e-11, 
    6.064112068580257e-11, 6.0252581024444967e-11, 5.986932698324993e-11, 
    5.9498569556208609e-11, 5.9145849949894329e-11, 5.8814648617518319e-11, 
    5.8506173499895172e-11, 5.82193694485418e-11, 5.7951114148935899e-11, 
    5.7696575675063919e-11, 5.7449715879001516e-11, 5.7203843594186021e-11, 
    5.6952195911223909e-11, 5.6688474982017512e-11, 5.6407300257641404e-11, 
    5.610454536978417e-11, 5.5777554383031143e-11, 5.5425216217471231e-11, 
    5.5047934476265823e-11, 5.464748962496734e-11, 5.4226837141310921e-11, 
    5.3789870591098682e-11, 5.334117610529109e-11, 5.2885774107589128e-11, 
    5.2428911742709612e-11, 5.1975878024400849e-11, 5.1531851065650816e-11, 
    5.1101786381540392e-11, 5.0690325888855265e-11, 5.0301714604478024e-11, 
    4.9939735288140831e-11, 4.9607634682571413e-11, 4.9308045662452826e-11, 
    4.9042899454582294e-11, 4.8813339335295696e-11, 4.8619635002003036e-11, 
    4.8461124536887589e-11, 4.8336159912974936e-11, 4.8242118656687716e-11, 
    4.8175441242875828e-11, 4.8131736839241526e-11, 4.8105917787148054e-11, 
    4.8092390290542998e-11, 4.8085266510492195e-11, 4.8078593603669179e-11, 
    4.8066568763411945e-11, 4.8043733753045958e-11, 4.8005151398876892e-11, 
    4.7946524870523064e-11, 4.7864277242547926e-11, 4.7755612603499994e-11, 
    4.7618521301907804e-11, 4.7451797378589359e-11, 4.7255030769747053e-11, 
    4.7028617641045421e-11, 4.6773762478360937e-11, 4.6492499626667457e-11, 
    4.6187702546620267e-11, 4.5863095380925267e-11, 4.5523227864526431e-11, 
    4.5173430867373202e-11, 4.481971569672803e-11, 4.4468640443194777e-11, 
    4.4127112916526446e-11, 4.3802161088505883e-11, 4.3500658146764113e-11, 
    4.3229040192243829e-11, 4.299298944410733e-11, 4.2797147472629545e-11, 
    4.2644832517892416e-11, 4.2537805755849127e-11, 4.2476070397102817e-11, 
    4.2457758717594122e-11, 4.2479069319264468e-11, 4.253432394500563e-11, 
    4.2616090326252754e-11, 4.271543912163928e-11, 4.2822262966921979e-11, 
    4.292572763465783e-11, 4.3014754351164562e-11, 4.3078580466377919e-11, 
    4.3107312358317722e-11, 4.3092473793176383e-11, 4.3027471178112575e-11, 
    4.2907990341511197e-11, 4.2732231806421332e-11, 4.2501038091219022e-11, 
    4.2217825237000437e-11, 4.1888396412098423e-11, 4.1520575412179005e-11, 
    4.1123764824647615e-11, 4.0708385881914339e-11, 4.0285317448262178e-11, 
    3.9865282801956287e-11, 3.945834273067887e-11, 3.9073406078835652e-11, 
    3.8717916084196009e-11, 3.839761941825638e-11, 3.8116529229311132e-11, 
    3.7876994805298919e-11, 3.7679940053863866e-11, 3.7525173013117718e-11, 
    3.7411811768717977e-11, 3.7338676576024793e-11, 3.7304734014756374e-11, 
    3.7309412594563887e-11, 3.7352881989400484e-11, 3.7436153199074693e-11, 
    3.7561089770018457e-11, 3.7730221097307001e-11, 3.7946499046471889e-11, 
    3.8212875776064749e-11, 3.8531899873170975e-11, 3.890521077603743e-11, 
    3.9333113882595163e-11, 3.9814168450584129e-11, 4.0344912153203767e-11, 
    4.0919645649387137e-11, 4.1530409809747194e-11, 4.2167041973586359e-11, 
    4.2817414302000669e-11, 4.3467742634619049e-11, 4.4103037960113219e-11, 
    4.4707583733112025e-11, 4.5265525165367858e-11, 4.5761400498364273e-11, 
    4.6180750265591683e-11, 4.6510636115840171e-11, 4.6740157916630074e-11, 
    4.6860855122915681e-11, 4.6867084005915038e-11, 4.6756211157391784e-11, 
    4.6528783092609017e-11, 4.6188502409391918e-11, 4.5742149907787316e-11, 
    4.5199324343139877e-11, 4.457213012421544e-11, 4.3874728185244922e-11, 
    4.3122844431205669e-11, 4.2333197499293541e-11, 4.1522943140921431e-11, 
    4.0709062461287798e-11, 3.9907845082961735e-11, 3.9134368974774016e-11, 
    3.8402101192598448e-11, 3.7722537908142115e-11, 3.7104989389411685e-11, 
    3.6556408928357224e-11, 3.6081373775745337e-11, 3.5682097325857607e-11, 
    3.5358579347859738e-11, 3.5108751948845075e-11, 3.4928736658617085e-11, 
    3.4813089558559609e-11, 3.475509624988107e-11, 3.4747048932876987e-11, 
    3.4780563044822582e-11, 3.4846822648907424e-11, 3.4936876593680881e-11, 
    3.5041875211069763e-11, 3.5153333420131587e-11, 3.5263340882604582e-11, 
    3.5364801303742544e-11, 3.5451626876770012e-11, 3.5518946256324818e-11, 
    3.5563250680813478e-11, 3.5582538922935072e-11, 3.5576370400710723e-11, 
    3.5545886666977228e-11, 3.5493704098576352e-11, 3.5423747529550905e-11, 
    3.5340964141698189e-11, 3.5250968946980403e-11, 3.5159583005274546e-11, 
    3.5072376795091798e-11, 3.4994157421996112e-11, 3.4928546248512078e-11, 
    3.4877579020071116e-11, 3.484148010958335e-11, 3.481852914279562e-11, 
    3.4805138655863041e-11, 3.4796060566115812e-11, 3.4784781584365429e-11, 
    3.4763996782404755e-11, 3.4726217160789261e-11, 3.4664372566639693e-11, 
    3.4572441516929609e-11, 3.4445972127338558e-11, 3.4282541979596198e-11, 
    3.4082039137909763e-11, 3.3846802961655119e-11, 3.35815702666691e-11, 
    3.329326520848054e-11, 3.2990615986364297e-11, 3.2683666484956509e-11, 
    3.2383169894075888e-11, 3.2099957927148594e-11, 3.1844286213599479e-11, 
    3.1625242653750007e-11, 3.1450210399689824e-11, 3.1324473553151714e-11, 
    3.1250934653437786e-11, 3.1229999807455946e-11, 3.1259599156736061e-11, 
    3.1335366510324399e-11, 3.1450907953904804e-11, 3.159819485632153e-11, 
    3.1767993136793484e-11, 3.195035329821458e-11, 3.2135063733735484e-11, 
    3.2312105839662086e-11, 3.2472064928638827e-11, 3.2606484626804333e-11, 
    3.2708128533317412e-11, 3.2771206885517239e-11, 3.2791516150990454e-11, 
    3.2766524070186531e-11, 3.2695365782238275e-11, 3.2578811614727096e-11, 
    3.2419150849795268e-11, 3.2220041907041661e-11, 3.1986302133528699e-11, 
    3.1723680783834364e-11, 3.143857832625437e-11, 3.1137784272003251e-11, 
    3.0828195535189168e-11, 3.0516575124006551e-11, 3.0209330807758728e-11, 
    2.991235443914972e-11, 2.9630902414771594e-11, 2.9369541203753246e-11, 
    2.9132121367618054e-11, 2.8921810005204478e-11, 2.8741115820487277e-11, 
    2.8591941715804473e-11, 2.8475612231614205e-11, 2.8392890700257673e-11, 
    2.8343963635040799e-11, 2.8328428165136403e-11, 2.834524296139988e-11, 
    2.8392708361157302e-11, 2.8468469546465948e-11, 2.8569562342609541e-11, 
    2.8692503488533756e-11, 2.8833458004127203e-11, 2.8988459714633272e-11, 
    2.9153673406447232e-11, 2.9325681711348164e-11, 2.9501774392516095e-11, 
    2.9680173841755041e-11, 2.9860221981788985e-11, 3.0042435471923798e-11, 
    3.0228470574856324e-11, 3.0420935482576982e-11, 3.0623108935318985e-11, 
    3.0838538979557721e-11, 3.1070597399482041e-11, 3.1321982875341538e-11, 
    3.1594259700592337e-11, 3.1887454400141238e-11, 3.2199766957786489e-11, 
    3.2527390296569455e-11, 3.2864518679052405e-11, 3.3203484417956664e-11, 
    3.3535068344670326e-11, 3.3848923328594865e-11, 3.4134119435620616e-11, 
    3.4379705255748606e-11, 3.4575323418465806e-11, 3.4711776676324375e-11, 
    3.4781539400918751e-11, 3.4779152325328167e-11, 3.47015217212121e-11, 
    3.4548058191551852e-11, 3.432069966870528e-11, 3.4023788771770735e-11, 
    3.3663846650187944e-11, 3.324923108732484e-11, 3.2789752526159897e-11, 
    3.229619529171634e-11, 3.177986162910973e-11, 3.1252090956589045e-11, 
    3.0723826406370962e-11, 3.0205191691293295e-11, 2.9705169930884443e-11, 
    2.9231334977662376e-11, 2.8789683469657613e-11, 2.8384540443077344e-11, 
    2.8018591426165573e-11, 2.7692963367673163e-11, 2.7407413248474644e-11, 
    2.7160577642727782e-11, 2.6950276412251417e-11, 2.6773800781535805e-11, 
    2.6628244547262677e-11, 2.6510766479533911e-11, 2.64188349193631e-11, 
    2.635035303218073e-11, 2.6303748296905441e-11, 2.627794898357674e-11, 
    2.6272316619304182e-11, 2.6286487351628751e-11, 2.6320227462937195e-11, 
    2.637324493324449e-11, 2.6445063716346453e-11, 2.6534896211714535e-11, 
    2.6641603175221836e-11, 2.6763665445625553e-11, 2.6899231210903637e-11, 
    2.7046150788063484e-11, 2.7202049539188584e-11, 2.7364341713369299e-11, 
    2.7530268064499418e-11, 2.7696846923083565e-11, 2.7860850639105908e-11, 
    2.8018730106585674e-11, 2.8166588144862124e-11, 2.8300148462500743e-11, 
    2.841482891494866e-11, 2.8505830978703832e-11, 2.8568355512352742e-11, 
    2.8597853216491766e-11, 2.8590365195062177e-11, 2.8542834149814326e-11, 
    2.8453459179002226e-11, 2.8321961870162345e-11, 2.8149806902679098e-11, 
    2.794026125240452e-11, 2.7698364583365826e-11, 2.7430712988699893e-11, 
    2.7145133305908622e-11, 2.6850186192471617e-11, 2.6554603955516986e-11, 
    2.6266630810542495e-11, 2.5993386371738032e-11, 2.5740213125628647e-11, 
    2.551016382922913e-11, 2.530359686995885e-11, 2.5117981226489206e-11, 
    2.4947885468359042e-11, 2.4785236118740642e-11, 2.4619752339972389e-11, 
    2.4439623969450799e-11, 2.4232302462823406e-11, 2.3985432958500956e-11, 
    2.3687766744446018e-11, 2.3330074885050617e-11, 2.2905916367659383e-11, 
    2.2412265115709665e-11, 2.1849884777679713e-11, 2.1223494695743215e-11, 
    2.0541654834313319e-11, 1.9816433517231599e-11, 1.9062840024813387e-11, 
    1.829812798497279e-11, 1.7540933892221922e-11, 1.681040293747717e-11, 
    1.6125293272810109e-11, 1.5503148339154064e-11, 1.4959543633457288e-11, 
    1.4507502626037035e-11, 1.4157032903824385e-11, 1.3914857897253647e-11, 
    1.3784296164583046e-11, 1.376532156744036e-11, 1.3854727012239104e-11, 
    1.4046432147863693e-11, 1.4331853316897465e-11, 1.4700339596966345e-11, 
    1.5139623503867549e-11, 1.5636298023171529e-11, 1.6176246230466142e-11, 
    1.6745089235330715e-11, 1.7328573719971229e-11, 1.7912963215905876e-11, 
    1.8485389816452244e-11, 1.903421058787683e-11, 1.9549322597570832e-11, 
    2.0022480899935932e-11, 2.0447563314564537e-11, 2.0820795913779859e-11, 
    2.1140881753788805e-11, 2.1409034440194113e-11, 2.1628878038985338e-11, 
    2.1806200403700623e-11, 2.1948539788270659e-11, 2.2064644283122312e-11, 
    2.2163802198994952e-11, 2.2255110546501936e-11, 2.234671563283453e-11, 
    2.2445113127277299e-11, 2.2554564002119515e-11, 2.2676694653850923e-11, 
    2.2810308571638827e-11, 2.2951462982748854e-11, 2.3093788971804593e-11, 
    2.3229046661434529e-11, 2.3347844177424084e-11, 2.3440478134531214e-11, 
    2.3497784455915739e-11, 2.3511943681632592e-11, 2.3477130745070814e-11, 
    2.3389979410010101e-11, 2.3249808223343954e-11, 2.305859623656159e-11, 
    2.2820720710903657e-11, 2.2542521295615841e-11, 2.2231708916958639e-11, 
    2.1896733077190974e-11, 2.1546151282295873e-11, 2.1188079047740883e-11, 
    2.0829741972505292e-11, 2.0477208857304276e-11, 2.0135259426599916e-11, 
    1.9807407631720803e-11, 1.9496053194322594e-11, 1.9202698538695735e-11, 
    1.892820523557299e-11, 1.8673053325270697e-11, 1.843754539185942e-11, 
    1.8221964738500795e-11, 1.8026656605355992e-11, 1.7852052473617734e-11, 
    1.7698623790307861e-11, 1.7566824706299361e-11, 1.7457011039624566e-11, 
    1.7369363798881078e-11, 1.7303847172020146e-11, 1.7260189513592329e-11, 
    1.723788890977098e-11, 1.7236248032004441e-11, 1.7254426720138886e-11, 
    1.7291506672387635e-11, 1.7346533562194999e-11, 1.7418576623331012e-11, 
    1.7506770013726435e-11, 1.7610342295977193e-11, 1.7728658468223925e-11, 
    1.7861235668693766e-11, 1.8007781493812896e-11, 1.8168207505700017e-11, 
    1.8342633916776864e-11, 1.8531373859451992e-11, 1.8734878616316873e-11, 
    1.8953649499124749e-11, 1.9188100022985742e-11, 1.943837955593905e-11, 
    1.9704177643499992e-11, 1.9984526058265905e-11, 2.0277606066730887e-11, 
    2.058061755837073e-11, 2.0889721141218651e-11, 2.120005628442843e-11, 
    2.1505887496729531e-11, 2.1800830268045234e-11, 2.2078159997596007e-11, 
    2.2331188439459992e-11, 2.2553669157053549e-11, 2.2740178609237734e-11, 
    2.2886464987202094e-11, 2.2989703041288015e-11, 2.3048657259930021e-11, 
    2.30637223855807e-11, 2.303685785921294e-11, 2.2971410322459019e-11, 
    2.2871875660785465e-11, 2.274358762421495e-11, 2.2592409894632152e-11, 
    2.2424415366701145e-11, 2.2245613609843748e-11, 2.2061725092585318e-11, 
    2.1878004478777222e-11, 2.1699122695528149e-11, 2.1529119406966458e-11, 
    2.1371369821805359e-11, 2.1228593527855475e-11, 2.1102860092346217e-11, 
    2.0995632716791286e-11, 2.0907773491733231e-11, 2.0839580363809658e-11, 
    2.0790814484234304e-11, 2.0760724997600788e-11, 2.0748103882209775e-11, 
    2.0751352547098457e-11, 2.0768549180468262e-11, 2.0797556824584141e-11, 
    2.0836103899887906e-11, 2.0881876703931422e-11, 2.0932573118553401e-11, 
    2.0985946979802521e-11, 2.103979997548626e-11, 2.1091929687128599e-11, 
    2.1140052620604338e-11, 2.1181716671328906e-11, 2.1214199287984999e-11, 
    2.1234442059033976e-11, 2.1239020170291358e-11, 2.1224197928343556e-11, 
    2.1186035262016673e-11, 2.1120580471308726e-11, 2.1024118490149877e-11, 
    2.0893464298321804e-11, 2.0726246768093583e-11, 2.0521188333986249e-11, 
    2.0278296566637294e-11, 1.9998999696861179e-11, 1.9686152387472932e-11, 
    1.9343964617560035e-11, 1.8977814952000584e-11, 1.859400997852207e-11, 
    1.8199491829985326e-11, 1.7801537138608404e-11, 1.7407459695957777e-11, 
    1.7024372693612467e-11, 1.6658968705033752e-11, 1.6317356768624013e-11, 
    1.6004931659370446e-11, 1.5726257423988679e-11, 1.5484944358890383e-11, 
    1.5283524263408241e-11, 1.5123266739629762e-11, 1.5004026426806815e-11, 
    1.4924032350762746e-11, 1.487973411589337e-11, 1.4865671787638983e-11, 
    1.4874467511896925e-11, 1.4896915242877987e-11, 1.4922228989212049e-11, 
    1.4938436782023596e-11, 1.493293630221727e-11, 1.4893144524659119e-11, 
    1.4807261158984819e-11, 1.4665014932524423e-11, 1.445840554156848e-11, 
    1.4182319126475732e-11, 1.3835006130937587e-11, 1.3418342935714937e-11, 
    1.2937898338516057e-11, 1.2402738050942591e-11, 1.1825041355969885e-11, 
    1.1219505164511199e-11, 1.0602619440705767e-11, 9.9918341364319937e-12, 
    9.4046948636177682e-12, 8.8579940525333402e-12, 8.3669882996285724e-12, 
    7.9447163225528475e-12, 7.6014870130115886e-12, 7.3445085131920902e-12, 
    7.1777147127386764e-12, 7.1017596246449404e-12, 7.1141904219681389e-12, 
    7.2097529623245716e-12, 7.38084358270024e-12, 7.618027596630516e-12, 
    7.9106200875337897e-12, 8.2472900768875463e-12, 8.6166360856647565e-12, 
    9.0077254432365305e-12, 9.4105545722031545e-12, 9.8164148128972205e-12, 
    1.0218157073589553e-11, 1.0610340526831508e-11, 1.0989270653151677e-11, 
    1.1352915452518181e-11, 1.1700760478843659e-11, 1.203354881988969e-11, 
    1.235296750640934e-11, 1.2661287343192899e-11, 1.296099019480258e-11, 
    1.3254379857623493e-11, 1.3543220089535726e-11, 1.3828409113978984e-11, 
    1.4109726631148243e-11, 1.4385642227887195e-11, 1.4653232574867401e-11, 
    1.4908190648675937e-11, 1.5144950289847508e-11, 1.5356911092643123e-11, 
    1.5536778830761048e-11, 1.567697479789603e-11, 1.5770135546090563e-11, 
    1.5809639532311578e-11, 1.5790152223263306e-11, 1.5708147985273652e-11, 
    1.5562360062045824e-11, 1.5354143059436683e-11, 1.5087684412548495e-11, 
    1.4770058919797831e-11, 1.4411093244631686e-11, 1.402304029965543e-11, 
    1.3620058420567352e-11, 1.3217551294410465e-11, 1.2831360382492796e-11, 
    1.2476899352200619e-11, 1.2168294422442086e-11, 1.1917563531890664e-11, 
    1.1733937792254128e-11, 1.1623358489426912e-11, 1.158819426435169e-11, 
    1.1627203869699004e-11, 1.1735739930685423e-11, 1.1906169882370818e-11, 
    1.2128462731432982e-11, 1.2390892594144238e-11, 1.2680791839605017e-11, 
    1.2985274243628392e-11, 1.3291888022732732e-11, 1.3589151236815888e-11, 
    1.3866930721549908e-11, 1.4116692249247263e-11, 1.4331598522263913e-11, 
    1.4506523720877546e-11, 1.4637974508224567e-11, 1.472398782267474e-11, 
    1.4764027224040115e-11, 1.4758898605017397e-11, 1.4710656085306905e-11, 
    1.4622565115587393e-11, 1.4499038543454892e-11, 1.4345561399098511e-11, 
    1.4168571937502567e-11, 1.3975282270772753e-11, 1.3773410374984991e-11, 
    1.357085885524142e-11, 1.3375302864519623e-11, 1.3193764664091216e-11, 
    1.3032129448690711e-11, 1.2894720379280129e-11, 1.27839025258525e-11, 
    1.269978725540924e-11, 1.2640063060330333e-11, 1.2599979208120438e-11, 
    1.2572475517791523e-11, 1.25485115895611e-11, 1.2517541216446485e-11, 
    1.2468148016581177e-11, 1.2388784527937292e-11, 1.2268603183627756e-11, 
    1.2098288168578985e-11, 1.1870868685220479e-11, 1.1582436752802404e-11, 
    1.1232721648608721e-11, 1.0825435889641356e-11, 1.0368416149312223e-11, 
    9.8734871175567975e-12, 9.3560707233985361e-12, 8.834528243775466e-12, 
    8.3293102007046055e-12, 7.8619147634598452e-12, 7.4537597850977756e-12, 
    7.1250066479193712e-12, 6.8934438135586356e-12, 6.7734532170935874e-12, 
    6.775191491900701e-12, 6.9039756903031953e-12, 7.1599555456276553e-12, 
    7.5380826411169692e-12, 8.0283788573579459e-12, 8.6164568962632262e-12, 
    9.2843162631735068e-12, 1.0011305767846303e-11, 1.0775220334044583e-11, 
    1.155343317350632e-11, 1.2324019066124262e-11, 1.3066761500349511e-11, 
    1.3764018687926945e-11, 1.4401364649228083e-11, 1.4968015209834343e-11, 
    1.5456979995929563e-11, 1.5865009449529698e-11, 1.619230104659134e-11, 
    1.6442051608466635e-11, 1.6619896338647424e-11, 1.6733266014696856e-11, 
    1.6790737552731071e-11, 1.6801416823695364e-11, 1.6774381420833238e-11, 
    1.6718222963144932e-11, 1.6640692658481126e-11, 1.6548466363651284e-11, 
    1.6447001630845975e-11, 1.6340503819370795e-11, 1.6231984539066025e-11, 
    1.6123383401078262e-11, 1.601574662802983e-11, 1.5909462399150534e-11, 
    1.580451681413185e-11, 1.5700773956152244e-11, 1.5598260614511485e-11, 
    1.5497442703085502e-11, 1.539945710543572e-11, 1.5306308299670196e-11, 
    1.5220991470252266e-11, 1.5147524546976055e-11, 1.5090880366051723e-11, 
    1.5056800296075553e-11, 1.5051498075220691e-11, 1.5081254165628233e-11, 
    1.5151911790173077e-11, 1.526832765398033e-11, 1.5433786706709534e-11, 
    1.5649460487131546e-11, 1.5913933036455457e-11, 1.6222869720868296e-11, 
    1.6568862043315865e-11, 1.6941497504085491e-11, 1.7327663245537619e-11, 
    1.7712087636150826e-11, 1.8078114306472272e-11, 1.8408635065810992e-11, 
    1.86871489272099e-11, 1.8898840694524869e-11, 1.9031627494471988e-11, 
    1.9077044399060556e-11, 1.9030925325548619e-11, 1.8893780695391173e-11, 
    1.867088220550987e-11, 1.8371973868137309e-11, 1.801067884873643e-11, 
    1.7603616102430049e-11, 1.7169298822869191e-11, 1.6726907939580378e-11, 
    1.6295022202322258e-11, 1.5890420369358513e-11, 1.5527039149787362e-11, 
    1.5215163215871182e-11, 1.4960918465520355e-11, 1.4766085192935057e-11, 
    1.4628249480913466e-11, 1.4541242525337473e-11, 1.4495867483431053e-11, 
    1.4480782610311671e-11, 1.4483493839914719e-11, 1.4491344252751407e-11, 
    1.4492442001991016e-11, 1.4476428627324488e-11, 1.4435019332394712e-11, 
    1.4362327484644304e-11, 1.4254950358921688e-11, 1.4111819784818881e-11, 
    1.3933903005252889e-11, 1.3723778787920942e-11, 1.3485169150711438e-11, 
    1.3222498142446447e-11, 1.294049604450391e-11, 1.2643914757898204e-11, 
    1.2337363610532132e-11, 1.2025235371618923e-11, 1.1711710925252478e-11, 
    1.1400818171287103e-11, 1.1096497990891491e-11, 1.080263563894124e-11, 
    1.0523049263677505e-11, 1.0261403755358532e-11, 1.0021086278537308e-11, 
    9.8050293860170363e-12, 9.6155204710000143e-12, 9.4540448555914024e-12, 
    9.321161038629163e-12, 9.2164578863014663e-12, 9.138590972947804e-12, 
    9.0854026051121522e-12, 9.0540993728647585e-12, 9.041482804214343e-12, 
    9.0441952805049284e-12, 9.0589529656436385e-12, 9.0827383075850507e-12, 
    9.1129411882677012e-12, 9.1474414064638947e-12, 9.1846232326372842e-12, 
    9.2233416804074807e-12, 9.2628618779406891e-12, 9.3027620431747189e-12, 
    9.3428505360121523e-12, 9.383104112982276e-12, 9.4236090465440401e-12, 
    9.4645529183591333e-12, 9.5062333145843928e-12, 9.5490814144848921e-12, 
    9.5937144769346435e-12, 9.6409765384077536e-12, 9.6919856951688728e-12, 
    9.7481609205419724e-12, 9.8112360383845528e-12, 9.883240956072004e-12, 
    9.9664677436380525e-12, 1.0063396922505959e-11, 1.0176591564132839e-11, 
    1.0308571239212565e-11, 1.0461651943558666e-11, 1.0637749395288765e-11, 
    1.0838190343354407e-11, 1.1063501053483608e-11, 1.1313225654779787e-11, 
    1.1585770826287282e-11, 1.1878315593310933e-11, 1.2186779927370115e-11, 
    1.2505902869235619e-11, 1.2829395150503608e-11, 1.3150197916771716e-11, 
    1.3460825494237053e-11, 1.375376208692082e-11, 1.4021891774127006e-11, 
    1.4258935602092301e-11, 1.445983345673378e-11, 1.4621065812679139e-11, 
    1.4740853861674713e-11, 1.481924647357887e-11, 1.4858052937361145e-11, 
    1.4860638654179869e-11, 1.4831592503908086e-11, 1.4776303272886966e-11, 
    1.4700436679270332e-11, 1.4609419498182354e-11, 1.4507935135755892e-11, 
    1.439948648138034e-11, 1.4286067752743044e-11, 1.416798726883633e-11, 
    1.4043847630110754e-11, 1.3910700575835034e-11, 1.3764355815470796e-11, 
    1.3599833320298352e-11, 1.3411891053463458e-11, 1.319562055466233e-11, 
    1.294702617404727e-11, 1.2663538562387208e-11, 1.2344432377133116e-11, 
    1.1991087667901625e-11, 1.1607075611879489e-11, 1.1198064771312228e-11, 
    1.0771538052019703e-11, 1.0336360633965472e-11, 9.9022013447338374e-12, 
    9.4788961563253582e-12, 9.0757672910047746e-12, 8.7009837935415036e-12, 
    8.3610029720354514e-12, 8.0601516214729813e-12, 7.8003881061728896e-12, 
    7.5812618960177032e-12, 7.4000881096344738e-12, 7.2523114711797825e-12, 
    7.1320361792656886e-12, 7.0326634635055394e-12, 6.9475842991673238e-12, 
    6.8708464390045292e-12, 6.7977075151453328e-12, 6.7250626082423494e-12, 
    6.6516394802128686e-12, 6.5779923991646721e-12, 6.5062585070529883e-12, 
    6.4397385781655105e-12, 6.3823333588402572e-12, 6.3379362741537823e-12, 
    6.3098299981290604e-12, 6.3002049229718232e-12,
  // Sqw-total(5, 0-1999)
    0.034019537256470077, 0.034007828788687716, 0.033972748552126869, 
    0.033914432287486723, 0.033833106777954897, 0.033729089851719594, 
    0.033602788958014267, 0.033454697341395286, 0.033285387096825395, 
    0.033095498880826101, 0.032885728690369209, 0.032656812774467761, 
    0.032409512276273748, 0.032144599495737898, 0.031862847636568423, 
    0.031565025537172567, 0.031251898228248878, 0.030924233310712628, 
    0.030582812245065424, 0.03022844483694764, 0.0298619846269477, 
    0.02948434263938091, 0.029096497053264093, 0.028699496808703297, 
    0.028294457881000778, 0.027882551834227901, 0.027464987180911882, 
    0.027042984904165051, 0.026617750143416597, 0.026190442437220973, 
    0.025762147025226143, 0.025333849540626209, 0.024906416009403163, 
    0.02448057947266542, 0.024056933839487888, 0.02363593484520091, 
    0.023217907320651782, 0.022803057450727127, 0.022391488377606312, 
    0.021983217422001208, 0.021578193356716516, 0.021176312537158189, 
    0.020777433204462337, 0.020381387835085106, 0.019987993912237514, 
    0.019597063844417943, 0.019208414886744164, 0.018821879805936848, 
    0.018437318692392173, 0.018054631831233431, 0.017673773000068334, 
    0.01729476207925916, 0.016917695545993122, 0.016542753350563336, 
    0.016170200870300067, 0.015800385080267015, 0.015433724700186495, 
    0.015070694771621965, 0.014711806773445473, 0.0143575858920166, 
    0.014008547349129792, 0.013665173721050245, 0.013327894966700036, 
    0.012997072473525684, 0.012672987904960907, 0.012355837084039803, 
    0.012045728657578548, 0.011742686917440317, 0.011446657942593964, 
    0.011157518168466447, 0.010875084560844926, 0.010599125723999247, 
    0.01032937345372298, 0.010065534407738738, 0.009807301674885506, 
    0.0095543660666708458, 0.0093064269357482372, 0.0090632022669127708, 
    0.0088244377171059745, 0.008589914232060061, 0.0083594538622672725, 
    0.0081329234520512682, 0.0079102359814308063, 0.007691349488089849, 
    0.007476263664946076, 0.0072650143935141971, 0.0070576666127006565, 
    0.0068543060212474666, 0.0066550301623630424, 0.0064599394419112789, 
    0.0062691285940026532, 0.006082679040651507, 0.0059006525066380025, 
    0.0057230861564247807, 0.0055499894235061156, 0.0053813426074613155, 
    0.0052170972216575807, 0.0050571779857175245, 0.0049014862729046512, 
    0.0047499047464001579, 0.0046023028546160211, 0.0044585428098219112, 
    0.0043184856519432827, 0.0041819970044602497, 0.0040489521633395179, 
    0.0039192402210590262, 0.0037927670109242566, 0.0036694567542071917, 
    0.0035492523946673263, 0.0034321147018707122, 0.0033180203074623859, 
    0.0032069589002503285, 0.0030989298424912203, 0.002993938480128321, 
    0.0028919924059640223, 0.0027930979014877161, 0.0026972567367491477, 
    0.0026044634555140661, 0.0025147032219310361, 0.0024279502607810807, 
    0.0023441668897046597, 0.0022633031197500843, 0.0021852967888227322, 
    0.0021100741878242115, 0.0020375511370325965, 0.0019676344662007753, 
    0.0019002238426813773, 0.0018352138763997046, 0.0017724964099007868, 
    0.0017119628795225609, 0.0016535066151115046, 0.0015970249362003805, 
    0.0015424209069544875, 0.0014896046331634792, 0.0014384940219128121, 
    0.001389014974980966, 0.0013411010443834612, 0.0012946926349610966, 
    0.0012497358862042414, 0.0012061813964140641, 0.0011639829619897273, 
    0.0011230964915291627, 0.0010834792205000777, 0.0010450893026386773, 
    0.001007885796405732, 0.00097182900724435497, 0.00093688109713728853, 
    0.00090300683853856685, 0.00087017437410031879, 0.00083835584772125381, 
    0.00080752779440401538, 0.00077767121197279529, 0.00074877128109683154, 
    0.00072081674500082545, 0.00069379900084758138, 0.00066771098638118698, 
    0.0006425459650254942, 0.00061829631911652818, 0.00059495245492613706, 
    0.0005725019066504471, 0.00055092870257577523, 0.00053021302862743178, 
    0.00051033119584097987, 0.00049125589194616657, 0.0004729566755095216, 
    0.00045540065543067616, 0.00043855328968593263, 0.00042237923498092395, 
    0.00040684318271855952, 0.0003919106252869935, 0.00037754850873810515, 
    0.00036372574198417231, 0.00035041354725299075, 0.00033758565043576124, 
    0.00032521832209369514, 0.00031329028950664606, 0.00030178254679878285, 
    0.00029067809372190892, 0.0002799616342430639, 0.00026961926403345999, 
    0.00025963817181394558, 0.00025000637391058136, 0.00024071249497257155, 
    0.00023174560124953337, 0.00022309508668811852, 0.00021475060687272101, 
    0.000206702051862591, 0.00019893954650974894, 0.00019145346597829608, 
    0.00018423445488996676, 0.00017727344060304462, 0.00017056163426682744, 
    0.00016409051702699653, 0.000157851812558731, 0.00015183745041927224, 
    0.00014603952704998131, 0.00014045027226306347, 0.00013506202857658256, 
    0.00012986724890600874, 0.00012485851521662421, 0.00012002857730219618, 
    0.00011537040749490699, 0.00011087726441857372, 0.00010654275733887229, 
    0.00010236090248691458, 9.8326163931573171e-05, 9.4433473892220789e-05, 
    9.0678230372471548e-05, 8.7056273108619326e-05, 8.3563841531108265e-05, 
    8.0197520305171226e-05, 7.6954178808270391e-05, 7.3830910587196821e-05, 
    7.0824977594883786e-05, 6.7933762162948125e-05, 6.5154727629731431e-05, 
    6.2485386714738108e-05, 5.9923275433541794e-05, 5.7465929771228358e-05, 
    5.5110862516791305e-05, 5.2855538495128582e-05, 5.0697347699789139e-05, 
    4.8633577243916139e-05, 4.6661384322926246e-05, 4.4777773273325128e-05, 
    4.2979580156496936e-05, 4.1263468030484893e-05, 3.9625935239931053e-05, 
    3.8063337782442375e-05, 3.6571925293381052e-05, 3.5147888649299587e-05, 
    3.3787415842774739e-05, 3.2486751806988077e-05, 3.1242257394049173e-05, 
    3.0050462786659928e-05, 2.8908111230194331e-05, 2.7812190021009423e-05, 
    2.6759947040000473e-05, 2.5748892605168498e-05, 2.477678785717259e-05, 
    2.3841622121852634e-05, 2.2941582586071842e-05, 2.2075020093992179e-05, 
    2.1240414895434428e-05, 2.0436345781200384e-05, 1.9661465299933102e-05, 
    1.8914482775324477e-05, 1.8194155763677498e-05, 1.7499289540100754e-05, 
    1.6828743297464308e-05, 1.6181441073932084e-05, 1.5556385048166676e-05, 
    1.4952668767495269e-05, 1.4369488080216064e-05, 1.3806147971221896e-05, 
    1.3262064076379947e-05, 1.2736758290890565e-05, 1.2229848515156825e-05, 
    1.1741033134377601e-05, 1.127007126633725e-05, 1.0816760115103158e-05, 
    1.0380910939057378e-05, 9.9623251912950282e-06, 9.5607723403731562e-06, 
    9.1759707458321133e-06, 8.8075727620306773e-06, 8.4551549818065355e-06, 
    8.1182142157116102e-06, 7.7961694378326012e-06, 7.4883695302485825e-06, 
    7.1941062451939273e-06, 6.9126314115626952e-06, 6.6431770774016435e-06, 
    6.3849770457320367e-06, 6.1372881587568088e-06, 5.8994097379286334e-06, 
    5.6706997922753347e-06, 5.45058694591912e-06, 5.2385774650191243e-06, 
    5.0342572329969918e-06, 4.8372889709687718e-06, 4.6474053775873946e-06, 
    4.4643991289075257e-06, 4.2881108174804068e-06, 4.1184159206268929e-06, 
    3.9552117927922547e-06, 3.7984055059319911e-06, 3.6479031542453859e-06, 
    3.5036010266272397e-06, 3.3653788601787099e-06, 3.2330952325271193e-06, 
    3.1065850351297892e-06, 2.9856588863636992e-06, 2.8701042845860699e-06, 
    2.759688255618624e-06, 2.6541612121925948e-06, 2.5532617113107903e-06, 
    2.4567217742545755e-06, 2.3642724264801094e-06, 2.2756491280313883e-06, 
    2.1905967993336003e-06, 2.108874202298907e-06, 2.0302575041852218e-06, 
    1.9545429242477249e-06, 1.8815484295305934e-06, 1.8111145005081444e-06, 
    1.7431040243004693e-06, 1.6774013959088555e-06, 1.6139109194248652e-06, 
    1.5525546104417091e-06, 1.493269512338628e-06, 1.4360046585568289e-06, 
    1.380717837805512e-06, 1.3273723463049988e-06, 1.2759339307178905e-06, 
    1.2263681298823124e-06, 1.1786382036728133e-06, 1.132703791389195e-06, 
    1.0885203705856562e-06, 1.0460394996948415e-06, 1.0052097348164242e-06, 
    9.6597802943579609e-07, 9.2829136754622348e-07, 8.9209835839813108e-07, 
    8.5735053767499936e-07, 8.2400317515514123e-07, 7.9201547224540811e-07, 
    7.6135013233716949e-07, 7.3197238455932489e-07, 7.0384862329368964e-07, 
    6.7694487748699046e-07, 6.5122534016543509e-07, 6.2665116749577152e-07, 
    6.031797058013915e-07, 5.8076423310225813e-07, 5.593542241203374e-07, 
    5.3889607577892132e-07, 5.193341766025995e-07, 5.0061217292158976e-07, 
    4.8267428076075548e-07, 4.6546650972463943e-07, 4.4893769917911334e-07, 
    4.3304030731768497e-07, 4.1773093368491901e-07, 4.0297058722474704e-07, 
    3.8872473305813374e-07, 3.7496315975672477e-07, 3.6165970886320331e-07, 
    3.4879190204414016e-07, 3.3634049438717373e-07, 3.2428897713118221e-07, 
    3.1262305265976583e-07, 3.0133010763652247e-07, 2.9039871610307973e-07, 
    2.7981820897146191e-07, 2.6957834794676244e-07, 2.596691366588085e-07, 
    2.5008079028214814e-07, 2.4080386632041417e-07, 2.3182953778160981e-07, 
    2.2314996737528705e-07, 2.1475872340459174e-07, 2.0665116641148046e-07, 
    1.9882473445206527e-07, 1.9127906292914455e-07, 1.8401589304872312e-07, 
    1.7703874681485486e-07, 1.7035237437139615e-07, 1.6396200612825542e-07, 
    1.5787246570779997e-07, 1.5208721633396603e-07, 1.466074229268594e-07, 
    1.4143111307052643e-07, 1.3655251414025206e-07, 1.3196163063159216e-07, 
    1.2764410827846851e-07, 1.2358140920976684e-07, 1.1975129873770198e-07, 
    1.161286188946858e-07, 1.1268630011774974e-07, 1.0939654063771867e-07, 
    1.0623206699511262e-07, 1.0316737894515309e-07, 1.0017988113530865e-07, 
    9.7250811593355094e-08, 9.436589465244101e-08, 9.1515670428973302e-08, 
    8.8695483568622872e-08, 8.5905145364759026e-08, 8.3148313599432903e-08, 
    8.043165818135909e-08, 7.776389671282022e-08, 7.5154789276111607e-08, 
    7.2614177559445685e-08, 7.0151139655283791e-08, 6.7773312606650027e-08, 
    6.5486411723822135e-08, 6.3293953699499686e-08, 6.1197171125295205e-08, 
    5.9195092414381545e-08, 5.7284753090243622e-08, 5.5461502769346021e-08, 
    5.3719374440927196e-08, 5.2051488345321844e-08, 5.0450468483814442e-08, 
    4.8908855331449241e-08, 4.7419501107046562e-08, 4.5975935182069385e-08, 
    4.4572685920861656e-08, 4.3205543834254052e-08, 4.1871749304312834e-08, 
    4.0570088980885011e-08, 3.9300887623735511e-08, 3.8065888348069173e-08, 
    3.6868022291148898e-08, 3.5711078956154507e-08, 3.4599298328688442e-08, 
    3.3536915173079854e-08, 3.2527691995598294e-08, 3.157448042295132e-08, 
    3.0678849168971838e-08, 2.9840811921165885e-08, 2.9058679300246799e-08, 
    2.8329048136017759e-08, 2.7646928204279051e-08, 2.7005994349741127e-08, 
    2.6398940256850096e-08, 2.581790177739485e-08, 2.5254911999353004e-08, 
    2.4702349203897504e-08, 2.4153340929445521e-08, 2.3602093947330229e-08, 
    2.3044128509273006e-08, 2.2476406287717785e-08, 2.1897352266239327e-08, 
    2.1306781539985979e-08, 2.0705749740801612e-08, 2.0096351467325957e-08, 
    1.9481492439327428e-08, 1.8864659633830024e-08, 1.8249708651179158e-08, 
    1.7640681116924557e-08, 1.7041656959439253e-08, 1.6456639587772977e-08, 
    1.5889466030153917e-08, 1.5343731170998004e-08, 1.4822714412218281e-08, 
    1.4329299526331769e-08, 1.3865882472214501e-08, 1.3434267714911162e-08, 
    1.3035559091441215e-08, 1.2670056455216629e-08, 1.233717233968513e-08, 
    1.2035384147322918e-08, 1.1762235656845276e-08, 1.1514398040587055e-08, 
    1.1287794662677702e-08, 1.1077787389367032e-08, 1.0879414702874675e-08, 
    1.0687665893460385e-08, 1.0497770332122449e-08, 1.0305478402835079e-08, 
    1.0107310225805867e-08, 9.900750964467693e-09, 9.6843760418898059e-09, 
    9.4578964287475698e-09, 9.2221214149499864e-09, 8.9788442590986787e-09, 
    8.7306626046816972e-09, 8.4807511635944529e-09, 8.2326069881822977e-09, 
    7.9897887995374948e-09, 7.7556701443465564e-09, 7.5332231926313613e-09, 
    7.3248452521362731e-09, 7.1322353209529179e-09, 6.9563228932186268e-09, 
    6.7972473292675044e-09, 6.6543827842690464e-09, 6.5264020291606179e-09, 
    6.4113714648108347e-09, 6.3068699374876257e-09, 6.2101241911793361e-09, 
    6.1181547861208311e-09, 6.0279264807923533e-09, 5.9364976895567414e-09, 
    5.8411632526971207e-09, 5.7395848407088754e-09, 5.6299028988852553e-09, 
    5.5108244715486e-09, 5.3816814913431769e-09, 5.2424556951246946e-09, 
    5.0937677303270721e-09, 4.9368305636720833e-09, 4.7733694948675332e-09, 
    4.6055137625762709e-09, 4.4356666180632717e-09, 4.2663625969303432e-09, 
    4.1001213333931698e-09, 3.9393075488503697e-09, 3.7860060206359074e-09, 
    3.6419191514502039e-09, 3.508292730803965e-09, 3.3858735623536818e-09, 
    3.2749000923877157e-09, 3.1751252511972092e-09, 3.0858684202987158e-09, 
    3.0060919038591045e-09, 2.9344957484075148e-09, 2.8696239616629111e-09, 
    2.8099744708050782e-09, 2.7541053210174247e-09, 2.7007298267195526e-09, 
    2.6487944921528296e-09, 2.5975346460009859e-09, 2.5465045918853099e-09, 
    2.4955808532640159e-09, 2.4449393390549304e-09, 2.395009063172245e-09, 
    2.346407069820857e-09, 2.2998604393867732e-09, 2.2561223065763512e-09, 
    2.2158890284254947e-09, 2.1797254079949596e-09, 2.1480038631580162e-09, 
    2.1208621828059727e-09, 2.0981826095063958e-09, 2.0795932360177687e-09, 
    2.0644906211581427e-09, 2.0520810336621913e-09, 2.0414361443855169e-09, 
    2.0315582437816414e-09, 2.0214494022598257e-09, 2.0101792503220511e-09, 
    1.9969462675817134e-09, 1.9811285180080459e-09, 1.9623206179065272e-09, 
    1.9403550947015705e-09, 1.9153073286088348e-09, 1.887484618515751e-09, 
    1.857400755452577e-09, 1.82573848134033e-09, 1.7933026972083935e-09, 
    1.7609678646535611e-09, 1.7296230312503546e-09, 1.7001180754594073e-09, 
    1.6732142841652259e-09, 1.6495421832534642e-09, 1.6295687372974071e-09, 
    1.6135754493939226e-09, 1.6016480198798357e-09, 1.5936775446814111e-09, 
    1.58937237860227e-09, 1.5882793042928558e-09, 1.5898120598665431e-09, 
    1.5932851455054423e-09, 1.5979506077405072e-09, 1.6030357523632039e-09, 
    1.6077797892657038e-09, 1.6114679014704454e-09, 1.6134613693699076e-09, 
    1.6132228992572301e-09, 1.6103364020584529e-09, 1.6045208144477531e-09, 
    1.5956375796530813e-09, 1.5836917483440707e-09, 1.5688266250051354e-09, 
    1.5513122314156366e-09, 1.5315280057558478e-09, 1.5099405855545078e-09, 
    1.4870776816814739e-09, 1.463499528772138e-09, 1.4397694657260616e-09, 
    1.4164254746257314e-09, 1.393954334849397e-09, 1.3727699926508979e-09, 
    1.3531973240528176e-09, 1.3354621149408881e-09, 1.3196874568205198e-09, 
    1.305896443907969e-09, 1.2940203823025735e-09, 1.2839115871217802e-09, 
    1.2753594134468346e-09, 1.2681082879168402e-09, 1.2618763093469121e-09, 
    1.2563733868136712e-09, 1.2513178341138881e-09, 1.2464508073090405e-09, 
    1.241548015423383e-09, 1.2364285245422914e-09, 1.2309604406250952e-09, 
    1.2250636016123893e-09, 1.2187092376597292e-09, 1.2119168747973086e-09, 
    1.2047485708924578e-09, 1.1973008468827372e-09, 1.1896946102453305e-09, 
    1.1820636163940686e-09, 1.1745420176829214e-09, 1.1672518388807295e-09, 
    1.1602911263794774e-09, 1.1537237688119942e-09, 1.1475717598133539e-09, 
    1.1418107023175012e-09, 1.1363689955232888e-09, 1.1311309843774909e-09, 
    1.1259438380052772e-09, 1.1206277349132995e-09, 1.1149884196227253e-09, 
    1.1088311250612665e-09, 1.1019745392121345e-09, 1.0942636476060564e-09, 
    1.0855802235460476e-09, 1.0758502171648024e-09, 1.0650473895945089e-09, 
    1.0531931486393011e-09, 1.0403527234954237e-09, 1.0266283878787053e-09, 
    1.0121504585402289e-09, 9.9706718943452801e-10, 9.8153447984837316e-10, 
    9.6570645387418733e-10, 9.4972757061795367e-10, 9.3372688685734279e-10, 
    9.178146306399731e-10, 9.0208113297950117e-10, 8.865977574012181e-10, 
    8.7141948620029227e-10, 8.5658847037951734e-10, 8.4213809835820433e-10, 
    8.28096865926304e-10, 8.1449173182317214e-10, 8.0135047840844949e-10, 
    7.8870300943612663e-10, 7.7658145355178841e-10, 7.650192573072129e-10, 
    7.5404936717900928e-10, 7.4370191724683831e-10, 7.3400157295867824e-10, 
    7.2496501438813363e-10, 7.1659868422629798e-10, 7.0889714530930382e-10, 
    7.0184208800323856e-10, 6.9540216025241024e-10, 6.8953350604386316e-10, 
    6.841810642517654e-10, 6.7928039099742796e-10, 6.7476000855737933e-10, 
    6.7054401362026878e-10, 6.6655492176896104e-10, 6.627165623388311e-10, 
    6.5895697489235716e-10, 6.5521111273916769e-10, 6.5142337906577867e-10, 
    6.4754972679991256e-10, 6.4355932305989594e-10, 6.3943547465719115e-10, 
    6.3517583382342722e-10, 6.3079163514160649e-10, 6.2630602230660155e-10, 
    6.2175139556312405e-10, 6.1716603575538016e-10, 6.1259012082477555e-10, 
    6.0806159243888002e-10, 6.0361213917335195e-10, 5.9926383163997951e-10, 
    5.9502665508338565e-10, 5.9089733391969459e-10, 5.8685951271363493e-10, 
    5.8288538874488265e-10, 5.7893854462704918e-10, 5.7497780255594863e-10, 
    5.709615978876891e-10, 5.6685251808477167e-10, 5.6262145135615208e-10, 
    5.5825103806185553e-10, 5.5373797748217966e-10, 5.4909412071455683e-10, 
    5.4434610997563087e-10, 5.3953376044926981e-10, 5.3470721406409043e-10, 
    5.2992322419125307e-10, 5.2524076678556441e-10, 5.2071645067697531e-10, 
    5.1639998498322905e-10, 5.1233011977243491e-10, 5.0853130482441894e-10, 
    5.0501140429553572e-10, 5.0176052814308614e-10, 4.9875122468572341e-10, 
    4.959398966773403e-10, 4.9326948681911273e-10, 4.906731252421173e-10, 
    4.8807860163171209e-10, 4.8541323526835416e-10, 4.8260886355107928e-10, 
    4.7960648457388372e-10, 4.7636029998915917e-10, 4.7284073677106768e-10, 
    4.6903632573172266e-10, 4.649542007150712e-10, 4.6061928652846871e-10, 
    4.5607218497284487e-10, 4.513660338160148e-10, 4.4656253781829733e-10, 
    4.4172761551475414e-10, 4.3692692316654105e-10, 4.3222173609013896e-10, 
    4.2766540702558777e-10, 4.2330074622765213e-10, 4.1915839809561737e-10, 
    4.152563727859144e-10, 4.1160057991423937e-10, 4.0818636218862791e-10, 
    4.0500068685836061e-10, 4.0202488676820539e-10, 3.992375579137869e-10, 
    3.9661744178862695e-10, 3.9414595422055128e-10, 3.918092551155622e-10, 
    3.8959961320084347e-10, 3.875160675275787e-10, 3.8556423600331188e-10, 
    3.8375543704088655e-10, 3.821050925422743e-10, 3.8063065287165335e-10, 
    3.7934913001400798e-10, 3.7827457145933635e-10, 3.7741560078696487e-10, 
    3.7677335589410985e-10, 3.763399434231692e-10, 3.76097670046809e-10, 
    3.7601903924497091e-10, 3.7606765712395732e-10, 3.7619984779975702e-10, 
    3.7636697209169121e-10, 3.7651811572375619e-10, 3.7660300247071725e-10, 
    3.76574785572416e-10, 3.763925565929051e-10, 3.7602328148446349e-10, 
    3.7544314167188011e-10, 3.7463811823573388e-10, 3.736039497632942e-10, 
    3.7234544416621811e-10, 3.7087538634012201e-10, 3.6921311201783701e-10, 
    3.6738297654173954e-10, 3.6541278994555508e-10, 3.63332392984085e-10, 
    3.6117235190867545e-10, 3.5896288073806971e-10, 3.5673289935265741e-10, 
    3.5450927060224012e-10, 3.5231612496464396e-10, 3.5017430617008548e-10, 
    3.4810085195186876e-10, 3.4610862516287086e-10, 3.4420599784598302e-10, 
    3.4239673621283797e-10, 3.4068001971922041e-10, 3.3905071503795737e-10, 
    3.3749981584449916e-10, 3.3601512340392021e-10, 3.3458205304575809e-10, 
    3.3318459381175772e-10, 3.3180625277527678e-10, 3.3043101992031553e-10, 
    3.2904420194690304e-10, 3.2763313980332909e-10, 3.2618769111122237e-10, 
    3.2470056434650577e-10, 3.2316741662633174e-10, 3.215868076373286e-10, 
    3.1995999609112901e-10, 3.1829066542235781e-10, 3.1658456409123138e-10, 
    3.1484917702265905e-10, 3.1309335187970547e-10, 3.1132699544210969e-10, 
    3.0956075567529657e-10, 3.0780574179153614e-10, 3.0607319781507334e-10, 
    3.0437417265520739e-10, 3.0271910295393821e-10, 3.0111735996372582e-10, 
    2.9957670362639883e-10, 2.981027349613087e-10, 2.9669828868379202e-10, 
    2.953629438260893e-10, 2.940925927374108e-10, 2.9287923109244374e-10, 
    2.9171095181334184e-10, 2.9057224743943678e-10, 2.8944456964753728e-10, 
    2.8830721805614064e-10, 2.8713840552744431e-10, 2.8591654000915759e-10, 
    2.8462151884262056e-10, 2.832360125910331e-10, 2.8174655024318523e-10, 
    2.8014436960176646e-10, 2.7842588255848058e-10, 2.7659279061827883e-10, 
    2.7465175296507861e-10, 2.7261372473320918e-10, 2.7049295457564331e-10, 
    2.6830581338728607e-10, 2.6606949551008141e-10, 2.6380078869349052e-10, 
    2.6151497211076937e-10, 2.5922498130151515e-10, 2.5694087787445518e-10, 
    2.5466969998524823e-10, 2.5241564577893616e-10, 2.5018060524333949e-10, 
    2.4796491709070486e-10, 2.457683162711176e-10, 2.4359089597542352e-10, 
    2.4143404972888614e-10, 2.3930120897778907e-10, 2.3719836456578531e-10, 
    2.3513424537603319e-10, 2.3312019040540989e-10, 2.3116965409243209e-10, 
    2.2929745296485516e-10, 2.2751876806121312e-10, 2.2584804539374692e-10, 
    2.2429785632504025e-10, 2.2287786511827417e-10, 2.2159398271343285e-10, 
    2.2044779953929002e-10, 2.194363207999129e-10, 2.1855208657783763e-10, 
    2.1778357748100073e-10, 2.1711593788151738e-10, 2.1653188226630585e-10, 
    2.1601273701277046e-10, 2.1553947553640866e-10, 2.1509370839512699e-10, 
    2.146584751561286e-10, 2.142188622867279e-10, 2.1376235320862715e-10, 
    2.1327896352479989e-10, 2.1276114578848594e-10, 2.1220355669341704e-10, 
    2.1160271094568351e-10, 2.1095661763519214e-10, 2.1026441779730902e-10, 
    2.0952610059200949e-10, 2.0874229614325564e-10, 2.0791417302083423e-10, 
    2.0704338660586993e-10, 2.0613211098651507e-10, 2.0518306740140555e-10, 
    2.0419956852599452e-10, 2.0318551449815524e-10, 2.0214536826392051e-10, 
    2.010840596357228e-10, 2.0000686850958833e-10, 1.9891927030192431e-10, 
    1.9782677945535061e-10, 1.9673478007625765e-10, 1.9564839581305927e-10, 
    1.9457236499534971e-10, 1.9351097407672438e-10, 1.9246798681561699e-10, 
    1.9144664281280727e-10, 1.9044964400214589e-10, 1.8947919437835367e-10, 
    1.885370216642042e-10, 1.8762443669282324e-10, 1.8674236778244562e-10, 
    1.8589141761302048e-10, 1.8507187048623346e-10, 1.8428370931270503e-10, 
    1.8352657873075256e-10, 1.8279973404893522e-10, 1.8210192166005437e-10, 
    1.8143125549841255e-10, 1.8078503994299168e-10, 1.8015960985610107e-10, 
    1.7955014369342238e-10, 1.7895053655790407e-10, 1.7835331519584583e-10, 
    1.7774964574761478e-10, 1.7712940832756948e-10, 1.7648142027989273e-10, 
    1.7579374418889293e-10, 1.7505413597527378e-10, 1.7425055367389747e-10, 
    1.7337177737040533e-10, 1.7240803736121633e-10, 1.7135167012899838e-10, 
    1.7019770779284328e-10, 1.6894442240301829e-10, 1.6759369386730853e-10, 
    1.6615127506725308e-10, 1.6462683800599662e-10, 1.6303386034991292e-10, 
    1.6138928293064709e-10, 1.5971303345276033e-10, 1.5802734655585173e-10, 
    1.5635600077393338e-10, 1.5472342019670135e-10, 1.5315375756348112e-10, 
    1.5166992331890671e-10, 1.502926589292005e-10, 1.490396356035592e-10, 
    1.4792466770545763e-10, 1.4695704023269606e-10, 1.4614102441708612e-10, 
    1.4547559290426566e-10, 1.4495442017283507e-10, 1.4456612697755101e-10, 
    1.4429487115226389e-10, 1.4412118149491836e-10, 1.4402308582630385e-10, 
    1.4397738983226357e-10, 1.4396107942941649e-10, 1.4395267754403143e-10, 
    1.4393349190785447e-10, 1.4388857978140058e-10, 1.4380740527465515e-10, 
    1.4368404176172962e-10, 1.4351698644306983e-10, 1.4330855033520121e-10, 
    1.4306393720028357e-10, 1.4279007942866682e-10, 1.4249441038709275e-10, 
    1.4218366115825693e-10, 1.4186285625142179e-10, 1.4153457796019981e-10, 
    1.411986030797781e-10, 1.4085187094634683e-10, 1.4048884666407297e-10, 
    1.4010213399525373e-10, 1.3968331003881337e-10, 1.3922381466657187e-10, 
    1.3871584174657097e-10, 1.3815307694301521e-10, 1.3753126017855473e-10, 
    1.3684846406977123e-10, 1.3610515062101754e-10, 1.3530396364701406e-10, 
    1.3444935912597458e-10, 1.3354709105944658e-10, 1.3260368066113705e-10, 
    1.3162589909116774e-10, 1.3062037535037145e-10, 1.2959330436576113e-10, 
    1.2855038023118866e-10, 1.2749681809654251e-10, 1.2643759121566128e-10, 
    1.2537770560699503e-10, 1.2432256520298611e-10, 1.2327828212446919e-10, 
    1.2225195563276196e-10, 1.2125180140394475e-10, 1.2028717462949648e-10, 
    1.1936838569172019e-10, 1.1850641112731536e-10, 1.1771241837108642e-10, 
    1.1699724209169068e-10, 1.163707462874846e-10, 1.1584123782394707e-10, 
    1.1541486677248615e-10, 1.1509515957905239e-10, 1.1488262816070236e-10, 
    1.147745633272404e-10, 1.1476495519890018e-10, 1.1484460823742749e-10, 
    1.1500137337851828e-10, 1.1522054202446361e-10, 1.1548534513962061e-10, 
    1.1577755136576848e-10, 1.1607808603599259e-10, 1.1636773794721377e-10, 
    1.1662780228347756e-10, 1.1684076403234119e-10, 1.1699088254666191e-10, 
    1.1706476045817903e-10, 1.1705177867716813e-10, 1.1694448331406217e-10, 
    1.1673880280384714e-10, 1.1643418139561762e-10, 1.1603351746226627e-10, 
    1.1554300200199398e-10, 1.1497173650566216e-10, 1.1433125254473078e-10, 
    1.1363485207673675e-10, 1.1289688158671668e-10, 1.1213188467932568e-10, 
    1.1135379120021456e-10, 1.1057510446211359e-10, 1.0980623225444327e-10, 
    1.0905493855286887e-10, 1.0832605212604587e-10, 1.07621381586804e-10, 
    1.0693992545726389e-10, 1.0627830644743123e-10, 1.0563144327596455e-10, 
    1.0499335219604876e-10, 1.0435806418858823e-10, 1.0372049423043941e-10, 
    1.0307726837169822e-10, 1.0242730492110533e-10, 1.0177222463234218e-10, 
    1.01116414764494e-10, 1.004668342059483e-10, 9.9832528189622849e-11, 
    9.9223919978922606e-11, 9.8651926818791622e-11, 9.8127038205426386e-11, 
    9.7658382039507876e-11, 9.7252951074746125e-11, 9.6914971605570485e-11, 
    9.6645559345435315e-11, 9.6442608258786671e-11, 9.6300975070158377e-11, 
    9.6212871465803723e-11, 9.6168468995903379e-11, 9.6156598761164344e-11, 
    9.6165526693018113e-11, 9.6183679157385285e-11, 9.6200339255257361e-11, 
    9.6206167150447623e-11, 9.6193629616917686e-11, 9.6157231997834195e-11, 
    9.6093638305297935e-11, 9.6001619383587434e-11, 9.5881935046060061e-11, 
    9.5737090210762593e-11, 9.5571078933109195e-11, 9.5389057639415704e-11, 
    9.5197034588222504e-11, 9.5001526398320498e-11, 9.4809264828528783e-11, 
    9.4626866304517845e-11, 9.446057342450152e-11, 9.4315967199355641e-11, 
    9.4197748005710507e-11, 9.4109494875749405e-11, 9.4053492317038542e-11, 
    9.4030548639421836e-11, 9.403987552204885e-11, 9.4078966735106361e-11, 
    9.4143549235386662e-11, 9.4227546686531977e-11, 9.4323131348907996e-11, 
    9.4420808047480138e-11, 9.4509611535913769e-11, 9.457735520121139e-11, 
    9.4611004865277936e-11, 9.4597112558202869e-11, 9.4522364373388406e-11, 
    9.4374153168334091e-11, 9.4141215011241069e-11, 9.3814238882963102e-11, 
    9.338646426255929e-11, 9.2854154661992891e-11, 9.2217006980329933e-11, 
    9.1478355476888277e-11, 9.0645261327627373e-11, 8.9728384491023492e-11, 
    8.8741716624068394e-11, 8.7702110224163834e-11, 8.6628703821952001e-11, 
    8.5542197589742144e-11, 8.4464063786225179e-11, 8.3415687964441263e-11, 
    8.2417507438576046e-11, 8.148816277638802e-11, 8.0643730004789066e-11, 
    7.9897030951268608e-11, 7.9257134823915413e-11, 7.8728984190613449e-11, 
    7.8313280275151193e-11, 7.8006557376100988e-11, 7.7801500375545664e-11, 
    7.7687449259502274e-11, 7.7651096932252904e-11, 7.7677283982084153e-11, 
    7.77498790556081e-11, 7.7852633554519364e-11, 7.7969981749013413e-11, 
    7.8087706556804835e-11, 7.8193467891962433e-11, 7.8277089617921437e-11, 
    7.8330721846603096e-11, 7.8348781449522302e-11, 7.8327782723203791e-11, 
    7.826604855727221e-11, 7.8163380599139872e-11, 7.8020702195079572e-11, 
    7.7839733801251066e-11, 7.7622701587068318e-11, 7.737211053227589e-11, 
    7.7090562816265412e-11, 7.6780636511287301e-11, 7.6444790057912229e-11, 
    7.6085301326753145e-11, 7.5704218134884671e-11, 7.5303320792052622e-11, 
    7.4884098821637757e-11, 7.4447749640018745e-11, 7.3995190344783463e-11, 
    7.3527114253601755e-11, 7.3044086045867534e-11, 7.2546663409055951e-11, 
    7.2035554307357526e-11, 7.1511793735483572e-11, 7.0976895537969559e-11, 
    7.0433000226066777e-11, 6.9882963395248616e-11, 6.9330390606381176e-11, 
    6.8779583649221097e-11, 6.8235430892403455e-11, 6.7703218343814668e-11, 
    6.7188396497226881e-11, 6.6696301556545318e-11, 6.6231872004357428e-11, 
    6.5799368637889072e-11, 6.5402120793010774e-11, 6.5042303590315668e-11, 
    6.4720777793429071e-11, 6.4436968432405867e-11, 6.4188818058808977e-11, 
    6.3972797908484394e-11, 6.3783992283433116e-11, 6.3616262324386939e-11, 
    6.3462491095710551e-11, 6.3314908046543542e-11, 6.316549561635889e-11, 
    6.3006468229623568e-11, 6.2830779361467906e-11, 6.2632640678763169e-11, 
    6.2408018421381999e-11, 6.2155009221417874e-11, 6.1874113244813232e-11, 
    6.1568317414090884e-11, 6.1242973330593437e-11, 6.0905468108297052e-11, 
    6.056470279598998e-11, 6.0230398988312506e-11, 5.9912312698840535e-11, 
    5.9619420461338413e-11, 5.9359142635539975e-11, 5.9136694630499791e-11, 
    5.8954612907166044e-11, 5.8812520620057491e-11, 5.8707129200871687e-11, 
    5.8632491215977548e-11, 5.8580463993215144e-11, 5.854134758273492e-11, 
    5.8504624711411489e-11, 5.8459747602360638e-11, 5.8396898757921083e-11, 
    5.8307668278105542e-11, 5.8185598450057333e-11, 5.8026571167125849e-11, 
    5.782901808247954e-11, 5.7593939921907944e-11, 5.7324756772391472e-11, 
    5.7027017587542033e-11, 5.6707976416163651e-11, 5.6376075572436713e-11, 
    5.6040381983008394e-11, 5.5710005952627164e-11, 5.5393532192194148e-11, 
    5.5098511699255453e-11, 5.4831037604524372e-11, 5.4595418128373922e-11, 
    5.4393988109251379e-11, 5.4227044743805327e-11, 5.4092909420288921e-11, 
    5.3988109896806938e-11, 5.3907636504332236e-11, 5.3845274069658998e-11, 
    5.3793939775740436e-11, 5.3746009763486263e-11, 5.3693615047829835e-11, 
    5.3628864544044066e-11, 5.3544009947672805e-11, 5.3431546680053581e-11, 
    5.3284274671826407e-11, 5.3095354144314514e-11, 5.2858376991080065e-11, 
    5.2567499841786357e-11, 5.2217647320443378e-11, 5.1804813503265484e-11, 
    5.1326440982436267e-11, 5.0781845719891775e-11, 5.0172673932127632e-11, 
    4.9503296636964188e-11, 4.8781114983426289e-11, 4.801669351175412e-11, 
    4.7223693873980022e-11, 4.641855168728648e-11, 4.5619928359483599e-11, 
    4.4847914104944046e-11, 4.4123080175546078e-11, 4.3465392795204274e-11, 
    4.2893121219047829e-11, 4.2421800279036344e-11, 4.2063349346902387e-11, 
    4.1825397670769268e-11, 4.1710903192092995e-11, 4.1718050078930289e-11, 
    4.1840455458223181e-11, 4.2067631342556694e-11, 4.238566786315011e-11, 
    4.2778053182137617e-11, 4.3226579306732593e-11, 4.3712228561331036e-11, 
    4.4216004490098584e-11, 4.4719635148141977e-11, 4.520613838992912e-11, 
    4.5660209451303214e-11, 4.6068469452116518e-11, 4.6419555162701187e-11, 
    4.6704138011331724e-11, 4.6914835579336856e-11, 4.7046134637632789e-11, 
    4.7094281763670886e-11, 4.7057230303158806e-11, 4.6934597477048376e-11, 
    4.6727686635595726e-11, 4.6439523218215441e-11, 4.6074920041048908e-11, 
    4.5640508542741976e-11, 4.5144763734198146e-11, 4.4597931329252045e-11, 
    4.4011893900308289e-11, 4.3399922732059573e-11, 4.2776343369047964e-11, 
    4.2156071373738683e-11, 4.1554112614475639e-11, 4.0984970705515886e-11, 
    4.0462079274961001e-11, 3.9997234115297084e-11, 3.9600118472027794e-11, 
    3.9277921588039273e-11, 3.9035112754232037e-11, 3.8873357507837995e-11, 
    3.8791630068437757e-11, 3.8786431582093941e-11, 3.8852204452798486e-11, 
    3.8981782743298603e-11, 3.9166952263470083e-11, 3.939898624370192e-11, 
    3.966918192764594e-11, 3.9969286052575929e-11, 4.0291867985780432e-11, 
    4.0630515059821682e-11, 4.0979959398346834e-11, 4.1336011256610646e-11, 
    4.1695438052860653e-11, 4.2055704672740799e-11, 4.2414694490889528e-11, 
    4.277035978396098e-11, 4.3120428390107557e-11, 4.3462110126157795e-11, 
    4.3791919417911757e-11, 4.4105561104715883e-11, 4.4397967815185175e-11, 
    4.466340809937956e-11, 4.4895754992520284e-11, 4.5088788239381159e-11, 
    4.5236591549434023e-11, 4.5333947034141716e-11, 4.5376723125356486e-11, 
    4.5362171961374632e-11, 4.528918000103778e-11, 4.5158333739926961e-11, 
    4.4971926466487525e-11, 4.4733782822616316e-11, 4.4449034760017525e-11, 
    4.4123763512070966e-11, 4.3764660502186353e-11, 4.3378649079210963e-11, 
    4.2972583451309806e-11, 4.2552981040141563e-11, 4.2125899676910406e-11, 
    4.1696847426124049e-11, 4.1270845298492137e-11, 4.0852509499470104e-11, 
    4.0446211265589267e-11, 4.0056201685018974e-11, 3.968674709931344e-11, 
    3.9342156050099829e-11, 3.9026765043969419e-11, 3.8744793649770742e-11, 
    3.850014931569598e-11, 3.8296116242502685e-11, 3.8135049215388263e-11, 
    3.8018027482929335e-11, 3.7944577191978286e-11, 3.7912447855545772e-11, 
    3.7917541057624173e-11, 3.7953929985725095e-11, 3.8014077385105807e-11, 
    3.8089165387047848e-11, 3.8169573136557342e-11, 3.8245423662421981e-11, 
    3.8307198793248216e-11, 3.8346319651351744e-11, 3.835570778252289e-11, 
    3.8330190895100333e-11, 3.8266815922899475e-11, 3.8164950711049096e-11, 
    3.8026254074506716e-11, 3.7854427822758958e-11, 3.765487866820475e-11, 
    3.7434228831991681e-11, 3.719980217343852e-11, 3.6959055454765094e-11, 
    3.6719086195268888e-11, 3.6486171461319042e-11, 3.6265450155947086e-11, 
    3.6060691641789043e-11, 3.5874233636688804e-11, 3.5707008871450612e-11, 
    3.5558713176956078e-11, 3.542804020424913e-11, 3.5313009304098403e-11, 
    3.5211277030366331e-11, 3.5120503830769294e-11, 3.5038658641764456e-11, 
    3.4964309722316788e-11, 3.4896805745009913e-11, 3.483641986001892e-11, 
    3.4784359091252275e-11, 3.4742714049492404e-11, 3.4714274601469145e-11, 
    3.4702289515124804e-11, 3.471013046635089e-11, 3.4740931599979452e-11, 
    3.4797183818627204e-11, 3.4880372825662789e-11, 3.4990641509610901e-11, 
    3.5126570064492109e-11, 3.5285031327745188e-11, 3.546122754218174e-11, 
    3.5648822078426564e-11, 3.5840247215674668e-11, 3.6027097649827184e-11, 
    3.6200635966511458e-11, 3.6352311006783442e-11, 3.6474297044385281e-11, 
    3.6559965637021716e-11, 3.6604294141668973e-11, 3.6604106058157492e-11, 
    3.6558212295279448e-11, 3.6467381488973729e-11, 3.6334194736866025e-11, 
    3.6162730067684894e-11, 3.5958210253908225e-11, 3.5726552804079819e-11, 
    3.5473930952639098e-11, 3.5206312710023059e-11, 3.4929088337990192e-11, 
    3.4646744492289677e-11, 3.4362663550586781e-11, 3.4079024828356494e-11, 
    3.3796841993632255e-11, 3.3516116778004581e-11, 3.323612672454492e-11, 
    3.2955791516355389e-11, 3.2674135786839212e-11, 3.2390762708629486e-11, 
    3.2106344441853131e-11, 3.1823017613577333e-11, 3.1544705120846218e-11, 
    3.1277248674110726e-11, 3.1028377431398957e-11, 3.0807434603032147e-11, 
    3.0624923634720899e-11, 3.0491838653312506e-11, 3.0418872695209237e-11, 
    3.0415531103000564e-11, 3.0489263117105714e-11, 3.0644650408032512e-11, 
    3.0882784471337677e-11, 3.1200864264616623e-11, 3.1592087399920533e-11, 
    3.2045832963202108e-11, 3.2548161484449543e-11, 3.3082579990856223e-11, 
    3.3631019785703616e-11, 3.4174940640406344e-11, 3.4696495299824654e-11, 
    3.5179610967802579e-11, 3.5610952242087958e-11, 3.5980636557312783e-11, 
    3.6282689677461882e-11, 3.6515153684480829e-11, 3.6679900376128708e-11, 
    3.678211923333416e-11, 3.6829569973970908e-11, 3.6831630846244509e-11, 
    3.6798268009440076e-11, 3.6738999385815382e-11, 3.6661951447097927e-11, 
    3.6573091376856414e-11, 3.6475718474036183e-11, 3.6370241747237797e-11, 
    3.6254264807042116e-11, 3.6122972552558714e-11, 3.5969773619882124e-11, 
    3.5787091686139243e-11, 3.5567287545323799e-11, 3.530356233254256e-11, 
    3.4990776406091283e-11, 3.4626085698915637e-11, 3.4209364796375229e-11, 
    3.3743353882324028e-11, 3.3233561414526421e-11, 3.2687910520457222e-11, 
    3.2116223158269635e-11, 3.152956587805825e-11, 3.0939574256462307e-11, 
    3.035778206571732e-11, 2.9795049651380739e-11, 2.9261135031363749e-11, 
    2.8764417054894575e-11, 2.8311763628975895e-11, 2.7908569500432265e-11, 
    2.7558886529577407e-11, 2.7265639296694392e-11, 2.7030853662780092e-11, 
    2.6855893162221733e-11, 2.6741617741352151e-11, 2.6688495218848339e-11, 
    2.6696626145456764e-11, 2.6765690582653566e-11, 2.6894802717457615e-11, 
    2.7082353905573365e-11, 2.7325810091162466e-11, 2.7621542959384931e-11, 
    2.7964672069649462e-11, 2.8349004223825756e-11, 2.8767041816725236e-11, 
    2.9210108288953516e-11, 2.9668549015988266e-11, 3.0132051458780519e-11, 
    3.0590018963706009e-11, 3.1032010502021793e-11, 3.1448164096539466e-11, 
    3.1829630116307037e-11, 3.2168912260562742e-11, 3.246013962484826e-11, 
    3.2699214948328825e-11, 3.2883847233474951e-11, 3.3013442352434272e-11, 
    3.3088907568626094e-11, 3.3112347035870487e-11, 3.3086717533915201e-11, 
    3.3015460884504561e-11, 3.2902161439582594e-11, 3.2750250614022636e-11, 
    3.2562808624131619e-11, 3.2342441514452479e-11, 3.2091281575411655e-11, 
    3.1811073666311603e-11, 3.1503359270685499e-11, 3.1169677613304058e-11, 
    3.0811823598361013e-11, 3.043207044470365e-11, 3.003336032855862e-11, 
    2.9619404002718311e-11, 2.9194708297792557e-11, 2.8764485794736075e-11, 
    2.8334482686588546e-11, 2.7910704416302298e-11, 2.7499089284781408e-11, 
    2.7105137810620044e-11, 2.6733549574283525e-11, 2.6387863163918688e-11, 
    2.6070175734874983e-11, 2.5780926573830114e-11, 2.5518793456689509e-11, 
    2.528068697499133e-11, 2.5061878493356735e-11, 2.4856224286385024e-11, 
    2.465651153394456e-11, 2.445487776182002e-11, 2.4243314455929041e-11, 
    2.4014178909439144e-11, 2.3760739236642396e-11, 2.3477673304939545e-11, 
    2.3161517253720102e-11, 2.2811001093310254e-11, 2.2427282850076983e-11, 
    2.2014028397121256e-11, 2.157734269184079e-11, 2.1125548801211844e-11, 
    2.0668834464039445e-11, 2.0218742725985013e-11, 1.9787592436088704e-11, 
    1.9387825808862803e-11, 1.903132017217137e-11, 1.8728708164435396e-11, 
    1.848876489972801e-11, 1.8317854512306086e-11, 1.8219525121043892e-11, 
    1.8194232176110224e-11, 1.8239256773298045e-11, 1.8348772864192023e-11, 
    1.8514136634855122e-11, 1.87243187027654e-11, 1.8966509809286493e-11, 
    1.9226825091042752e-11, 1.9491109029850068e-11, 1.9745728894069021e-11, 
    1.9978373757528434e-11, 2.0178753576076178e-11, 2.0339183331843437e-11, 
    2.0455000389477871e-11, 2.0524810192741518e-11, 2.0550509192627982e-11, 
    2.0537145369569419e-11, 2.049257601821987e-11, 2.0426986867057971e-11, 
    2.0352271279167717e-11, 2.0281335988246279e-11, 2.0227344253136285e-11, 
    2.0202966426159715e-11, 2.021962500140366e-11, 2.0286834527902353e-11, 
    2.041160424681837e-11, 2.0597990342743616e-11, 2.0846765696743996e-11, 
    2.1155271518702362e-11, 2.1517444731601377e-11, 2.1924025428893151e-11, 
    2.2362921355613353e-11, 2.2819758668488026e-11, 2.3278537682239765e-11, 
    2.3722402589581651e-11, 2.4134449856770389e-11, 2.4498551471104226e-11, 
    2.4800126444587759e-11, 2.5026830699228201e-11, 2.5169102665897823e-11, 
    2.5220558568277126e-11, 2.5178203461093567e-11, 2.5042456892420478e-11, 
    2.4816991724659979e-11, 2.4508434765887943e-11, 2.4125902090423505e-11, 
    2.3680481481542485e-11, 2.3184637935246111e-11, 2.2651629991019573e-11, 
    2.2094931062176887e-11, 2.1527739614236534e-11, 2.096254307435044e-11, 
    2.0410797614215783e-11, 1.9882694253959051e-11, 1.9387018430802353e-11, 
    1.893107898733881e-11, 1.8520716513245971e-11, 1.8160320801422127e-11, 
    1.7852909032190481e-11, 1.7600184898025894e-11, 1.7402623665614443e-11, 
    1.7259535631086198e-11, 1.7169144891231176e-11, 1.7128660358535823e-11, 
    1.7134361199160037e-11, 1.7181701570494428e-11, 1.7265435505842387e-11, 
    1.7379760549245374e-11, 1.7518501440669174e-11, 1.7675309968045225e-11, 
    1.7843904739927645e-11, 1.8018297239398437e-11, 1.8193053837128114e-11, 
    1.8363540585121464e-11, 1.8526148482545089e-11, 1.8678491261367924e-11, 
    1.881954842437934e-11, 1.8949753454671261e-11, 1.9070994620638706e-11, 
    1.9186531248968325e-11, 1.9300827271575053e-11, 1.941928162438368e-11, 
    1.9547908303989599e-11, 1.9692933094072801e-11, 1.9860388331028379e-11, 
    2.0055692471577991e-11, 2.0283293499368442e-11, 2.0546337743390885e-11, 
    2.084646322358504e-11, 2.1183673741590611e-11, 2.1556306056896547e-11, 
    2.1961109741666921e-11, 2.2393378417737794e-11, 2.2847126520561112e-11, 
    2.331530970866946e-11, 2.3790030799770494e-11, 2.4262755995320222e-11, 
    2.4724509367596161e-11, 2.5166075148430131e-11, 2.5578202663406137e-11, 
    2.5951839049566724e-11, 2.6278398723629133e-11, 2.6550074025863655e-11, 
    2.6760184735997772e-11, 2.6903552237763193e-11, 2.6976864521165584e-11, 
    2.6979007463430289e-11, 2.6911306545718087e-11, 2.6777666010802856e-11, 
    2.6584541422154851e-11, 2.6340747770768088e-11, 2.6057112201685263e-11, 
    2.5745947652970095e-11, 2.5420401252078403e-11, 2.5093728149225377e-11, 
    2.4778531695229051e-11, 2.4486036324897061e-11, 2.422544536106479e-11, 
    2.40034568792713e-11, 2.3823930205304233e-11, 2.3687782019013293e-11, 
    2.3593074165418917e-11, 2.3535296234136984e-11, 2.3507811114089782e-11, 
    2.3502421934705883e-11, 2.3509992240943954e-11, 2.3521088548427122e-11, 
    2.3526582211017845e-11, 2.3518172130445111e-11, 2.3488773515216583e-11, 
    2.3432800513927364e-11, 2.3346292744771459e-11, 2.3226933249339301e-11, 
    2.3073947982127867e-11, 2.2887931187163071e-11, 2.2670629555709757e-11, 
    2.2424700555644877e-11, 2.2153465370952567e-11, 2.1860694686910774e-11, 
    2.155040564180314e-11, 2.1226694792322325e-11, 2.0893592544040532e-11, 
    2.0554936073452274e-11, 2.0214262504661811e-11, 1.9874719093279525e-11, 
    1.9538995758919438e-11, 1.9209291647929461e-11, 1.8887317907847225e-11, 
    1.8574360568633974e-11, 1.8271389622365606e-11, 1.7979219390774753e-11, 
    1.7698705313946013e-11, 1.7430945338463538e-11, 1.7177450655195424e-11, 
    1.6940264049818848e-11, 1.6721964404927704e-11, 1.6525557351002801e-11, 
    1.6354231060225331e-11, 1.6210973444423868e-11, 1.609811526415223e-11, 
    1.6016810492434406e-11, 1.5966523660221124e-11, 1.5944616252161691e-11, 
    1.5946065843780506e-11, 1.5963396311971683e-11, 1.5986825597816742e-11, 
    1.6004675232853223e-11, 1.6003988196603759e-11, 1.5971332573641022e-11, 
    1.5893732407230388e-11, 1.5759623150723928e-11, 1.5559767371428953e-11, 
    1.5288054598065151e-11, 1.4942085343210611e-11, 1.4523526577789119e-11, 
    1.4038180062636309e-11, 1.3495758344107971e-11, 1.2909401412319964e-11, 
    1.2294949114202879e-11, 1.1670029716242445e-11, 1.1053043058587156e-11, 
    1.0462094909937264e-11, 9.9139799177069203e-12, 9.4232588724018868e-12, 
    9.0015221074324143e-12, 8.6568785999647739e-12, 8.3936924679970673e-12, 
    8.2125913585602303e-12, 8.1107329692420917e-12, 8.0822913928968634e-12, 
    8.1191152610649009e-12, 8.2115104578019428e-12, 8.3490501490454319e-12, 
    8.5213644530941249e-12, 8.7188447231457546e-12, 8.9332008302226395e-12, 
    9.1578634240440788e-12, 9.3881845300047035e-12, 9.6214668980578123e-12, 
    9.8568265556100897e-12, 1.0094925702199275e-11, 1.0337588307873246e-11, 
    1.0587364139825938e-11, 1.084706411097673e-11, 1.1119290638254734e-11, 
    1.1405983528691678e-11, 1.170803656769049e-11, 1.2024964321887296e-11, 
    1.2354672937941578e-11, 1.2693315155835335e-11, 1.3035283092439324e-11, 
    1.3373322024752615e-11, 1.3698794273050064e-11, 1.40020641836294e-11, 
    1.4273020226165451e-11, 1.450168762374774e-11, 1.4678898584113947e-11, 
    1.4796976664541449e-11, 1.4850361127594552e-11, 1.4836137776258986e-11, 
    1.4754407158188581e-11, 1.4608442694389018e-11, 1.4404643367829909e-11, 
    1.4152235848930377e-11, 1.3862788935725571e-11, 1.3549530663710603e-11, 
    1.3226560767328202e-11, 1.290800084326595e-11, 1.2607164720882873e-11, 
    1.2335788253674706e-11, 1.2103424759499e-11, 1.1916983561005255e-11, 
    1.1780500296998746e-11, 1.1695104979016937e-11, 1.1659198293150291e-11, 
    1.1668794454267894e-11, 1.1718018958240581e-11, 1.1799673612892697e-11, 
    1.1905870828246864e-11, 1.2028633521625727e-11, 1.2160463381402709e-11, 
    1.2294785567525868e-11, 1.2426288784119209e-11, 1.2551112215096572e-11, 
    1.2666880063757633e-11, 1.2772592709300488e-11, 1.2868400570294024e-11, 
    1.2955275382090793e-11, 1.3034636510754046e-11, 1.310795923430771e-11, 
    1.3176427569615237e-11, 1.3240639171029603e-11, 1.3300428340949565e-11, 
    1.335480922769174e-11, 1.3402059793051129e-11, 1.3439898462169318e-11, 
    1.3465807215388341e-11, 1.3477387184191484e-11, 1.3472768040046663e-11, 
    1.3450976016061329e-11, 1.3412248805003623e-11, 1.3358217826228238e-11, 
    1.3291952518041507e-11, 1.3217818297253174e-11, 1.3141177625752308e-11, 
    1.3067901203169307e-11, 1.3003784611480974e-11, 1.2953880241963566e-11, 
    1.2921830543246822e-11, 1.2909285550988235e-11, 1.291546484893589e-11, 
    1.293692030410005e-11, 1.2967576086571857e-11, 1.2999022909512325e-11, 
    1.3021095499163584e-11, 1.3022649313558846e-11, 1.2992520334882939e-11, 
    1.2920531542071361e-11, 1.279847949559752e-11, 1.2621007319288177e-11, 
    1.2386265580679555e-11, 1.2096287079456583e-11, 1.1757076787566483e-11, 
    1.1378372820986607e-11, 1.0973128719590555e-11, 1.0556745481639034e-11, 
    1.0146141576804284e-11, 9.7587314506162722e-12, 9.4113942263089479e-12, 
    9.1195204190784339e-12, 8.8962004324503021e-12, 8.7515796199418426e-12, 
    8.6924589562331522e-12, 8.7221006653263555e-12, 8.8402650948005542e-12, 
    9.043453595140172e-12, 9.3253211208146854e-12, 9.677201207787806e-12, 
    1.0088737405898277e-11, 1.0548542017909042e-11, 1.1044859357218137e-11, 
    1.156616955347888e-11, 1.2101722598982382e-11, 1.2641956539922324e-11, 
    1.3178790630900164e-11, 1.3705782738085877e-11, 1.4218155599929377e-11, 
    1.4712693140868839e-11, 1.518755995078618e-11, 1.5642019668686625e-11, 
    1.6076134038037964e-11, 1.6490450927164173e-11, 1.6885702295381314e-11, 
    1.7262544648137452e-11, 1.7621361972885104e-11, 1.796212582023777e-11, 
    1.8284332838173268e-11, 1.8586998787177017e-11, 1.8868725841379568e-11, 
    1.9127798690364663e-11, 1.9362332287979134e-11, 1.9570445298922547e-11, 
    1.9750437000899601e-11, 1.9900953244619306e-11, 2.002114732743251e-11, 
    2.0110789923432359e-11, 2.0170341755446986e-11, 2.0200972951896767e-11, 
    2.0204526771053901e-11, 2.018342545949128e-11, 2.014054070653229e-11, 
    2.0079040780354146e-11, 2.0002219311685267e-11, 1.9913332784640817e-11, 
    1.9815461210805861e-11, 1.9711394997204107e-11, 1.9603548559140902e-11, 
    1.9493906249561164e-11, 1.9383983908317286e-11, 1.9274803435568245e-11, 
    1.9166876613011554e-11, 1.9060182574009603e-11, 1.8954159661013663e-11, 
    1.8847702017647543e-11, 1.8739187059583232e-11, 1.86265274189909e-11, 
    1.850727423630717e-11, 1.8378752644267752e-11, 1.8238249246834456e-11, 
    1.8083204371755093e-11, 1.7911427790143474e-11, 1.7721281380468806e-11, 
    1.7511835155237598e-11, 1.7282946474625784e-11, 1.7035284076634337e-11, 
    1.6770284093345151e-11, 1.6490040853490543e-11, 1.619715541617443e-11, 
    1.5894572291766205e-11, 1.5585404235221982e-11, 1.5272800555230123e-11, 
    1.4959836716087369e-11, 1.4649466291308378e-11, 1.4344507534543512e-11, 
    1.4047673311145353e-11, 1.3761628682420859e-11, 1.3489047932754029e-11, 
    1.3232664512862726e-11, 1.2995284774528437e-11, 1.2779778017562122e-11, 
    1.2589003379922175e-11, 1.2425693959591865e-11, 1.2292296936229186e-11, 
    1.2190792861270823e-11, 1.2122509170340935e-11, 1.2087917182908764e-11, 
    1.2086492509858295e-11, 1.2116618631633109e-11, 1.2175555987199471e-11, 
    1.2259493962616235e-11, 1.2363680843836517e-11, 1.2482624789434065e-11, 
    1.2610349974662198e-11, 1.2740674182806661e-11, 1.2867494267410864e-11, 
    1.298505320614108e-11, 1.308815699377936e-11, 1.3172322678206393e-11, 
    1.323387570485662e-11, 1.3269989584977235e-11, 1.3278675057957753e-11, 
    1.32587548972815e-11, 1.3209825341577425e-11, 1.3132256635562787e-11, 
    1.3027205738336345e-11, 1.2896651021451494e-11, 1.2743462176546949e-11, 
    1.2571441365423485e-11, 1.2385342705091334e-11, 1.2190818527541445e-11, 
    1.1994275967191639e-11, 1.1802623937419473e-11, 1.162290254468656e-11, 
    1.1461837352686766e-11, 1.1325319784818559e-11, 1.121788768266554e-11, 
    1.1142246302688632e-11, 1.1098912066720176e-11, 1.1086002720033576e-11, 
    1.1099238043459688e-11, 1.1132160722698647e-11, 1.117656312514542e-11, 
    1.1223092019072378e-11, 1.1262006632389226e-11, 1.1283965776578719e-11, 
    1.1280823274927512e-11, 1.1246324529852184e-11, 1.1176640663873284e-11, 
    1.1070711210556953e-11, 1.0930353141471766e-11, 1.0760138381374362e-11, 
    1.0567067367027308e-11, 1.0360072411049244e-11, 1.0149410130447949e-11, 
    9.9459947121567843e-12, 9.760740648103908e-12, 9.6039388713459306e-12, 
    9.4847431522865393e-12, 9.4107502075794509e-12, 9.387705226584531e-12, 
    9.4193289135437466e-12, 9.507252564369247e-12, 9.6510469297857984e-12, 
    9.8483381296093571e-12, 1.009498447850252e-11, 1.0385314613975201e-11, 
    1.0712407169745295e-11, 1.1068404318071326e-11, 1.144484848060777e-11, 
    1.1833043830068242e-11, 1.2224391898845677e-11, 1.2610724597284315e-11, 
    1.2984586685596814e-11, 1.3339467059532192e-11, 1.3669953196298606e-11, 
    1.3971816933134002e-11, 1.4242013096193046e-11, 1.4478609441150739e-11, 
    1.4680646352698949e-11, 1.4847960715369518e-11, 1.4980976475265472e-11, 
    1.5080481900570601e-11, 1.5147415749243253e-11, 1.518268322384226e-11, 
    1.5186993872272839e-11, 1.516075148035668e-11, 1.5103976977614489e-11, 
    1.5016296015242171e-11, 1.4896960202731058e-11, 1.4744927036571829e-11, 
    1.4558979909131817e-11, 1.4337882746040619e-11, 1.4080565654926925e-11, 
    1.378633369552004e-11, 1.3455072783981005e-11, 1.3087453282446409e-11, 
    1.2685105314279834e-11, 1.2250750061572929e-11, 1.1788278037869148e-11, 
    1.1302756081736526e-11, 1.0800362969853639e-11, 1.028824019237512e-11, 
    9.7742700645194174e-12, 9.2667815370644017e-12, 8.7742096208815827e-12, 
    8.3047175545396197e-12, 7.865808993080825e-12, 7.4639758220331159e-12, 
    7.1043689795826777e-12, 6.7905671970410354e-12, 6.5244233428175129e-12, 
    6.3060292228398355e-12, 6.1337732671822751e-12, 6.004523821664387e-12, 
    5.9138841984094434e-12, 5.8565094509949207e-12, 5.8264667198360423e-12, 
    5.8175928333333669e-12, 5.8238228309140479e-12, 5.8394845885720506e-12, 
    5.8595178282188603e-12, 5.8796442047705337e-12, 5.8964701792630594e-12, 
    5.9075494111877925e-12, 5.9114064535140851e-12,
  // Sqw-total(6, 0-1999)
    0.027516003292299508, 0.027513148260365917, 0.027504524394755259, 
    0.02748995904305554, 0.02746917624026737, 0.027441813052599198, 
    0.02740743999727811, 0.027365583543813802, 0.027315748700648616, 
    0.02725743996478612, 0.027190179392486091, 0.027113521135029801, 
    0.027027062361702769, 0.026930450960735392, 0.026823390697603818, 
    0.026705644592524183, 0.026577037175570008, 0.026437456048023417, 
    0.0262868529045466, 0.026125243936872163, 0.025952709411915527, 
    0.025769392227756434, 0.025575495391497661, 0.025371278587879097, 
    0.025157054245847014, 0.024933183684241411, 0.024700073962374433, 
    0.024458175941037059, 0.024207983778101346, 0.023950035684054623, 
    0.023684915321797558, 0.023413252843576055, 0.023135724305324248, 
    0.02285304815373496, 0.022565977678178008, 0.022275288750346955, 
    0.021981762789935199, 0.021686165611606332, 0.021389223523195701, 
    0.021091598648964625, 0.020793865847932747, 0.02049649371469927, 
    0.020199831953594101, 0.019904106912616182, 0.019609426298813487, 
    0.019315793155067845, 0.019023128169673352, 0.018731298438079538, 
    0.018440150022277519, 0.01814954116148754, 0.017859372849901387, 
    0.017569613741889079, 0.017280316951698169, 0.016991627214016983, 
    0.016703777953475982, 0.016417078937920576, 0.016131896216741479, 
    0.01584862683937896, 0.015567671310794784, 0.01528940681867855, 
    0.015014163965551046, 0.014742209116351721, 0.014473733631479168, 
    0.014208850326511816, 0.013947596618409518, 0.013689943103148779, 
    0.013435805846445926, 0.013185060496824904, 0.012937556439651101, 
    0.012693129549921587, 0.012451612588468136, 0.012212842825286027, 
    0.011976666973564372, 0.011742943906282133, 0.01151154586035545, 
    0.01128235889989641, 0.011055283328133325, 0.010830234546520904, 
    0.010607144610241957, 0.010385964472793704, 0.010166666691355545, 
    0.0099492482079255162, 0.0097337327419476198, 0.0095201723275600645, 
    0.0093086475918645606, 0.0090992664836307222, 0.0088921613072508333, 
    0.0086874840786493636, 0.0084854003846157548, 0.008286082082760219, 
    0.0080896993145028878, 0.0078964124060853565, 0.007706364289750303, 
    0.0075196740768608611, 0.0073364323479540106, 0.0071566985890802199, 
    0.0069805010060082504, 0.0068078387053471523, 0.0066386859716806041, 
    0.0064729981266575991, 0.0063107182656501415, 0.0061517840616126555, 
    0.0059961338250171135, 0.0058437111186726287, 0.0056944674347916601, 
    0.0055483627203019867, 0.0054053638443434769, 0.005265441392813504, 
    0.0051285654047599381, 0.0049947008002877366, 0.004863803271006756, 
    0.0047358163119685104, 0.0046106698865354071, 0.0044882809649730076, 
    0.0043685559042163126, 0.0042513943817439823, 0.0041366943965090008, 
    0.0040243577290282571, 0.003914295221596328, 0.0038064312944399827, 
    0.0037007072386067851, 0.003597082997397404, 0.0034955373376098766, 
    0.00339606649328079, 0.0032986815163035051, 0.003203404675755691, 
    0.0031102653044114159, 0.0030192954976240786, 0.0029305260333283259, 
    0.0028439828130090682, 0.0027596840345963901, 0.0026776382118187145, 
    0.002597843061631259, 0.0025202852007487724, 0.0024449405302191668, 
    0.0023717751468667141, 0.0023007466032535229, 0.0022318053422419881, 
    0.0021648961550324503, 0.0020999595478977274, 0.0020369329468489347, 
    0.001975751714741117, 0.0019163499956115489, 0.0018586614309839804, 
    0.0018026198087231649, 0.0017481597052315878, 0.0016952171672847181, 
    0.0016437304539870024, 0.001593640827538321, 0.0015448933501834372, 
    0.0014974376203102714, 0.0014512283684136379, 0.0014062258365712338, 
    0.0013623958833525684, 0.0013197097868814969, 0.0012781437567845834, 
    0.001237678204139581, 0.0011982968502528919, 0.0011599857742667528, 
    0.0011227325026877022, 0.0010865252304157074, 0.0010513522353296589, 
    0.0010172015121100147, 0.00098406061245085732, 0.00095191664504075998, 
    0.00092075636548668107, 0.00089056627737028817, 0.00086133267177832559, 
    0.00083304155207613499, 0.00080567841926389887, 0.00077922792544352429, 
    0.00075367343290378157, 0.00072899653901598721, 0.00070517663901473085, 
    0.00068219059835541139, 0.00066001259436293221, 0.00063861416580908881, 
    0.00061796448264277788, 0.00059803082064276744, 0.00057877920137954083, 
    0.00056017513985067401, 0.00054218443254820561, 0.00052477391814122383, 
    0.00050791215065476775, 0.00049156993911034458, 0.00047572072546953878, 
    0.00046034079154769767, 0.00044540930272596595, 0.00043090820976849183, 
    0.00041682203867872788, 0.00040313760204805683, 0.00038984366434353295, 
    0.00037693058923425366, 0.00036438999086693338, 0.00035221440444932803, 
    0.00034039698578090262, 0.000328931245200158, 0.00031781081898613685, 
    0.00030702928026342537, 0.00029657999130496953, 0.00028645599907366936, 
    0.00027664997526164939, 0.0002671542006009636, 0.0002579605908141321, 
    0.00024906075857096017, 0.00024044610280612733, 0.00023210791441504261, 
    0.00022403748630050866, 0.00021622621636574208, 0.00020866569437736328, 
    0.00020134776731060058, 0.00019426458217887703, 0.0001874086095867237, 
    0.00018077265447056089, 0.00017434986202359681, 0.00016813372630200991, 
    0.00016211810656672739, 0.00015629725255073538, 0.00015066583540492844, 
    0.00014521897708090635, 0.00013995226831073644, 0.00013486176483626006, 
    0.00012994395338964838, 0.00012519568290934681, 0.0001206140619029649, 
    0.00011619632873208907, 0.00011193970675772179, 0.00010784125972987204, 
    0.00010389776382474473, 0.00010010561108893909, 9.6460755001722621e-05, 
    9.2958703126219574e-05, 8.9594555393839829e-05, 8.6363080561715935e-05, 
    8.3258818788040361e-05, 8.0276195782647e-05, 7.7409633894372408e-05, 
    7.465364764699035e-05, 7.2002915102686071e-05, 6.9452321237147639e-05, 
    6.6996974375411499e-05, 6.4632200859509486e-05, 6.235352589380446e-05, 
    6.0156649632526773e-05, 5.8037427034162894e-05, 5.5991858089678807e-05, 
    5.4016092209431848e-05, 5.2106447398424493e-05, 5.025944191303093e-05, 
    4.8471833825639798e-05, 4.674066260589828e-05, 4.5063286552047023e-05, 
    4.3437410582586658e-05, 4.1861100302327341e-05, 4.0332780077476321e-05, 
    3.8851214767911799e-05, 3.741547648126166e-05, 3.6024899027966526e-05, 
    3.4679023560236347e-05, 3.3377539168296939e-05, 3.2120222060575471e-05, 
    3.0906876504537663e-05, 2.9737280099122261e-05, 2.8611135325468294e-05, 
    2.7528028773237659e-05, 2.648739901220808e-05, 2.5488513765111309e-05, 
    2.4530456796707289e-05, 2.3612124702805482e-05, 2.2732233506359883e-05, 
    2.1889334609689372e-05, 2.1081839213691775e-05, 2.0308049829820465e-05, 
    1.956619704243894e-05, 1.8854479301093951e-05, 1.8171103305563332e-05, 
    1.751432253696499e-05, 1.6882471702368451e-05, 1.6273995274876212e-05, 
    1.5687468874061797e-05, 1.5121612867363917e-05, 1.457529820300124e-05, 
    1.4047545036329543e-05, 1.3537515135599617e-05, 1.3044499323182201e-05, 
    1.2567901329049474e-05, 1.2107219424777277e-05, 1.1662027105543346e-05, 
    1.123195392885625e-05, 1.0816667434781587e-05, 1.0415856881440101e-05, 
    1.0029219342381973e-05, 9.6564485279509172e-06, 9.2972265105922661e-06, 
    8.9512183511433401e-06, 8.6180694470424409e-06, 8.2974052628281401e-06, 
    7.9888329769376907e-06, 7.6919445008056453e-06, 7.4063203111735327e-06, 
    7.1315335852621698e-06, 6.8671542353819951e-06, 6.6127525835383522e-06, 
    6.3679025735571931e-06, 6.1321845572825051e-06, 5.9051877898876697e-06, 
    5.6865128095966202e-06, 5.4757738578692215e-06, 5.2726014251477197e-06, 
    5.0766449064602064e-06, 4.8875752443825141e-06, 4.70508735142237e-06, 
    4.528902057938195e-06, 4.3587673373816858e-06, 4.1944586151427121e-06, 
    4.0357780613847888e-06, 3.882552881500397e-06, 3.7346327309244235e-06, 
    3.5918864724032393e-06, 3.4541985511333224e-06, 3.3214652781026209e-06, 
    3.1935912877767115e-06, 3.0704863794238243e-06, 2.9520628760634975e-06, 
    2.8382335533281044e-06, 2.7289101165194409e-06, 2.6240021453514147e-06, 
    2.5234163887622001e-06, 2.4270562765090162e-06, 2.3348215193370021e-06, 
    2.2466076900925946e-06, 2.1623057112238768e-06, 2.0818012137013596e-06, 
    2.0049737759287366e-06, 1.9316960933583197e-06, 1.8618331682716824e-06, 
    1.7952416386792646e-06, 1.7317693835869325e-06, 1.6712555434056968e-06, 
    1.6135310783529842e-06, 1.5584199520816573e-06, 1.5057409762448487e-06, 
    1.4553102874571143e-06, 1.4069443601933412e-06, 1.3604633948380439e-06, 
    1.3156948698510336e-06, 1.2724770168759576e-06, 1.2306619737193149e-06, 
    1.1901183919252195e-06, 1.1507333216469931e-06, 1.1124132588962849e-06, 
    1.075084311887464e-06, 1.0386915134594696e-06, 1.0031973685971675e-06, 
    9.6857977237100236e-07, 9.3482946258537629e-07, 9.0194718162654216e-07, 
    8.6994071777800699e-07, 8.3882198034976513e-07, 8.0860424194712038e-07, 
    7.7929965777989206e-07, 7.5091715033118675e-07, 7.2346072765712455e-07, 
    6.9692828563688276e-07, 6.7131092550411384e-07, 6.4659279751232492e-07, 
    6.2275145669030853e-07, 5.9975868896404422e-07, 5.7758173585615952e-07, 
    5.5618481790864025e-07, 5.3553083404806355e-07, 5.1558310119364675e-07, 
    4.9630699770914974e-07, 4.7767138770477817e-07, 4.5964972853199533e-07, 
    4.4222079882311367e-07, 4.2536902279507134e-07, 4.090844039160008e-07, 
    3.933621111106179e-07, 3.7820178105836945e-07, 3.6360660830064713e-07, 
    3.4958229315271818e-07, 3.3613590758544357e-07, 3.232747270013596e-07, 
    3.1100506411683085e-07, 2.99331134995611e-07, 2.8825398686528308e-07, 
    2.7777052358831364e-07, 2.6787267389428779e-07, 2.5854675688931046e-07, 
    2.4977310355940314e-07, 2.4152598938835214e-07, 2.3377391850358547e-07, 
    2.2648027527044004e-07, 2.1960432624311739e-07, 2.1310251943413446e-07, 
    2.0692999350740658e-07, 2.0104218367297385e-07, 1.9539639728076958e-07, 
    1.8995323433249038e-07, 1.8467774550415375e-07, 1.7954025128967073e-07, 
    1.7451678498131394e-07, 1.6958916433588595e-07, 1.6474473447973638e-07, 
    1.5997585366215935e-07, 1.5527920897373673e-07, 1.5065505105420375e-07, 
    1.461064251719483e-07, 1.416384554687339e-07, 1.3725771313103546e-07, 
    1.3297167433397084e-07, 1.2878825330035798e-07, 1.247153842908244e-07, 
    1.2076062399126226e-07, 1.1693075312720984e-07, 1.132313696834871e-07, 
    1.0966648343445192e-07, 1.0623813756733871e-07, 1.0294609545015029e-07, 
    9.9787635236664373e-08, 9.6757492123590083e-08, 9.3847976585175689e-08, 
    9.1049279880295947e-08, 8.8349957197516698e-08, 8.5737557997430282e-08, 
    8.3199355038268466e-08, 8.0723111383950036e-08, 7.8297819332902195e-08, 
    7.5914347968069947e-08, 7.3565945502277274e-08, 7.1248558013810028e-08, 
    6.8960944551273143e-08, 6.6704588376627683e-08, 6.4483422106643967e-08, 
    6.2303399753708052e-08, 6.0171958853649199e-08, 5.8097421417069725e-08, 
    5.6088382417993457e-08, 5.415313041898229e-08, 5.2299136919174811e-08, 
    5.0532641139491359e-08, 4.8858345644348313e-08, 4.7279227593909577e-08, 
    4.579646067662759e-08, 4.4409435562693093e-08, 4.3115861613753899e-08, 
    4.1911930752441101e-08, 4.0792524546803013e-08, 3.975144824063097e-08, 
    3.8781678954509536e-08, 3.7875619522421304e-08, 3.7025352774699975e-08, 
    3.6222893561326056e-08, 3.5460436180893628e-08, 3.473059398595727e-08, 
    3.4026625228002953e-08, 3.3342636347613923e-08, 3.2673750859202294e-08, 
    3.2016230678103232e-08, 3.1367536950734765e-08, 3.0726320477466149e-08, 
    3.0092336831140131e-08, 2.9466288340707588e-08, 2.8849602665166436e-08, 
    2.8244165280810892e-08, 2.765202873451275e-08, 2.7075125054705993e-08, 
    2.6515007562291763e-08, 2.5972645444954586e-08, 2.5448288302016496e-08, 
    2.4941410126365321e-08, 2.4450733177166916e-08, 2.3974323975133397e-08, 
    2.3509746361175678e-08, 2.3054252052743167e-08, 2.260498682652058e-08, 
    2.2159191333800304e-08, 2.1714378356716272e-08, 2.126847326797142e-08, 
    2.0819909802778276e-08, 2.0367679186492291e-08, 1.9911335371040827e-08, 
    1.9450963125957185e-08, 1.8987117794359202e-08, 1.8520746468912221e-08, 
    1.8053099614443118e-08, 1.7585640838094374e-08, 1.7119960293381393e-08, 
    1.6657695327283411e-08, 1.6200459905261708e-08, 1.5749783336901795e-08, 
    1.5307057888564969e-08, 1.4873495086579986e-08, 1.4450090700145927e-08, 
    1.4037599280240668e-08, 1.3636519559987456e-08, 1.3247092658781594e-08, 
    1.2869314832204625e-08, 1.2502966120863375e-08, 1.2147655074074649e-08, 
    1.1802878405846892e-08, 1.1468092571067964e-08, 1.1142792793171946e-08, 
    1.0826593384639292e-08, 1.051930259080419e-08, 1.0220984663060299e-08, 
    9.932002625209608e-09, 9.6530362552576307e-09, 9.3850719743296317e-09, 
    9.1293634673987709e-09, 8.8873646765121296e-09, 8.6606391042493886e-09, 
    8.4507517481798289e-09, 8.2591513114560163e-09, 8.0870514233694038e-09, 
    7.9353194020785217e-09, 7.8043805905696303e-09, 7.6941447083355626e-09, 
    7.6039590424536916e-09, 7.5325910821649064e-09, 7.4782413643568586e-09, 
    7.4385852893476795e-09, 7.4108414405566688e-09, 7.3918626013306633e-09, 
    7.3782452652370759e-09, 7.3664527790125642e-09, 7.3529472842516263e-09, 
    7.3343252236462267e-09, 7.3074512642100973e-09, 7.2695850119344006e-09, 
    7.2184948941576137e-09, 7.1525532469323919e-09, 7.0708070016301445e-09, 
    6.9730186636201442e-09, 6.8596735450984371e-09, 6.7319506677268704e-09, 
    6.5916570827215919e-09, 6.4411277226632844e-09, 6.2830958395886224e-09, 
    6.1205414330425345e-09, 5.9565273718528502e-09, 5.7940340910758848e-09, 
    5.6358043394104194e-09, 5.484208554869953e-09, 5.3411399641368273e-09, 
    5.2079456879917846e-09, 5.0853972321586652e-09, 4.9737001152938341e-09, 
    4.8725393284065564e-09, 4.7811544069117156e-09, 4.6984361150535375e-09, 
    4.6230354730637981e-09, 4.553476025684704e-09, 4.4882608223599011e-09, 
    4.4259673272258356e-09, 4.3653251982285737e-09, 4.3052741881409664e-09, 
    4.245001243868181e-09, 4.1839577500707341e-09, 4.1218589320690943e-09, 
    4.0586684291361354e-09, 3.9945711499560951e-09, 3.9299376813879402e-09, 
    3.8652830580550065e-09, 3.8012225585443384e-09, 3.7384265645816205e-09, 
    3.6775764650126607e-09, 3.6193231524403781e-09, 3.5642497928028586e-09, 
    3.512840197267909e-09, 3.4654542906166608e-09, 3.4223117015546542e-09, 
    3.3834844446883434e-09, 3.3488989489185378e-09, 3.3183473237359231e-09, 
    3.2915068796888317e-09, 3.2679664647653815e-09, 3.2472573643583646e-09, 
    3.2288863095394133e-09, 3.2123677129524347e-09, 3.1972524980734495e-09, 
    3.1831510350524071e-09, 3.1697484347871717e-09, 3.1568110576848536e-09, 
    3.1441841381063574e-09, 3.1317811210810632e-09, 3.1195663417145581e-09, 
    3.1075331028835575e-09, 3.0956798493646659e-09, 3.0839870399590871e-09, 
    3.0723974206614243e-09, 3.060801744834414e-09, 3.0490315826925475e-09, 
    3.0368598954089054e-09, 3.0240093732618569e-09, 3.0101675893344079e-09, 
    2.995007478797719e-09, 2.9782109549701739e-09, 2.9594934410185651e-09, 
    2.938626808807267e-09, 2.9154586985942841e-09, 2.8899263879256974e-09, 
    2.8620641741750979e-09, 2.8320036696880517e-09, 2.7999672988452002e-09, 
    2.7662556192365233e-09, 2.7312298032923933e-09, 2.6952906814283939e-09, 
    2.658856118990092e-09, 2.6223382973675185e-09, 2.5861225055664674e-09, 
    2.5505486282383625e-09, 2.5158964604445917e-09, 2.4823754281860578e-09, 
    2.450119161935035e-09, 2.419184904456059e-09, 2.3895575898037741e-09, 
    2.3611580192036848e-09, 2.3338544804167893e-09, 2.3074768283078384e-09, 
    2.2818320878530008e-09, 2.2567203985922963e-09, 2.2319503401333227e-09, 
    2.2073525884078543e-09, 2.1827911987679476e-09, 2.1581718376085503e-09, 
    2.1334467752261567e-09, 2.108616454498258e-09, 2.0837279506082904e-09, 
    2.0588705808205678e-09, 2.0341692970985275e-09, 2.0097763772681248e-09, 
    1.9858621222193598e-09, 1.9626050926838243e-09, 1.9401825325565925e-09, 
    1.9187613599365234e-09, 1.8984902467893516e-09, 1.8794929856880894e-09, 
    1.8618634743778623e-09, 1.8456623477672693e-09, 1.8309153549695196e-09, 
    1.8176133169890198e-09, 1.8057135646627502e-09, 1.7951424915377771e-09, 
    1.7857990024329697e-09, 1.7775584318840245e-09, 1.7702767141800599e-09, 
    1.7637944714463642e-09, 1.7579409489949211e-09, 1.7525376807985989e-09, 
    1.7474019654908516e-09, 1.7423501563885578e-09, 1.7372009993615697e-09, 
    1.731778973779177e-09, 1.7259177977361526e-09, 1.7194639450328108e-09, 
    1.7122801817688354e-09, 1.7042488597234331e-09, 1.6952748387997017e-09, 
    1.6852877608528663e-09, 1.6742436049200059e-09, 1.6621252998876884e-09, 
    1.6489424821684473e-09, 1.6347303272221019e-09, 1.6195476759689674e-09, 
    1.6034745022978389e-09, 1.5866090361928419e-09, 1.5690646013056229e-09, 
    1.5509664670956941e-09, 1.5324487188925788e-09, 1.5136513680663861e-09, 
    1.4947176389255855e-09, 1.4757915136841279e-09, 1.4570154229624023e-09, 
    1.438528109549278e-09, 1.4204624784921434e-09, 1.4029434809070256e-09, 
    1.3860858607574825e-09, 1.3699918527448929e-09, 1.3547487706264497e-09, 
    1.3404266369969779e-09, 1.3270759031291759e-09, 1.3147255209052238e-09, 
    1.3033814866593541e-09, 1.2930261261526504e-09, 1.2836182341921713e-09, 
    1.2750942732901758e-09, 1.2673705953858022e-09, 1.2603467524853275e-09, 
    1.253909654776464e-09, 1.2479384577126703e-09, 1.2423097854111398e-09, 
    1.2369030541307529e-09, 1.231605474681825e-09, 1.226316499311346e-09, 
    1.2209513694781042e-09, 1.2154437013282242e-09, 1.2097468979109203e-09, 
    1.203834485412913e-09, 1.1976993547210756e-09, 1.1913521000581474e-09, 
    1.1848185304835312e-09, 1.1781366219959408e-09, 1.171352986278522e-09, 
    1.1645191500839518e-09, 1.1576877128560533e-09, 1.1509086654182062e-09, 
    1.1442259533910015e-09, 1.1376745297719144e-09, 1.1312780002768015e-09, 
    1.1250470416494976e-09, 1.1189786571860827e-09, 1.1130563883619596e-09, 
    1.1072514064290472e-09, 1.1015245067925966e-09, 1.0958288213765429e-09, 
    1.0901131297924324e-09, 1.0843254676622708e-09, 1.0784168757736615e-09, 
    1.0723449349574846e-09, 1.0660769115506648e-09, 1.0595921964323941e-09, 
    1.0528839499310131e-09, 1.0459597463778289e-09, 1.0388412302251371e-09, 
    1.0315627478179308e-09, 1.024169127239701e-09, 1.0167127040230875e-09, 
    1.0092498956970426e-09, 1.0018375397653379e-09, 9.9452932255601513e-10, 
    9.8737252585311526e-10, 9.8040538589124053e-10, 9.7365516542933403e-10, 
    9.6713713474263846e-10, 9.6085438961897865e-10, 9.547985601036098e-10, 
    9.489512004439471e-10, 9.4328580739883886e-10, 9.3777018898665802e-10, 
    9.3236907702212911e-10, 9.2704674208577187e-10, 9.2176949646355748e-10, 
    9.1650789157779582e-10, 9.1123855398989659e-10, 9.0594551965215614e-10, 
    9.0062104812956055e-10, 8.9526582452724567e-10, 8.898886167512812e-10, 
    8.8450532909711298e-10, 8.7913759499238659e-10, 8.7381094151003946e-10, 
    8.6855271791294285e-10, 8.6338989790458713e-10, 8.5834697570758343e-10, 
    8.53444079213092e-10, 8.4869549436045783e-10, 8.4410866209107291e-10, 
    8.3968375559624866e-10, 8.354137874463597e-10, 8.3128526256577582e-10, 
    8.2727922248090987e-10, 8.2337262438793818e-10, 8.1953986562975996e-10, 
    8.1575439028313866e-10, 8.119901923166584e-10, 8.082231987786331e-10, 
    8.0443241302493236e-10, 8.0060083505113455e-10, 7.9671605883416972e-10, 
    7.9277065639215786e-10, 7.8876224559747405e-10, 7.846933482712971e-10, 
    7.8057099003652115e-10, 7.7640613159908709e-10, 7.7221290626709716e-10, 
    7.6800776914916007e-10, 7.6380852533844769e-10, 7.5963338538761826e-10, 
    7.5549999610334872e-10, 7.5142457988790091e-10, 7.4742115142803587e-10, 
    7.4350088366788868e-10, 7.3967161057507171e-10, 7.3593748563962269e-10, 
    7.322987696125229e-10, 7.2875178516298558e-10, 7.2528895810644917e-10, 
    7.2189903045322092e-10, 7.1856737917827655e-10, 7.1527648857940675e-10, 
    7.1200655818706224e-10, 7.0873628222157122e-10, 7.0544374761753222e-10, 
    7.021074966732782e-10, 6.9870762881138525e-10, 6.9522697246427603e-10, 
    6.9165217897069571e-10, 6.8797470801333483e-10, 6.8419156542624931e-10, 
    6.8030576383625547e-10, 6.7632637529849956e-10, 6.7226821113047298e-10, 
    6.6815104477819598e-10, 6.6399848488027621e-10, 6.5983649128454867e-10, 
    6.5569172434539467e-10, 6.5158977991271629e-10, 6.475535277873901e-10, 
    6.4360164447545057e-10, 6.3974752641750532e-10, 6.3599863140020861e-10, 
    6.3235636557216984e-10, 6.2881646064406098e-10, 6.2536987704514176e-10, 
    6.220040463875915e-10, 6.1870442882234434e-10, 6.1545613143616451e-10, 
    6.1224551698907759e-10, 6.0906158209770788e-10, 6.0589703764276758e-10, 
    6.0274896327083244e-10, 5.9961903511821175e-10, 5.9651327336301096e-10, 
    5.9344142221903275e-10, 5.9041596496717544e-10, 5.8745093357568866e-10, 
    5.8456057052268918e-10, 5.8175800523835703e-10, 5.7905399760682805e-10, 
    5.764558938806927e-10, 5.7396681453065029e-10, 5.7158518847094192e-10, 
    5.6930458815047964e-10, 5.6711394618392202e-10, 5.6499805388662889e-10, 
    5.6293835976054678e-10, 5.6091394918219879e-10, 5.5890266698962506e-10, 
    5.5688224170860524e-10, 5.5483138859752026e-10, 5.5273073769135432e-10, 
    5.5056360382722078e-10, 5.4831648640509033e-10, 5.4597936372340821e-10, 
    5.4354572793284593e-10, 5.4101247154222171e-10, 5.3837960012494815e-10, 
    5.3564990836825567e-10, 5.3282860519683693e-10, 5.299229894685608e-10, 
    5.2694213766730628e-10, 5.2389668833848e-10, 5.2079861723933243e-10, 
    5.1766107502723025e-10, 5.144981693887477e-10, 5.1132473364063066e-10, 
    5.081559953229194e-10, 5.0500719408937631e-10, 5.0189310428060235e-10, 
    4.9882754067810429e-10, 4.9582281687416553e-10, 4.9288927530291211e-10, 
    4.9003486455718548e-10, 4.8726487751453066e-10, 4.8458179697518739e-10, 
    4.8198535594750137e-10, 4.7947272290119953e-10, 4.7703887486629007e-10, 
    4.7467705364475439e-10, 4.7237931821483872e-10, 4.7013710167241713e-10, 
    4.6794177200472129e-10, 4.6578508816238926e-10, 4.6365959199193044e-10, 
    4.6155885674184118e-10, 4.5947762967876957e-10, 4.5741182144124379e-10, 
    4.5535842738662972e-10, 4.5331532647991018e-10, 4.5128106200142076e-10, 
    4.4925455728983058e-10, 4.4723485360631118e-10, 4.4522085322840549e-10, 
    4.4321111898881899e-10, 4.4120368640604968e-10, 4.3919597739075474e-10, 
    4.3718475105319277e-10, 4.3516615579238748e-10, 4.3313581156628806e-10, 
    4.3108901458745645e-10, 4.290209505773937e-10, 4.2692700707379581e-10, 
    4.2480306664160406e-10, 4.2264585702832645e-10, 4.2045321822981297e-10, 
    4.1822436465679753e-10, 4.1596004254398622e-10, 4.1366260968045159e-10, 
    4.113359810377876e-10, 4.0898550984482341e-10, 4.0661773602484884e-10, 
    4.042401120002797e-10, 4.0186064494919532e-10, 3.9948756817479456e-10, 
    3.9712899838474663e-10, 3.94792665274661e-10, 3.9248566282314102e-10, 
    3.9021430089664095e-10, 3.8798399011489888e-10, 3.8579922129290237e-10, 
    3.8366356775617372e-10, 3.8157977546498937e-10, 3.7954984813607536e-10, 
    3.7757520167401418e-10, 3.7565680299430499e-10, 3.7379533233157412e-10, 
    3.7199130425743681e-10, 3.7024517731455568e-10, 3.6855737221170269e-10, 
    3.6692824607375481e-10, 3.6535795549811054e-10, 3.6384626929527083e-10, 
    3.6239226773865003e-10, 3.6099405866940197e-10, 3.5964844197608643e-10, 
    3.5835067354701312e-10, 3.570942697678134e-10, 3.5587100236669188e-10, 
    3.5467099451948382e-10, 3.5348303058424941e-10, 3.5229498372133724e-10, 
    3.5109438758722121e-10, 3.4986903302515204e-10, 3.4860761524829762e-10, 
    3.4730028300542493e-10, 3.4593911387067769e-10, 3.4451840237010037e-10, 
    3.4303481850800091e-10, 3.4148736638016096e-10, 3.3987723848613621e-10, 
    3.3820752088023053e-10, 3.3648289100894653e-10, 3.3470926894378159e-10, 
    3.3289354340009021e-10, 3.3104332582979171e-10, 3.2916681749054853e-10, 
    3.2727272585647339e-10, 3.253702595464774e-10, 3.2346910757423049e-10, 
    3.2157944516819043e-10, 3.1971183151991125e-10, 3.1787707793428781e-10, 
    3.160859820010936e-10, 3.1434900945239893e-10, 3.1267587357617042e-10, 
    3.1107513328359399e-10, 3.0955376579394367e-10, 3.0811684609125453e-10, 
    3.0676729517920394e-10, 3.0550578899385863e-10, 3.0433077107015069e-10, 
    3.032386200712497e-10, 3.0222386492431186e-10, 3.0127949480598731e-10, 
    3.0039722887686867e-10, 2.9956779518135002e-10, 2.9878110244907925e-10, 
    2.9802639819607195e-10, 2.9729232537000681e-10, 2.9656701367257191e-10, 
    2.9583813762809265e-10, 2.9509309045899117e-10, 2.943192391886144e-10, 
    2.9350432963844305e-10, 2.9263698169427757e-10, 2.9170733016769284e-10, 
    2.907076606651704e-10, 2.896330646752731e-10, 2.884819620257156e-10, 
    2.8725647314415827e-10, 2.859625223243413e-10, 2.8460969977607597e-10, 
    2.8321080755778138e-10, 2.8178117093591978e-10, 2.8033770640782113e-10, 
    2.7889788371822049e-10, 2.7747859389222437e-10, 2.7609508609321284e-10, 
    2.7476000086123733e-10, 2.7348262492805838e-10, 2.7226835203007216e-10, 
    2.711184747924101e-10, 2.700302229131259e-10, 2.6899711990085774e-10, 
    2.6800955811294702e-10, 2.670556044521385e-10, 2.6612193172813604e-10, 
    2.6519485399306002e-10, 2.642613524549473e-10, 2.6331006797194938e-10, 
    2.6233214733398864e-10, 2.6132193907913657e-10, 2.602774312553954e-10, 
    2.5920047836521815e-10, 2.5809670442576385e-10, 2.5697519857562926e-10, 
    2.5584792644917433e-10, 2.5472896532470406e-10, 2.5363358719414965e-10, 
    2.5257726483697029e-10, 2.5157463476692269e-10, 2.5063854555559386e-10, 
    2.4977918216208299e-10, 2.4900338343376706e-10, 2.4831412667242304e-10, 
    2.4771028681668973e-10, 2.471865909896526e-10, 2.4673386238016482e-10, 
    2.4633945787840407e-10, 2.4598793069287329e-10, 2.4566184014003773e-10, 
    2.4534268931530594e-10, 2.4501190512947178e-10, 2.4465183618652838e-10, 
    2.4424665848904849e-10, 2.4378318771437781e-10, 2.4325148969973207e-10, 
    2.4264530587365923e-10, 2.4196221657788109e-10, 2.4120359097137341e-10, 
    2.4037427874877053e-10, 2.3948213626784276e-10, 2.3853737600290637e-10, 
    2.3755184119040844e-10, 2.3653822855114825e-10, 2.3550935416084519e-10, 
    2.3447747817710568e-10, 2.334537668998302e-10, 2.3244787796888432e-10, 
    2.3146771479616182e-10, 2.3051930453544813e-10, 2.2960681815062528e-10, 
    2.2873266796192341e-10, 2.2789767471769294e-10, 2.2710125172142136e-10, 
    2.2634160434859853e-10, 2.2561588288307753e-10, 2.2492033121967038e-10, 
    2.2425037136956503e-10, 2.2360068232776518e-10, 2.2296522738960279e-10, 
    2.2233730116196164e-10, 2.217095527866962e-10, 2.2107405561577805e-10, 
    2.2042237923621852e-10, 2.1974573968407384e-10, 2.1903518410678541e-10, 
    2.1828186445600757e-10, 2.1747735791390631e-10, 2.1661408821317183e-10, 
    2.1568577260950506e-10, 2.1468793090302167e-10, 2.1361837526468485e-10, 
    2.1247767690754284e-10, 2.1126951225432207e-10, 2.1000089182450099e-10, 
    2.0868216893907575e-10, 2.07326833503201e-10, 2.059510550529843e-10, 
    2.0457297840005298e-10, 2.0321182471491833e-10, 2.0188683930619021e-10, 
    2.0061616221987057e-10, 1.9941574566182598e-10, 1.9829836512960717e-10, 
    1.97272865746e-10, 1.9634367642208102e-10, 1.9551066308550269e-10, 
    1.9476930657997866e-10, 1.9411121668060601e-10, 1.9352488928905779e-10, 
    1.9299666504038605e-10, 1.9251175671174872e-10, 1.9205527528894256e-10, 
    1.9161313982838042e-10, 1.9117282071389983e-10, 1.9072382314539651e-10, 
    1.9025795694435132e-10, 1.8976934290428176e-10, 1.8925423753461813e-10, 
    1.8871069686729282e-10, 1.8813816334628587e-10, 1.8753703018108802e-10, 
    1.8690823674044353e-10, 1.8625292700584281e-10, 1.8557221398398711e-10, 
    1.848670288313466e-10, 1.8413808114091835e-10, 1.8338588816877072e-10, 
    1.8261088650791959e-10, 1.8181358056651433e-10, 1.8099473457895309e-10, 
    1.8015557926683344e-10, 1.7929802904303519e-10, 1.7842486813536096e-10, 
    1.7753991980519291e-10, 1.7664813510944752e-10, 1.7575560193814072e-10, 
    1.7486943364157544e-10, 1.7399753637636257e-10, 1.7314822468322236e-10, 
    1.7232974544073493e-10, 1.7154969623099414e-10, 1.7081444711346655e-10, 
    1.7012856569250036e-10, 1.6949437915460233e-10, 1.6891168736018208e-10, 
    1.6837770180601715e-10, 1.6788720011910141e-10, 1.6743290598421555e-10, 
    1.6700603664674627e-10, 1.6659696139330698e-10, 1.6619586916022715e-10, 
    1.6579340441549792e-10, 1.6538115865375027e-10, 1.6495201539957786e-10, 
    1.6450030669817664e-10, 1.6402182767013098e-10, 1.6351372481676849e-10, 
    1.6297435620813654e-10, 1.624031438320459e-10, 1.6180050424411199e-10, 
    1.6116786710870796e-10, 1.6050778557319365e-10, 1.5982409417974102e-10, 
    1.5912209811242943e-10, 1.5840865308744479e-10, 1.5769215311471436e-10, 
    1.5698230355506389e-10, 1.5628969503342507e-10, 1.5562516294840917e-10, 
    1.5499900282076341e-10, 1.5442008256800324e-10, 1.5389499302978546e-10, 
    1.5342730538161923e-10, 1.5301706030182429e-10, 1.5266053850428374e-10, 
    1.5235038171679434e-10, 1.5207603742164522e-10, 1.5182451642617322e-10, 
    1.5158135618635742e-10, 1.5133173297441982e-10, 1.5106156397976653e-10, 
    1.5075854009825093e-10, 1.5041295635268422e-10, 1.5001829645202248e-10, 
    1.4957152151035539e-10, 1.4907306323663836e-10, 1.4852654827593484e-10, 
    1.4793830269963523e-10, 1.4731668721648187e-10, 1.4667135596561829e-10, 
    1.4601248293414592e-10, 1.4535003592076932e-10, 1.4469311434024208e-10, 
    1.4404941905452546e-10, 1.4342484257960186e-10, 1.4282321172817547e-10, 
    1.4224616046285807e-10, 1.4169315769271326e-10, 1.4116163705085185e-10, 
    1.4064726692850492e-10, 1.4014429910030147e-10, 1.3964599544996821e-10, 
    1.3914510094026468e-10, 1.3863432204745981e-10, 1.3810677702363288e-10, 
    1.375563939996824e-10, 1.3697819485949937e-10, 1.3636848415811983e-10, 
    1.3572489497898707e-10, 1.3504633246407851e-10, 1.3433279970700464e-10, 
    1.3358517643766215e-10, 1.328049632524755e-10, 1.3199406176068916e-10, 
    1.31154598973928e-10, 1.3028886020499977e-10, 1.2939932130377298e-10, 
    1.2848879184280489e-10, 1.2756062813060564e-10, 1.2661901894855017e-10, 
    1.2566925067179896e-10, 1.2471795189078297e-10, 1.2377322632978439e-10, 
    1.2284467120095554e-10, 1.2194321747121552e-10, 1.2108081765720023e-10, 
    1.2026995633409824e-10, 1.1952304243749094e-10, 1.1885168331220513e-10, 
    1.1826594456370617e-10, 1.1777361987830681e-10, 1.1737961260150216e-10, 
    1.1708544735649809e-10, 1.1688902519472387e-10, 1.1678458549231568e-10, 
    1.1676296135619815e-10, 1.1681204072178593e-10, 1.1691746772923456e-10, 
    1.1706347091562611e-10, 1.1723378563494355e-10, 1.1741254966077359e-10, 
    1.1758513824580639e-10, 1.177388259470065e-10, 1.1786326516671392e-10, 
    1.1795072200659253e-10, 1.1799611110925747e-10, 1.1799680727995419e-10, 
    1.1795233747318026e-10, 1.1786394590072045e-10, 1.1773415724130687e-10, 
    1.1756632556805828e-10, 1.1736427599276182e-10, 1.1713198864499542e-10, 
    1.1687340575340763e-10, 1.1659226802300216e-10, 1.1629204034547994e-10, 
    1.1597582277714417e-10, 1.1564628856656234e-10, 1.1530557255379207e-10, 
    1.1495516077879006e-10, 1.1459574437199005e-10, 1.1422710837948887e-10, 
    1.1384801378015294e-10, 1.1345620521980448e-10, 1.130484582659107e-10, 
    1.1262079519762505e-10, 1.1216877525106542e-10, 1.1168793490350723e-10, 
    1.1117426190018738e-10, 1.1062474470225804e-10, 1.1003786387010994e-10, 
    1.0941404921367496e-10, 1.0875596252959002e-10, 1.0806866403189325e-10, 
    1.0735953385175789e-10, 1.0663804187580228e-10, 1.0591529817662408e-10, 
    1.0520348114569673e-10, 1.0451513344062763e-10, 1.0386245571368068e-10, 
    1.0325656487844052e-10, 1.0270689073089981e-10, 1.0222063392385039e-10, 
    1.0180244243776231e-10, 1.0145422143297408e-10, 1.0117516673263746e-10, 
    1.0096192835790274e-10, 1.0080895283323462e-10, 1.007088985835572e-10, 
    1.0065314121126919e-10, 1.0063227012891783e-10, 1.0063659485948416e-10, 
    1.0065655032746125e-10, 1.006830673695865e-10, 1.00707791931475e-10, 
    1.0072323960655822e-10, 1.0072283115815677e-10, 1.0070086535664701e-10, 
    1.0065241486595244e-10, 1.0057323269449668e-10, 1.0045961716714765e-10, 
    1.0030835966601844e-10, 1.0011670532738959e-10, 9.9882415022431613e-11, 
    9.9603850980834397e-11, 9.9280167173231619e-11, 9.8911484446063428e-11, 
    9.8499119773481661e-11, 9.8045757572704404e-11, 9.7555608996176812e-11, 
    9.7034455673507651e-11, 9.6489644275586345e-11, 9.5929947912897876e-11, 
    9.5365358436038306e-11, 9.4806755123194672e-11, 9.4265534534346211e-11, 
    9.3753141336154992e-11, 9.3280605308190223e-11, 9.2858029203499791e-11, 
    9.249412368794522e-11, 9.2195727548229432e-11, 9.1967434772408162e-11, 
    9.181125857257347e-11, 9.1726428766302855e-11, 9.1709287238643553e-11, 
    9.1753361486299018e-11, 9.1849546487695732e-11, 9.1986492993639623e-11, 
    9.2151112884742646e-11, 9.2329250776751546e-11, 9.2506412032675711e-11, 
    9.2668583717553595e-11, 9.2803012207780557e-11, 9.2898952010910693e-11, 
    9.2948248966440342e-11, 9.2945794320494813e-11, 9.2889724048035371e-11, 
    9.2781439590093083e-11, 9.2625358937355994e-11, 9.2428505080300478e-11, 
    9.2199912850527375e-11, 9.194995415773276e-11, 9.1689580249536854e-11, 
    9.1429611373528647e-11, 9.1180055288002319e-11, 9.0949552800230596e-11, 
    9.0744918710583518e-11, 9.0570858039879665e-11, 9.0429781997702062e-11, 
    9.0321797707360013e-11, 9.0244790669804282e-11, 9.0194646253735864e-11, 
    9.0165522824756971e-11, 9.0150249282833629e-11, 9.014074073343591e-11, 
    9.0128505998135348e-11, 9.0105115518902267e-11, 9.0062721158687554e-11, 
    8.9994497726552562e-11, 8.9895047641388543e-11, 8.9760671378644809e-11, 
    8.9589542115784456e-11, 8.938170154990503e-11, 8.913892897392331e-11, 
    8.88644345874378e-11, 8.8562460851390471e-11, 8.8237761985365144e-11, 
    8.7895093808464972e-11, 8.753866943964783e-11, 8.7171746564743832e-11, 
    8.6796288971806618e-11, 8.641283846702585e-11, 8.6020527808257994e-11, 
    8.5617324278118585e-11, 8.5200388804378867e-11, 8.4766608237292955e-11, 
    8.431315702491818e-11, 8.3838108203266929e-11, 8.3340928064904959e-11, 
    8.2822891707002837e-11, 8.2287292534552761e-11, 8.1739468483106071e-11, 
    8.1186557690597392e-11, 8.0637099239043621e-11, 8.0100426295056152e-11, 
    7.9585975981282942e-11, 7.9102523722061718e-11, 7.8657499513385615e-11, 
    7.8256381772896401e-11, 7.7902310699682172e-11, 7.7595900887849225e-11, 
    7.7335344369340617e-11, 7.7116726486117151e-11, 7.6934602517512968e-11, 
    7.6782701081456967e-11, 7.6654762167808048e-11, 7.6545336964360716e-11, 
    7.6450556630984153e-11, 7.6368701520297972e-11, 7.6300596677864966e-11, 
    7.6249694817792849e-11, 7.6221930883177598e-11, 7.6225257681990421e-11, 
    7.6268990097294377e-11, 7.6362913152297913e-11, 7.6516323401754258e-11, 
    7.6736995981710942e-11, 7.7030244652639496e-11, 7.7398060701775654e-11, 
    7.7838505662802657e-11, 7.8345329290498055e-11, 7.8907920802084396e-11, 
    7.9511540318123985e-11, 8.0137899349512013e-11, 8.0765977900425084e-11, 
    8.1373110577348077e-11, 8.1936178598043422e-11, 8.2432919310960397e-11, 
    8.2843158108389892e-11, 8.3149978802353877e-11, 8.3340651629029756e-11, 
    8.3407336930753486e-11, 8.3347439416005612e-11, 8.3163663308914479e-11, 
    8.2863695295461166e-11, 8.2459624708530699e-11, 8.1967056134400483e-11, 
    8.1404074472519762e-11, 8.0790070315113448e-11, 8.0144573803402495e-11, 
    7.9486111792604436e-11, 7.8831255547889975e-11, 7.8193835184050634e-11, 
    7.7584439124238821e-11, 7.7010171099202248e-11, 7.6474708565795519e-11, 
    7.5978566711249691e-11, 7.5519620118103699e-11, 7.5093723101343189e-11, 
    7.4695443187128932e-11, 7.431875129995375e-11, 7.3957691101354402e-11, 
    7.3606898160148976e-11, 7.3262006317660874e-11, 7.2919853692115852e-11, 
    7.2578580566822947e-11, 7.2237555153578971e-11, 7.1897255617968222e-11, 
    7.1559054599971527e-11, 7.1225039303962723e-11, 7.0897823364972442e-11, 
    7.0580433571479984e-11, 7.027621235517432e-11, 6.9988797887826515e-11, 
    6.9722101380835644e-11, 6.9480304823139509e-11, 6.9267798614667075e-11, 
    6.908910369591988e-11, 6.8948678801113894e-11, 6.8850682639298381e-11, 
    6.8798658993431959e-11, 6.8795199341345423e-11, 6.8841553251780715e-11, 
    6.8937320840781996e-11, 6.9080176608602653e-11, 6.926574246743455e-11, 
    6.9487550023338505e-11, 6.9737204165735948e-11, 7.0004665696840757e-11, 
    7.0278704945453278e-11, 7.0547426409865556e-11, 7.0798904447237498e-11, 
    7.1021810649351181e-11, 7.1206047285178974e-11, 7.1343275106711514e-11, 
    7.1427372300476021e-11, 7.1454723611142881e-11, 7.1424379161214152e-11, 
    7.1338038581880565e-11, 7.11998983891803e-11, 7.1016323065587792e-11, 
    7.0795429158774522e-11, 7.0546538254596948e-11, 7.0279572884024141e-11, 
    7.0004400914423052e-11, 6.9730177606670462e-11, 6.9464702505108586e-11, 
    6.9213871875653595e-11, 6.8981197085164568e-11, 6.876751343418778e-11, 
    6.8570836329130429e-11, 6.8386452140823353e-11, 6.82071821679209e-11, 
    6.8023895099450937e-11, 6.7826168360949306e-11, 6.760310567985718e-11, 
    6.734420667694548e-11, 6.704025816313337e-11, 6.6684132923661231e-11, 
    6.6271453919313876e-11, 6.5801032018498198e-11, 6.5275057847098918e-11, 
    6.4699011385485318e-11, 6.4081311880547153e-11, 6.3432705542586007e-11, 
    6.2765491960490108e-11, 6.2092622461090291e-11, 6.1426779000019552e-11, 
    6.0779491106961968e-11, 6.01604072927973e-11, 5.9576732380235246e-11, 
    5.9032926191034271e-11, 5.8530639057870348e-11, 5.8068912472395557e-11, 
    5.7644575533422338e-11, 5.7252825857016557e-11, 5.6887909223424907e-11, 
    5.654384365102825e-11, 5.6215091281447781e-11, 5.5897157659901437e-11, 
    5.5587038382023635e-11, 5.5283497170160375e-11, 5.4987148834811907e-11, 
    5.4700379083234217e-11, 5.4427068172548299e-11, 5.417220828237705e-11, 
    5.3941419091554504e-11, 5.3740409119982952e-11, 5.3574429960335953e-11, 
    5.3447768243953894e-11, 5.3363288916622019e-11, 5.3322093248185626e-11, 
    5.3323263999939752e-11, 5.3363763726581955e-11, 5.3438437064778524e-11, 
    5.354016557764878e-11, 5.3660137186762267e-11, 5.3788238465461432e-11, 
    5.3913538509399371e-11, 5.4024866664921977e-11, 5.4111422398333485e-11, 
    5.4163424664980733e-11, 5.4172734449418426e-11, 5.4133426123870573e-11, 
    5.4042264291756305e-11, 5.3899051164446411e-11, 5.3706796274369838e-11, 
    5.3471708596003562e-11, 5.3202979382380351e-11, 5.2912364033954429e-11, 
    5.2613573925240193e-11, 5.2321507050238974e-11, 5.2051367273809479e-11, 
    5.1817720563781391e-11, 5.1633537330801999e-11, 5.1509314720264878e-11, 
    5.1452312859193437e-11, 5.1465993107904488e-11, 5.1549684059210239e-11, 
    5.1698520969977466e-11, 5.1903693535436785e-11, 5.2152969118487248e-11, 
    5.2431465963832891e-11, 5.2722654420681274e-11, 5.3009481662800836e-11, 
    5.3275546152056938e-11, 5.3506225185590439e-11, 5.3689656303088327e-11, 
    5.3817488495261039e-11, 5.388533058184303e-11, 5.3892861541302428e-11, 
    5.3843585649544242e-11, 5.374427532807512e-11, 5.3604138667910623e-11, 
    5.3433810931489327e-11, 5.32442772922842e-11, 5.3045814520566842e-11, 
    5.2847085525727732e-11, 5.2654456432750046e-11, 5.2471600532410265e-11, 
    5.2299418773098061e-11, 5.213627087147793e-11, 5.1978474866729361e-11, 
    5.1820999456270361e-11, 5.1658285388310889e-11, 5.1485062471926289e-11, 
    5.1297099056560309e-11, 5.1091800489041844e-11, 5.0868580400758314e-11, 
    5.0628998137092786e-11, 5.0376656906547649e-11, 5.0116876861829738e-11, 
    4.985620527310419e-11, 4.9601822888341856e-11, 4.9360915560863872e-11, 
    4.9140070097296337e-11, 4.8944773608087555e-11, 4.8779029140781016e-11, 
    4.8645127481663929e-11, 4.8543583054505381e-11, 4.8473222414572991e-11, 
    4.8431405031977404e-11, 4.8414342901749655e-11, 4.8417495057269928e-11, 
    4.8436001380402917e-11, 4.8465118714811488e-11, 4.8500639162506767e-11, 
    4.8539245055166379e-11, 4.8578805821675548e-11, 4.8618563063805798e-11, 
    4.8659208710356452e-11, 4.8702832744703348e-11, 4.8752746832896361e-11, 
    4.8813181356819917e-11, 4.8888878978018778e-11, 4.8984605681170139e-11, 
    4.9104637876647136e-11, 4.9252252494308522e-11, 4.9429272206817898e-11, 
    4.963572558828383e-11, 4.9869643281560886e-11, 5.0127010594879344e-11, 
    5.0401903919751728e-11, 5.068676596348182e-11, 5.0972810324829367e-11, 
    5.1250512384072523e-11, 5.1510141514800122e-11, 5.1742275981622912e-11, 
    5.1938283242922016e-11, 5.2090710738021264e-11, 5.2193593930608694e-11, 
    5.2242665670551888e-11, 5.2235478598441714e-11, 5.2171453940179434e-11, 
    5.2051882576201612e-11, 5.1879877371588704e-11, 5.1660311081921407e-11, 
    5.1399716478874375e-11, 5.1106170205980934e-11, 5.0789132714747596e-11, 
    5.0459236808238627e-11, 5.0128010420979317e-11, 4.9807536523308932e-11, 
    4.9510030200779001e-11, 4.9247345120678656e-11, 4.903042881412849e-11, 
    4.8868770133204981e-11, 4.8769830951102649e-11, 4.8738545849773337e-11, 
    4.8776901357231815e-11, 4.8883633478607342e-11, 4.9054092641411335e-11, 
    4.928028280980837e-11, 4.9551083361865589e-11, 4.9852668321984929e-11, 
    5.0169095448611732e-11, 5.0483030728370619e-11, 5.0776583363234106e-11, 
    5.103220269682939e-11, 5.1233571012560176e-11, 5.1366430267457019e-11, 
    5.1419308865907448e-11, 5.1384088619176518e-11, 5.1256365773500489e-11, 
    5.1035600253053735e-11, 5.072502907123445e-11, 5.0331376737307635e-11, 
    4.986436763595306e-11, 4.9336096957365434e-11, 4.8760305280606143e-11, 
    4.8151613374853119e-11, 4.7524771928591291e-11, 4.689396857097092e-11, 
    4.6272230887890636e-11, 4.5670960617694538e-11, 4.509959924866043e-11, 
    4.4565418264537438e-11, 4.4073458130030377e-11, 4.362655783164926e-11, 
    4.322549252494963e-11, 4.2869175020220616e-11, 4.2554909917009766e-11, 
    4.2278699268640359e-11, 4.2035551337036151e-11, 4.1819802708287009e-11, 
    4.162543893729494e-11, 4.1446376706756471e-11, 4.1276726561844707e-11, 
    4.1110997421660042e-11, 4.0944232953234133e-11, 4.0772105655932291e-11, 
    4.0590921194806237e-11, 4.0397565284990095e-11, 4.0189403207787618e-11, 
    3.9964152216500841e-11, 3.9719740835322763e-11, 3.9454175001232664e-11, 
    3.9165459063697413e-11, 3.8851553310033955e-11, 3.8510401743442247e-11, 
    3.8140038890634522e-11, 3.7738746028711029e-11, 3.7305249349816208e-11, 
    3.6838963087918256e-11, 3.6340212551625664e-11, 3.5810453893410011e-11, 
    3.5252442761756625e-11, 3.467033851532564e-11, 3.4069749717562239e-11, 
    3.3457690332566761e-11, 3.2842462888110083e-11, 3.2233477963225423e-11, 
    3.1641002731137431e-11, 3.1075871114960927e-11, 3.0549145539154564e-11, 
    3.0071759579679242e-11, 2.9654147441600573e-11, 2.9305873189774712e-11, 
    2.9035267896393078e-11, 2.884910050218133e-11, 2.8752284144033778e-11, 
    2.8747641777663393e-11, 2.8835745121003389e-11, 2.9014841195670192e-11, 
    2.9280869637043519e-11, 2.9627596745225794e-11, 3.0046838183365455e-11, 
    3.0528791975680804e-11, 3.1062437616676962e-11, 3.1635994669342804e-11, 
    3.2237407930530619e-11, 3.2854817746999253e-11, 3.3476977967358888e-11, 
    3.4093596434703352e-11, 3.4695570164823055e-11, 3.5275097350353434e-11, 
    3.5825647941799658e-11, 3.6341835173869029e-11, 3.68191826200401e-11, 
    3.7253845275860731e-11, 3.7642315349694951e-11, 3.7981165504354122e-11, 
    3.8266875348406987e-11, 3.8495773282127654e-11, 3.8664111283002011e-11, 
    3.876828148466955e-11, 3.880514224721923e-11, 3.8772436610112267e-11, 
    3.8669235006746832e-11, 3.8496356206809674e-11, 3.8256707351684476e-11, 
    3.7955490232400062e-11, 3.7600227527971652e-11, 3.7200620706527409e-11, 
    3.6768204199779372e-11, 3.6315853298127254e-11, 3.585716168188857e-11, 
    3.5405754480233251e-11, 3.4974598930520889e-11, 3.4575349438893052e-11, 
    3.4217788090487848e-11, 3.3909410394573693e-11, 3.3655138579680064e-11, 
    3.3457212374592798e-11, 3.3315229271414502e-11, 3.3226311921425165e-11, 
    3.3185394489584463e-11, 3.3185589988983975e-11, 3.3218608802267258e-11, 
    3.3275218696409768e-11, 3.3345696847138843e-11, 3.3420285488054904e-11, 
    3.3489602363508981e-11, 3.3545016600582912e-11, 3.3578973105760544e-11, 
    3.3585239881288954e-11, 3.3559091499522995e-11, 3.3497415225929561e-11, 
    3.3398731697307376e-11, 3.3263152974878649e-11, 3.3092270386069481e-11, 
    3.2889000734814233e-11, 3.2657388136317676e-11, 3.2402400054671419e-11, 
    3.2129725490925812e-11, 3.1845598573749324e-11, 3.1556617582422171e-11, 
    3.1269628380800929e-11, 3.0991604072776613e-11, 3.0729551347375441e-11, 
    3.0490410598218712e-11, 3.0280947775394907e-11, 3.0107607460780684e-11, 
    2.9976342186033267e-11, 2.9892387494078936e-11, 2.9860014460845509e-11, 
    2.9882235339622622e-11, 2.996052600749569e-11, 3.0094543794071528e-11, 
    3.02818984096359e-11, 3.0518003396816259e-11, 3.0796025040247965e-11, 
    3.1106950842596933e-11, 3.143981723177986e-11, 3.1782077143010574e-11, 
    3.2120124444714594e-11, 3.2439921352050802e-11, 3.2727751018704577e-11, 
    3.2970983500122887e-11, 3.3158854870153404e-11, 3.3283172263108358e-11, 
    3.3338899053519318e-11, 3.332453116458989e-11, 3.3242284054905735e-11, 
    3.3098009941403064e-11, 3.2900879951470065e-11, 3.2662820200747939e-11, 
    3.2397775383703011e-11, 3.2120827422665047e-11, 3.1847262264985798e-11, 
    3.1591647243684208e-11, 3.1367002180126435e-11, 3.1184107211284484e-11, 
    3.1051021909098002e-11, 3.0972820116067538e-11, 3.0951548987788898e-11, 
    3.0986414494822673e-11, 3.1074153263019358e-11, 3.1209522927850868e-11, 
    3.1385916955457419e-11, 3.15960021603707e-11, 3.1832360210977488e-11, 
    3.2088069199016456e-11, 3.2357216451308114e-11, 3.2635279612069663e-11, 
    3.2919393199237171e-11, 3.3208455397577086e-11, 3.3503104373782364e-11, 
    3.380552114082011e-11, 3.411913542339531e-11, 3.4448175249085913e-11, 
    3.4797159419488298e-11, 3.5170328531126049e-11, 3.5571070057029421e-11, 
    3.6001384209697888e-11, 3.6461448600667268e-11, 3.6949309064619421e-11, 
    3.7460758547571268e-11, 3.7989404990526651e-11, 3.8526961749221572e-11, 
    3.9063707840810171e-11, 3.9589126558387635e-11, 4.0092644973672168e-11, 
    4.0564418388809375e-11, 4.099606376873498e-11, 4.138130763047742e-11, 
    4.1716435277788022e-11, 4.2000524403462128e-11, 4.2235419690281251e-11, 
    4.2425454418081957e-11, 4.2576925989657838e-11, 4.2697395868913697e-11, 
    4.2794870557157895e-11, 4.2876951411176195e-11, 4.2950017901901047e-11, 
    4.301855512991827e-11, 4.308464550905391e-11, 4.3147711847220114e-11, 
    4.3204487781562056e-11, 4.3249246507849266e-11, 4.3274233497009323e-11, 
    4.3270277921589063e-11, 4.3227507735659118e-11, 4.3136127906060613e-11, 
    4.298717997179115e-11, 4.2773242665237521e-11, 4.2489015163255713e-11, 
    4.2131761685267694e-11, 4.1701575926572179e-11, 4.1201479208903938e-11, 
    4.063731816080765e-11, 4.0017515680943483e-11, 3.9352652046961122e-11, 
    3.8654935993505272e-11, 3.7937570840678113e-11, 3.7214075873729794e-11, 
    3.6497600643309588e-11, 3.5800270775085381e-11, 3.5132607811661901e-11, 
    3.4503090732604973e-11, 3.3917848329187294e-11, 3.3380562198417125e-11, 
    3.2892541256147853e-11, 3.2453000920214988e-11, 3.205949682485492e-11, 
    3.170849680609882e-11, 3.1396014199968098e-11, 3.111826950384843e-11, 
    3.0872281678878694e-11, 3.0656358997970169e-11, 3.0470429303591267e-11, 
    3.0316165920945808e-11, 3.0196915283686088e-11, 3.0117413730509198e-11, 
    3.0083348521853167e-11, 3.0100790641968478e-11, 3.0175539215097787e-11, 
    3.0312474782551062e-11, 3.0514945498646999e-11, 3.0784238028500133e-11, 
    3.1119181094926637e-11, 3.151588635657112e-11, 3.1967643620118335e-11, 
    3.2464976511243508e-11, 3.2995827373527258e-11, 3.3545882497191581e-11, 
    3.409901085560137e-11, 3.4637809394067452e-11, 3.5144219907123263e-11, 
    3.5600232442976385e-11, 3.5988640774590757e-11, 3.6293830534357124e-11, 
    3.6502555999407634e-11, 3.660468937759235e-11, 3.6593893410896455e-11, 
    3.6468151508366241e-11, 3.6230115063258924e-11, 3.5887235615348555e-11, 
    3.5451616823531576e-11, 3.4939589353241548e-11, 3.4371008033947118e-11, 
    3.3768279523366543e-11, 3.3155174952966082e-11, 3.255550574769775e-11, 
    3.1991742236270217e-11, 3.1483676872687967e-11, 3.1047230413736875e-11, 
    3.0693504762384181e-11, 3.0428156788685605e-11, 3.025115198982315e-11, 
    3.0156910094851853e-11, 3.0134861622940535e-11, 3.0170334505564761e-11, 
    3.0245723506012494e-11, 3.0341849996084428e-11, 3.0439372052329623e-11, 
    3.0520165222578567e-11, 3.0568547056848335e-11, 3.0572260161558025e-11, 
    3.0523161678616109e-11, 3.041756694440441e-11, 3.0256258179501294e-11, 
    3.0044173701088598e-11, 2.9789830283747707e-11, 2.9504539226541891e-11, 
    2.9201493380885675e-11, 2.8894798171789103e-11, 2.8598516739416859e-11, 
    2.8325793015039021e-11, 2.8088101720794448e-11, 2.7894641759030301e-11, 
    2.7751925611768603e-11, 2.7663537894805873e-11, 2.7630091797903993e-11, 
    2.7649352688367295e-11, 2.7716531511457476e-11, 2.7824714780105006e-11, 
    2.7965418704840722e-11, 2.812921701017915e-11, 2.8306424212258863e-11, 
    2.8487786847100558e-11, 2.8665120642523343e-11, 2.88318606589118e-11, 
    2.8983476604402401e-11, 2.9117705757391189e-11, 2.9234600513479149e-11, 
    2.9336362913691225e-11, 2.9426998907169037e-11, 2.9511814075042178e-11, 
    2.9596801129214641e-11, 2.9687987485347763e-11, 2.9790793253784977e-11, 
    2.9909459346260668e-11, 3.004659137750446e-11, 3.0202862111309049e-11, 
    3.037685381527461e-11, 3.0565064174034618e-11, 3.0762037566784342e-11, 
    3.0960605463743639e-11, 3.1152199204593715e-11, 3.1327220012998369e-11, 
    3.1475440625727995e-11, 3.1586435620305392e-11, 3.1650031989687424e-11, 
    3.165678544599014e-11, 3.1598478278083388e-11, 3.146862670602669e-11, 
    3.1262978291749475e-11, 3.0979967415660409e-11, 3.062108433718833e-11, 
    3.019111258252266e-11, 2.9698187393961361e-11, 2.9153635213959237e-11, 
    2.8571581015485803e-11, 2.796832111674902e-11, 2.7361499272342673e-11, 
    2.6769131671411431e-11, 2.620856421741825e-11, 2.5695447930131264e-11, 
    2.5242824881892797e-11, 2.486039885246254e-11, 2.4554063524769848e-11, 
    2.4325716491627731e-11, 2.4173371678381153e-11, 2.4091531489476117e-11, 
    2.4071793240067878e-11, 2.4103582276056436e-11, 2.4174974447588839e-11, 
    2.4273500688870888e-11, 2.438688582819779e-11, 2.4503659322471714e-11, 
    2.4613632760807591e-11, 2.4708225652234418e-11, 2.4780662655446041e-11, 
    2.4826075753515273e-11, 2.4841538163565154e-11,
  // Sqw-total(7, 0-1999)
    0.023501003581474594, 0.023501998820253334, 0.023504851600812806, 
    0.023509169258947426, 0.023514317535977821, 0.023519449823961161, 
    0.023523546080683272, 0.023525459454596429, 0.023523968213539262, 
    0.023517830231255071, 0.023505837088644191, 0.023486864824410047, 
    0.023459918543293778, 0.02342416846370815, 0.0233789755441993, 
    0.023323905533137974, 0.023258731084162942, 0.023183422405366243, 
    0.023098127693311776, 0.023003145278155918, 0.02289888991914402, 
    0.022785856002740343, 0.022664580489799906, 0.022535608333757774, 
    0.022399462766152688, 0.022256622350074348, 0.022107506077570203, 
    0.021952467081490613, 0.021791794797188364, 0.021625724697821747, 
    0.021454454091061535, 0.021278161954385172, 0.021097030445019229, 
    0.020911265584071886, 0.020721114704319366, 0.020526878571646857, 
    0.020328916624224237, 0.020127644481076467, 0.019923523690706428, 
    0.019717044541020731, 0.019508703543931624, 0.019298977851418847, 
    0.019088299275487254, 0.018877030715541494, 0.018665447617500646, 
    0.018453726610196255, 0.018241942733886053, 0.018030075773204209, 
    0.01781802523604456, 0.017605632594819322, 0.017392708637322538, 
    0.017179063252515243, 0.016964534762321799, 0.016749016024839272, 
    0.016532474955392503, 0.016314967778027691, 0.01609664413871903, 
    0.015877744072602992, 0.015658587609520002, 0.015439558428938464, 
    0.015221083370408358, 0.015003609741395731, 0.014787582254782151, 
    0.014573421124992233, 0.014361502432757963, 0.014152141423366344, 
    0.013945579015523729, 0.013741971530138224, 0.013541383530562287, 
    0.013343783691796072, 0.013149043745995336, 0.012956940721897682, 
    0.012767162833884429, 0.012579319416743368, 0.012392955200689918, 
    0.012207568965087902, 0.012022636220519857, 0.011837635100256906, 
    0.01165207416768624, 0.011465520446888052, 0.011277625732421104, 
    0.011088149183405987, 0.010896974378006788, 0.010704119385846171, 
    0.010509738965484487, 0.010314118646566187, 0.010117661134117512, 
    0.0099208660980183178, 0.0097243049165707928, 0.0095285922806439046, 
    0.0093343567084526822, 0.0091422119690038744, 0.0089527311846800215, 
    0.0087664250176344716, 0.0085837248893339615, 0.0084049716916397461, 
    0.0082304099743585966, 0.0080601871851171975, 0.0078943572288408953, 
    0.0077328874279926491, 0.0075756679067997892, 0.0074225224822130446, 
    0.0072732202957656233, 0.0071274876272421185, 0.006985019551012021, 
    0.0068454912880498917, 0.006708569237914597, 0.0065739217256683769, 
    0.0064412294661443034, 0.0063101956466804074, 0.0061805553884073019, 
    0.0060520842031556634, 0.0059246049571040696, 0.0057979928160558176, 
    0.0056721777003506668, 0.0055471439224881128, 0.0054229269023570552, 
    0.0052996071231802859, 0.0051773017658596626, 0.00505615469786756, 
    0.004936325657758615, 0.0048179795419167675, 0.0047012766562134142, 
    0.0045863646488933365, 0.0044733726147741411, 0.0043624075886045111, 
    0.0042535533664590603, 0.0041468713465935177, 0.0040424028965044476, 
    0.0039401726509175755, 0.0038401921322802871, 0.0037424631537305649, 
    0.0036469805958477702, 0.0035537343167973659, 0.0034627101321697937, 
    0.0033738899593757994, 0.0032872513413314459, 0.0032027666332101147, 
    0.0031204021513382228, 0.003040117550383727, 0.0029618656257115786, 
    0.0028855926476330481, 0.0028112392393886479, 0.0027387417253566244, 
    0.0026680338108057539, 0.0025990484156577691, 0.0025317194738285116, 
    0.002465983524581712, 0.0024017809579430951, 0.0023390568259155317, 
    0.0022777611876984129, 0.0022178490132361826, 0.002159279718868673, 
    0.0021020164464973109, 0.0020460252198702135, 0.0019912741164012388, 
    0.0019377325803259101, 0.0018853709748540811, 0.0018341604310225931, 
    0.0017840730043917773, 0.0017350821036918656, 0.00168716311428033, 
    0.0016402941093603919, 0.0015944565273366459, 0.0015496356962778053, 
    0.001505821105597822, 0.0014630063577646246, 0.0014211887742302787, 
    0.001380368673860772, 0.0013405483827700702, 0.0013017310662234117, 
    0.0012639194922901501, 0.0012271148413319508, 0.0011913156655205678, 
    0.0011565170806852002, 0.0011227102427075004, 0.0010898821270750917, 
    0.001058015597849493, 0.0010270897253811672, 0.00099708029363629823, 
    0.00096796042948526573, 0.00093970128762154912, 0.00091227273432409751, 
    0.00088564398833633159, 0.00085978419440591058, 0.00083466292122383171, 
    0.00081025058789696417, 0.00078651882998104076, 0.00076344081703000864, 
    0.00074099152937587677, 0.00071914799423849444, 0.00069788947267412384, 
    0.00067719758177211024, 0.00065705633294328811, 0.00063745206832029869, 
    0.00061837328338509292, 0.0005998103340897809, 0.00058175503926961815, 
    0.00056420020192311337, 0.00054713908379134776, 0.0005305648748069263, 
    0.00051447020127380724, 0.00049884671375940569, 0.00048368478810837095, 
    0.00046897336183990263, 0.00045469991499413014, 0.00044085059090405351, 
    0.00042741043993797562, 0.00041436375923213642, 0.000401694494664696, 
    0.00038938666821587313, 0.0003774247944117823, 0.00036579425339600954, 
    0.00035448159467438528, 0.00034347475389468618, 0.00033276317420556222, 
    0.00032233783280894796, 0.00031219118136595293, 0.00030231701517584639, 
    0.00029271029000163318, 0.00028336690684167479, 0.00027428348395938098, 
    0.00026545713250726528, 0.0002568852477977484, 0.00024856532349621318, 
    0.00024049479156609981, 0.00023267088736606998, 0.00022509053732521812, 
    0.00021775026622163174, 0.00021064612205979062, 0.00020377361840556184, 
    0.00019712769615647062, 0.00019070270842706761, 0.00018449243295460177, 
    0.00017849011583353868, 0.00017268854841614312, 0.00016708017610900087, 
    0.00016165723404646076, 0.00015641190087814144, 0.00015133645885697769, 
    0.00014642344665361084, 0.00014166579125861006, 0.00013705690710337276, 
    0.00013259075398335863, 0.00012826185008039552, 0.00012406524173033301, 
    0.00011999643682971859, 0.00011605131318512183, 0.00011222601604915127, 
    0.00010851686012779873, 0.00010492025031152175, 0.00010143263239512536, 
    9.8050480495751407e-05, 9.4770322367100356e-05, 9.1588798089134335e-05, 
    8.8502742475809012e-05, 8.5509277701217745e-05, 8.2605900641360589e-05, 
    7.9790549553420206e-05, 7.7061636966928028e-05, 7.4418039742084208e-05, 
    7.1859042612722207e-05, 6.9384237449901265e-05, 6.6993386167884196e-05, 
    6.468625989859193e-05, 6.2462470189223764e-05, 6.0321309161223668e-05, 
    5.8261614714249057e-05, 5.6281674141751698e-05, 5.4379175358197597e-05, 
    5.255120989147719e-05, 5.0794326515080593e-05, 4.9104629505486471e-05, 
    4.7477911538435912e-05, 4.5909808548316499e-05, 4.4395962650549035e-05, 
    4.2932179459238385e-05, 4.1514567654957351e-05, 4.0139651179632138e-05, 
    3.880444760031295e-05, 3.750650961065755e-05, 3.6243929975509326e-05, 
    3.5015313170256203e-05, 3.3819719304241871e-05, 3.2656587510115387e-05, 
    3.1525646782035435e-05, 3.0426822280632053e-05, 2.9360144485210797e-05, 
    2.8325667399465402e-05, 2.7323400475377357e-05, 2.6353257187132373e-05, 
    2.5415021438022825e-05, 2.4508331369895882e-05, 2.363267879114148e-05, 
    2.2787421427618077e-05, 2.1971804575983969e-05, 2.1184988500945888e-05, 
    2.0426078036008574e-05, 1.9694151259189905e-05, 1.898828474418671e-05, 
    1.8307573645065375e-05, 1.7651145674486286e-05, 1.7018168801697367e-05, 
    1.6407853164273909e-05, 1.581944820727868e-05, 1.5252236407693479e-05, 
    1.4705525098658235e-05, 1.4178637886398161e-05, 1.3670906974391652e-05, 
    1.3181667412298924e-05, 1.2710253914599084e-05, 1.2256000496920473e-05, 
    1.1818242802397084e-05, 1.1396322679416621e-05, 1.0989594353323882e-05, 
    1.0597431425242597e-05, 1.0219233927838985e-05, 9.8544347567534582e-06, 
    9.5025049481373022e-06, 9.1629574557706421e-06, 8.8353492606026143e-06, 
    8.5192817962314868e-06, 8.2143997777764853e-06, 7.9203885772334092e-06, 
    7.6369703026956003e-06, 7.3638987306234156e-06, 7.1009532288751981e-06, 
    6.8479318134691768e-06, 6.6046435137165941e-06, 6.3709002814495745e-06, 
    6.1465087595267321e-06, 5.9312623075004102e-06, 5.7249337454901491e-06, 
    5.5272693034060758e-06, 5.3379842365997421e-06, 5.1567604883344697e-06, 
    4.9832466483895054e-06, 4.8170602915880171e-06, 4.6577925984667907e-06, 
    4.5050149854107725e-06, 4.3582873209615933e-06, 4.217167194009587e-06, 
    4.0812196344906411e-06, 3.9500266712413063e-06, 3.8231961402574947e-06, 
    3.700369225518071e-06, 3.581226314855871e-06, 3.4654908791528854e-06, 
    3.35293122466485e-06, 3.2433601187836813e-06, 3.1366324376871944e-06, 
    3.0326411207780392e-06, 2.9313118283576553e-06, 2.8325967760603303e-06, 
    2.7364682516012169e-06, 2.6429123034523571e-06, 2.5519230264604454e-06, 
    2.463497765261743e-06, 2.3776334241152257e-06, 2.2943239304139234e-06, 
    2.2135587658444475e-06, 2.1353223725249762e-06, 2.0595941731602329e-06, 
    1.9863489219885995e-06, 1.9155571251260145e-06, 1.8471853286091637e-06, 
    1.7811961557491014e-06, 1.7175480681824115e-06, 1.6561949099918709e-06, 
    1.5970853597348742e-06, 1.5401624507674854e-06, 1.485363323875588e-06, 
    1.4326193486166048e-06, 1.381856698816247e-06, 1.3329974015843159e-06, 
    1.285960810570317e-06, 1.2406653918955654e-06, 1.1970306653195717e-06, 
    1.1549791182399691e-06, 1.1144379097064192e-06, 1.0753402037309858e-06, 
    1.0376260135137675e-06, 1.001242493543095e-06, 9.6614367923998889e-07, 
    9.322897346337692e-07, 8.9964582165443133e-07, 8.6818074202929053e-07, 
    8.378655214389684e-07, 8.0867210164309812e-07, 7.8057228154999355e-07, 
    7.5353700453389974e-07, 7.2753603382722135e-07, 7.0253799692373604e-07, 
    6.7851072401300893e-07, 6.554217615026922e-07, 6.3323891823236228e-07, 
    6.1193070183728519e-07, 5.9146652758557081e-07, 5.7181662716975116e-07, 
    5.5295164449413898e-07, 5.3484196837918778e-07, 5.1745690907941208e-07, 
    5.0076386519303916e-07, 4.8472764419283785e-07, 4.6931008863646772e-07, 
    4.5447012368195818e-07, 4.4016428426116632e-07, 4.2634771227805308e-07, 
    4.1297554532163855e-07, 4.0000456056720381e-07, 3.8739489840578581e-07, 
    3.7511167691140657e-07, 3.6312632040439268e-07, 3.514174616962235e-07, 
    3.3997133055321522e-07, 3.2878160295126136e-07, 3.1784874648053916e-07, 
    3.0717894937816583e-07, 2.9678275669239902e-07, 2.8667355479515825e-07, 
    2.7686604335144743e-07, 2.6737481600612637e-07, 2.582131407831802e-07, 
    2.4939199574607384e-07, 2.4091937957351874e-07, 2.3279988643559337e-07, 
    2.2503451234111997e-07, 2.1762064862055514e-07, 2.1055221581869049e-07, 
    2.0381989752824273e-07, 1.974114441701895e-07, 1.9131202957475787e-07, 
    1.855046539007093e-07, 1.7997059386391381e-07, 1.7468990282031951e-07, 
    1.6964196005947647e-07, 1.6480606050830525e-07, 1.6016202597244622e-07, 
    1.5569080838960957e-07, 1.5137504775377597e-07, 1.4719954352429789e-07, 
    1.4315160065115778e-07, 1.3922121906391859e-07, 1.3540110893621655e-07, 
    1.3168653029714466e-07, 1.2807497357103231e-07, 1.2456571362414557e-07, 
    1.2115928274181753e-07, 1.1785691483785533e-07, 1.1466001432157957e-07, 
    1.1156969735244866e-07, 1.0858644275050761e-07, 1.0570987500051013e-07, 
    1.0293868567031641e-07, 1.0027068304579926e-07, 9.7702945869230052e-08, 
    9.5232046155614719e-08, 9.2854300268484002e-08, 9.0566006272832251e-08, 
    8.8363630154912179e-08, 8.6243912126631769e-08, 8.4203877110749089e-08, 
    8.2240748101296314e-08, 8.0351776538893252e-08, 7.8534017272271213e-08, 
    7.6784086051696779e-08, 7.509794207729978e-08, 7.3470737105873132e-08, 
    7.1896764536543613e-08, 7.0369528893608307e-08, 6.8881938797563994e-08, 
    6.7426608528179233e-08, 6.5996236597480656e-08, 6.4584017928345887e-08, 
    6.3184040544463876e-08, 6.179161988720049e-08, 6.0403532770233806e-08, 
    5.9018127778505947e-08, 5.7635306216864943e-08, 5.6256385282388805e-08, 
    5.4883869141707935e-08, 5.3521162854006078e-08, 5.2172266392764861e-08, 
    5.0841482629515753e-08, 4.9533164287127675e-08, 4.8251513798011916e-08, 
    4.7000438071554906e-08, 4.5783450743443112e-08, 4.4603608165320993e-08, 
    4.3463463846663941e-08, 4.2365028090516202e-08, 4.1309725048073605e-08, 
    4.0298345702200546e-08, 3.9331001866063197e-08, 3.8407090471896458e-08, 
    3.7525279567424426e-08, 3.6683526136964368e-08, 3.5879132681734185e-08, 
    3.5108844179556675e-08, 3.4368981733619662e-08, 3.36556040985204e-08, 
    3.2964684975791348e-08, 3.2292292103449142e-08, 3.1634754708219341e-08, 
    3.0988807496973985e-08, 3.0351702678067083e-08, 2.9721284707045933e-08, 
    2.9096026206681832e-08, 2.8475026325844221e-08, 2.7857975483550535e-08, 
    2.7245091961006285e-08, 2.6637037133384178e-08, 2.6034816470795837e-08, 
    2.5439673787928543e-08, 2.4852985618102331e-08, 2.4276162125364364e-08, 
    2.3710559555227137e-08, 2.3157408025534723e-08, 2.2617756416445356e-08, 
    2.2092434626462417e-08, 2.1582031573302568e-08, 2.1086886367665952e-08, 
    2.0607089321924367e-08, 2.0142489812630916e-08, 1.9692708653053749e-08, 
    1.9257154143863439e-08, 1.8835042225599867e-08, 1.8425422564678498e-08, 
    1.8027212858196436e-08, 1.7639243636300197e-08, 1.7260314539975541e-08, 
    1.6889261352986668e-08, 1.6525030507349356e-08, 1.6166755687112756e-08, 
    1.5813829012780285e-08, 1.5465958684182837e-08, 1.5123205004681728e-08, 
    1.4785988626581435e-08, 1.4455067378973882e-08, 1.4131481861166359e-08, 
    1.3816473480528494e-08, 1.3511382274572212e-08, 1.3217534080583738e-08, 
    1.2936128160437993e-08, 1.2668135912698933e-08, 1.2414220032268296e-08, 
    1.2174680692780878e-08, 1.1949432348927047e-08, 1.1738011252401115e-08, 
    1.1539610983363181e-08, 1.1353140792887282e-08, 1.1177300331984533e-08, 
    1.1010663589913064e-08, 1.0851765305527441e-08, 1.0699183703208539e-08, 
    1.0551614786150064e-08, 1.0407934393683361e-08, 1.0267245627603928e-08, 
    1.0128910033647585e-08, 9.9925619238412245e-09, 9.8581056910362642e-09, 
    9.7256968209719847e-09, 9.5957076878028147e-09, 9.468680087672601e-09, 
    9.3452670149764716e-09, 9.2261670968141814e-09, 9.1120555813486442e-09, 
    9.0035164184564033e-09, 8.9009800217260576e-09, 8.8046713784079336e-09, 
    8.7145724360548689e-09, 8.6304020533203395e-09, 8.5516153858030372e-09, 
    8.4774233694063525e-09, 8.4068312564699276e-09, 8.3386937874262519e-09, 
    8.2717831342839579e-09, 8.2048647865930976e-09, 8.1367757129085985e-09, 
    8.0664990869681362e-09, 7.9932298818827359e-09, 7.9164265380244305e-09, 
    7.8358448002026758e-09, 7.7515514610796581e-09, 7.6639170533925035e-09, 
    7.5735884480246307e-09, 7.4814435272480325e-09, 7.3885316316778101e-09, 
    7.2960041431154784e-09, 7.2050403277803582e-09, 7.1167734106799794e-09, 
    7.0322218011387035e-09, 6.9522295320548943e-09, 6.8774193381997109e-09, 
    6.8081605399884729e-09, 6.7445530736556483e-09, 6.6864277359158523e-09, 
    6.6333619508021925e-09, 6.5847093656068963e-09, 6.5396411277245918e-09, 
    6.4971959852708678e-09, 6.4563362821882228e-09, 6.4160065441228857e-09, 
    6.3751915611219668e-09, 6.3329708057661273e-09, 6.2885665041289217e-09, 
    6.2413828128988947e-09, 6.1910342716364979e-09, 6.1373620079562932e-09, 
    6.0804370496564331e-09, 6.0205505573453684e-09, 5.9581916919658828e-09, 
    5.8940143514845553e-09, 5.8287948460627241e-09, 5.7633829624333647e-09, 
    5.6986494748516483e-09, 5.63543322974243e-09, 5.5744911962298566e-09, 
    5.5164544935233236e-09, 5.461793226269203e-09, 5.410792192690987e-09, 
    5.3635389442263177e-09, 5.319924644023428e-09, 5.2796574455486317e-09, 
    5.2422870830096999e-09, 5.2072387392294019e-09, 5.1738535153204621e-09, 
    5.141432636017526e-09, 5.1092821707443706e-09, 5.0767554041938358e-09, 
    5.043290043428418e-09, 5.0084382489472092e-09, 4.9718878090713891e-09, 
    4.9334737328749045e-09, 4.893179983296611e-09, 4.8511319212046904e-09, 
    4.8075803832319168e-09, 4.7628789462400725e-09, 4.7174560182503703e-09, 
    4.6717838186384134e-09, 4.6263461180865066e-09, 4.5816068023728781e-09, 
    4.5379809518853063e-09, 4.4958101248421347e-09, 4.4553430522916305e-09, 
    4.416722781819581e-09, 4.3799807765383544e-09, 4.3450382262816928e-09, 
    4.3117142355456639e-09, 4.2797403372095809e-09, 4.2487802127363587e-09, 
    4.218453366290609e-09, 4.1883610403517373e-09, 4.158112774623861e-09, 
    4.1273517216542128e-09, 4.0957771778874009e-09, 4.0631627647130553e-09, 
    4.0293692908831241e-09, 3.9943514689561172e-09, 3.958158344945779e-09, 
    3.9209275670623166e-09, 3.8828742194480481e-09, 3.8442751397248464e-09, 
    3.8054500657585595e-09, 3.7667409269011858e-09, 3.7284908190200492e-09, 
    3.6910239129265052e-09, 3.6546275995738815e-09, 3.6195377348028924e-09, 
    3.5859277671513348e-09, 3.55390205783498e-09, 3.5234936353471619e-09, 
    3.4946661737706772e-09, 3.4673199442617992e-09, 3.4413011417553172e-09, 
    3.4164140089356759e-09, 3.3924348632888186e-09, 3.3691272837832038e-09, 
    3.3462574081878072e-09, 3.3236085374507005e-09, 3.300994064362872e-09, 
    3.2782680232834169e-09, 3.2553325020764481e-09, 3.2321415682658809e-09, 
    3.2087013784515169e-09, 3.1850665680509067e-09, 3.1613331470194363e-09, 
    3.1376285199585678e-09, 3.1140992911837362e-09, 3.0908978905799649e-09, 
    3.0681689385393e-09, 3.0460364807359575e-09, 3.0245929652933171e-09, 
    3.0038908998128226e-09, 2.9839376985428068e-09, 2.9646941737714297e-09, 
    2.9460766303178643e-09, 2.9279624476335523e-09, 2.910198533322208e-09, 
    2.8926120346675301e-09, 2.8750223177645757e-09, 2.8572533514975767e-09, 
    2.8391454490292873e-09, 2.8205655878901844e-09, 2.8014155070604856e-09, 
    2.7816371782119844e-09, 2.7612153023844853e-09, 2.740176902383713e-09, 
    2.7185881375376932e-09, 2.6965488323241076e-09, 2.6741851533919289e-09, 
    2.651641149242131e-09, 2.6290696871679056e-09, 2.6066234987846592e-09, 
    2.5844467676060487e-09, 2.5626678185670655e-09, 2.5413931666259873e-09, 
    2.5207032340241021e-09, 2.5006497906553869e-09, 2.4812552317838595e-09, 
    2.4625135437694919e-09, 2.4443929013456295e-09, 2.426839578924669e-09, 
    2.4097830084734066e-09, 2.3931415615764997e-09, 2.3768287937188057e-09, 
    2.3607596905368837e-09, 2.344856637049245e-09, 2.3290546894218702e-09, 
    2.313305908077037e-09, 2.2975824241964219e-09, 2.281878140882564e-09, 
    2.2662088549259948e-09, 2.2506108987592231e-09, 2.235138265126599e-09, 
    2.2198584989949885e-09, 2.2048475233369831e-09, 2.190183837374356e-09, 
    2.1759424263178015e-09, 2.1621888862868592e-09, 2.1489741363191701e-09, 
    2.1363302128867504e-09, 2.124267370100317e-09, 2.1127728190710217e-09, 
    2.1018110790912437e-09, 2.0913260051615032e-09, 2.0812442063254537e-09, 
    2.0714796305813055e-09, 2.0619388446595103e-09, 2.0525266647022941e-09, 
    2.0431515998131254e-09, 2.0337308112084702e-09, 2.0241941708463517e-09, 
    2.0144872875910055e-09, 2.0045733151308461e-09, 1.9944336078053693e-09, 
    1.9840672482907021e-09, 1.9734896819776522e-09, 1.9627305679136546e-09, 
    1.9518311563356342e-09, 1.9408412961319269e-09, 1.929816336346271e-09, 
    1.918813977411066e-09, 1.9078912610819042e-09, 1.8971016988748405e-09, 
    1.8864926949606095e-09, 1.8761032355385912e-09, 1.8659620076614943e-09, 
    1.8560859524753069e-09, 1.8464794069361334e-09, 1.8371338332730674e-09, 
    1.8280283034992561e-09, 1.8191306727001752e-09, 1.8103995062502575e-09, 
    1.8017866329722712e-09, 1.7932402425699628e-09, 1.7847082920983938e-09, 
    1.776142056935796e-09, 1.7674994854931113e-09, 1.7587482002272821e-09, 
    1.749867809392695e-09, 1.7408514200834006e-09, 1.7317061413019546e-09, 
    1.7224526052133019e-09, 1.7131234515928006e-09, 1.7037609579554877e-09, 
    1.6944139474152818e-09, 1.6851342638905647e-09, 1.6759730184825708e-09, 
    1.6669770026434534e-09, 1.6581854411056371e-09, 1.6496274100452411e-09, 
    1.6413200353412758e-09, 1.6332676484323345e-09, 1.6254618658503851e-09, 
    1.6178826259980412e-09, 1.610499960274064e-09, 1.6032764408566797e-09, 
    1.59616997788386e-09, 1.5891368095233808e-09, 1.5821343909171203e-09, 
    1.5751240237963468e-09, 1.5680729867711671e-09, 1.5609561189724846e-09, 
    1.5537567068159118e-09, 1.5464667536441913e-09, 1.5390865822861136e-09, 
    1.5316239553278672e-09, 1.5240927436093603e-09, 1.5165113588686876e-09, 
    1.5089010282806514e-09, 1.5012841043179943e-09, 1.493682467162943e-09, 
    1.4861161710988331e-09, 1.4786023305906339e-09, 1.4711543613343327e-09, 
    1.4637814917414202e-09, 1.4564886325598652e-09, 1.4492764896147665e-09, 
    1.4421419643547707e-09, 1.435078720014404e-09, 1.4280779534400279e-09, 
    1.4211292431705084e-09, 1.414221501808015e-09, 1.4073439036197746e-09, 
    1.4004868189979541e-09, 1.3936426224535331e-09, 1.3868063973986936e-09, 
    1.3799764257119752e-09, 1.3731544814764258e-09, 1.3663458548936851e-09, 
    1.3595591493223161e-09, 1.3528057882628558e-09, 1.3460993406923195e-09, 
    1.339454618327256e-09, 1.3328866808806138e-09, 1.3264097334615083e-09, 
    1.3200360520622631e-09, 1.3137749526160725e-09, 1.307631917881041e-09, 
    1.3016078825305025e-09, 1.2956988024626544e-09, 1.2898954623937903e-09, 
    1.2841836362249463e-09, 1.2785445127122936e-09, 1.2729554681546273e-09, 
    1.2673910803958491e-09, 1.2618243979297593e-09, 1.2562283309085807e-09, 
    1.2505771586157598e-09, 1.2448479829614927e-09, 1.23902211054783e-09, 
    1.233086181639411e-09, 1.2270330662144442e-09, 1.2208623506634226e-09, 
    1.214580473714444e-09, 1.2082004124705864e-09, 1.2017410042347763e-09, 
    1.1952258749028046e-09, 1.1886821133241839e-09, 1.1821387230473188e-09, 
    1.1756250124671422e-09, 1.1691689689220544e-09, 1.1627958073040344e-09, 
    1.1565267019427595e-09, 1.1503778732439341e-09, 1.1443599796286173e-09, 
    1.1384779439788398e-09, 1.1327310956744672e-09, 1.1271136905349449e-09, 
    1.1216156529789983e-09, 1.1162235370519051e-09, 1.110921548190207e-09, 
    1.1056926058926975e-09, 1.1005192876347932e-09, 1.0953846867140091e-09, 
    1.0902730648358585e-09, 1.0851703557462107e-09, 1.0800644604234823e-09, 
    1.0749454333545971e-09, 1.0698055187391953e-09, 1.0646391506638057e-09, 
    1.0594428663955813e-09, 1.0542152375640058e-09, 1.0489567546924383e-09, 
    1.0436697355290376e-09, 1.0383581556726846e-09, 1.0330274923013758e-09, 
    1.0276844671990235e-09, 1.0223367636415469e-09, 1.0169926340946732e-09, 
    1.011660492169487e-09, 1.0063484280742772e-09, 1.0010637443944603e-09, 
    9.9581248490556937e-10, 9.9059905801707232e-10, 9.8542589883749393e-10, 
    9.8029331134847066e-10, 9.7519941854883032e-10, 9.7014030547528613e-10, 
    9.651103084372748e-10, 9.6010249104177603e-10, 9.5510923845190413e-10, 
    9.5012298828109357e-10, 9.4513697940302592e-10, 9.4014603884986517e-10, 
    9.3514726286949142e-10, 9.3014059643369644e-10, 9.2512918008550882e-10, 
    9.2011948834666244e-10, 9.1512117730486568e-10, 9.1014668316355577e-10, 
    9.0521055843419563e-10, 9.0032865313718889e-10, 8.9551713880863906e-10, 
    8.9079154416021195e-10, 8.8616580282257885e-10, 8.8165147228609166e-10, 
    8.7725710518094716e-10, 8.7298789784514989e-10, 8.6884553819987253e-10, 
    8.648283326124074e-10, 8.6093149442683227e-10, 8.5714763047286635e-10, 
    8.5346727979971262e-10, 8.498795478885084e-10, 8.4637269470215589e-10, 
    8.4293472059358971e-10, 8.3955383635686001e-10, 8.3621888991261752e-10, 
    8.3291964452497946e-10, 8.2964699012980538e-10, 8.2639302073046706e-10, 
    8.2315104134266517e-10, 8.1991543822666554e-10, 8.1668149883597198e-10, 
    8.1344513512815453e-10, 8.1020258375836622e-10, 8.0695006083406187e-10, 
    8.0368347143057321e-10, 8.003981518282083e-10, 7.9708876024629669e-10, 
    7.9374926389811354e-10, 7.9037314017404352e-10, 7.8695371099496669e-10, 
    7.8348467069595646e-10, 7.7996069065914666e-10, 7.763781272835063e-10, 
    7.727356719468982e-10, 7.6903495826015261e-10, 7.6528094472651035e-10, 
    7.614821359665731e-10, 7.5765046293332085e-10, 7.5380094235201618e-10, 
    7.4995102165735621e-10, 7.4611973515630804e-10, 7.423266690630119e-10, 
    7.3859089647121546e-10, 7.3492989151692547e-10, 7.3135860578306245e-10, 
    7.2788868616832488e-10, 7.2452798728476777e-10, 7.2128031642981299e-10, 
    7.1814549555141352e-10, 7.1511962424157256e-10, 7.1219558010615213e-10, 
    7.0936360583889168e-10, 7.066119994998767e-10, 7.0392775154651194e-10, 
    7.0129717392554489e-10, 6.987064060233993e-10, 6.9614187363763954e-10, 
    6.9359061998305474e-10, 6.9104061904576423e-10, 6.8848103688669935e-10, 
    6.8590250638456238e-10, 6.8329736808517198e-10, 6.8065995405122488e-10, 
    6.7798679748821971e-10, 6.7527682900886734e-10, 6.7253143525393859e-10, 
    6.6975442502793467e-10, 6.669517990607172e-10, 6.6413140262518547e-10, 
    6.6130239961512291e-10, 6.5847467532133211e-10, 6.5565815579936536e-10, 
    6.5286217188478304e-10, 6.5009485161268298e-10, 6.4736267418516366e-10, 
    6.4467014724569241e-10, 6.4201969281241334e-10, 6.3941166789329057e-10, 
    6.368445807224009e-10, 6.3431539733677385e-10, 6.3181997023126033e-10, 
    6.2935348037370665e-10, 6.2691091681107752e-10, 6.244875139234911e-10, 
    6.2207916032161647e-10, 6.19682709684198e-10, 6.1729624634352852e-10, 
    6.1491921669946263e-10, 6.1255250590456968e-10, 6.1019837551215738e-10, 
    6.0786034990771447e-10, 6.0554296508852356e-10, 6.032514897012119e-10, 
    6.0099154384633613e-10, 5.9876870513268619e-10, 5.9658808967377462e-10, 
    5.9445395216032524e-10, 5.9236930827513892e-10, 5.9033565455850448e-10, 
    5.8835274368611331e-10, 5.8641850588120407e-10, 5.8452905394776564e-10, 
    5.8267884482453465e-10, 5.8086092824500088e-10, 5.7906732665030103e-10, 
    5.7728947336659045e-10, 5.7551873026539896e-10, 5.7374690112204884e-10, 
    5.7196676032610653e-10, 5.7017249860981832e-10, 5.6836012274626652e-10, 
    5.6652769648311744e-10, 5.6467548112372071e-10, 5.628058959749325e-10, 
    5.6092334748295939e-10, 5.5903388591886378e-10, 5.5714477175357518e-10, 
    5.5526391899181106e-10, 5.533993208122092e-10, 5.5155845052739591e-10, 
    5.4974772669610416e-10, 5.4797205043996078e-10, 5.4623447871615736e-10, 
    5.4453602296488727e-10, 5.4287561751920947e-10, 5.4125020081741061e-10, 
    5.3965494394292366e-10, 5.3808353578282026e-10, 5.3652854414377867e-10, 
    5.3498177060755172e-10, 5.334346078854827e-10, 5.318783365954381e-10, 
    5.3030439602279823e-10, 5.287045833278577e-10, 5.2707123886769196e-10, 
    5.2539737970488737e-10, 5.2367685861495634e-10, 5.2190449791261822e-10, 
    5.2007626270675046e-10, 5.1818942030713025e-10, 5.1624271044232505e-10, 
    5.1423646863611324e-10, 5.1217271312828383e-10, 5.100551306927584e-10, 
    5.0788898495211681e-10, 5.0568088849929614e-10, 5.0343850787689346e-10, 
    5.0117015294553845e-10, 4.9888435157703357e-10, 4.9658940801554925e-10, 
    4.9429302202191031e-10, 4.9200197990328055e-10, 4.8972199615875279e-10, 
    4.8745766865069994e-10, 4.8521259478199262e-10, 4.8298958473929037e-10, 
    4.8079096258559577e-10, 4.786188877323629e-10, 4.7647565965603679e-10, 
    4.7436392688315733e-10, 4.7228680721046613e-10, 4.7024784940350263e-10, 
    4.6825088096825348e-10, 4.6629971644363087e-10, 4.6439779933707382e-10, 
    4.625477912929656e-10, 4.6075118655672904e-10, 4.5900796549839667e-10, 
    4.573163620226545e-10, 4.5567274043664532e-10, 4.5407161722107106e-10, 
    4.5250580187038567e-10, 4.5096668014031924e-10, 4.4944455148794986e-10, 
    4.4792908043539423e-10, 4.464097506120561e-10, 4.4487635752435791e-10, 
    4.4331946595832392e-10, 4.4173085289819452e-10, 4.4010388206874064e-10, 
    4.3843381521347246e-10, 4.3671803129802782e-10, 4.3495614794291501e-10, 
    4.3315001290310031e-10, 4.3130359458873116e-10, 4.2942272975403812e-10, 
    4.2751478259835339e-10, 4.2558820361181179e-10, 4.236520470139831e-10, 
    4.2171547096033953e-10, 4.1978728437831484e-10, 4.1787555589624079e-10, 
    4.1598734960437183e-10, 4.1412857852881588e-10, 4.1230399481911496e-10, 
    4.105172902073667e-10, 4.0877128889104815e-10, 4.0706815860697382e-10, 
    4.054096407687098e-10, 4.0379720798409738e-10, 4.0223217445113122e-10, 
    4.007156762828664e-10, 3.9924859777232052e-10, 3.9783140452910734e-10, 
    3.9646395599057151e-10, 3.9514530531902355e-10, 3.9387355539997313e-10, 
    3.9264577804988185e-10, 3.914580369149759e-10, 3.9030549830793922e-10, 
    3.8918265683166163e-10, 3.8808360055903759e-10, 3.8700234531655691e-10, 
    3.8593314541092056e-10, 3.8487078763103469e-10, 3.8381080116024493e-10, 
    3.8274959794008905e-10, 3.8168449540835687e-10, 3.806136485769964e-10, 
    3.7953588787738673e-10, 3.7845050561472299e-10, 3.7735697660735622e-10, 
    3.7625470352174314e-10, 3.7514275598173438e-10, 3.7401968614794255e-10, 
    3.7288340349376597e-10, 3.7173114781602152e-10, 3.705595466561742e-10, 
    3.6936478227504679e-10, 3.6814280889955943e-10, 3.6688965049657576e-10, 
    3.6560172296120254e-10, 3.6427617035128324e-10, 3.6291116385740602e-10, 
    3.6150617347436808e-10, 3.6006215106314444e-10, 3.5858164744627008e-10, 
    3.5706880931953327e-10, 3.55529298833183e-10, 3.5397009576838692e-10, 
    3.5239923056329932e-10, 3.5082542096832501e-10, 3.4925768376984255e-10, 
    3.4770488813091604e-10, 3.4617533299520468e-10, 3.446763276548517e-10, 
    3.43213845730594e-10, 3.4179222888511788e-10, 3.404140080880252e-10, 
    3.3907980598440267e-10, 3.3778837846060121e-10, 3.3653672622592602e-10, 
    3.3532033601481095e-10, 3.3413348132631267e-10, 3.3296960424622354e-10, 
    3.318217091963697e-10, 3.3068280560218684e-10, 3.2954629132754576e-10, 
    3.2840634818125331e-10, 3.2725823807136681e-10, 3.2609854291100078e-10, 
    3.2492529642500716e-10, 3.2373801356515887e-10, 3.2253759556015321e-10, 
    3.2132614867626889e-10, 3.201066721652153e-10, 3.1888270763549545e-10, 
    3.1765791967918669e-10, 3.1643570429670813e-10, 3.1521880411794079e-10, 
    3.1400904472339491e-10, 3.1280715812123103e-10, 3.1161277697302953e-10, 
    3.1042454948028268e-10, 3.0924042239866839e-10, 3.0805800708717885e-10, 
    3.068750342385245e-10, 3.0568979113381579e-10, 3.0450154235215189e-10, 
    3.0331080947074125e-10, 3.0211954569940548e-10, 3.009311010767789e-10, 
    2.9975004428155747e-10, 2.9858180129367023e-10, 2.9743219037491926e-10, 
    2.9630686850011305e-10, 2.9521079199305587e-10, 2.9414768743804924e-10, 
    2.9311966248549943e-10, 2.9212692819582947e-10, 2.9116771815689287e-10, 
    2.9023835553092059e-10, 2.8933351712249268e-10, 2.8844661243972974e-10, 
    2.8757030358373008e-10, 2.8669704571111587e-10, 2.8581968189265254e-10, 
    2.8493197483048828e-10, 2.8402908401735344e-10, 2.8310790598397693e-10, 
    2.8216730028874087e-10, 2.8120813769509911e-10, 2.8023321780449189e-10, 
    2.7924702378617938e-10, 2.7825537855294133e-10, 2.7726500311306531e-10, 
    2.7628305567702992e-10, 2.7531664661142454e-10, 2.743724262869853e-10, 
    2.7345622131058193e-10, 2.7257279686090808e-10, 2.7172568098136955e-10, 
    2.7091712269960776e-10, 2.7014808315537017e-10, 2.6941830013247319e-10, 
    2.687263339890418e-10, 2.6806962037891918e-10, 2.6744446362171811e-10, 
    2.6684601123971096e-10, 2.6626817974506171e-10, 2.6570360437933827e-10, 
    2.6514358000380183e-10, 2.645781184953935e-10, 2.639960645702832e-10, 
    2.6338538315058853e-10, 2.6273354791932687e-10, 2.6202808731685517e-10, 
    2.6125720478715427e-10, 2.6041047673234154e-10, 2.594795304347518e-10, 
    2.5845869575293493e-10, 2.5734550811796481e-10, 2.5614110810812621e-10, 
    2.5485040506120599e-10, 2.5348208805307191e-10, 2.520484054565184e-10, 
    2.5056478559898963e-10, 2.4904926891642875e-10, 2.4752184680453973e-10, 
    2.4600367391823249e-10, 2.4451626977483371e-10, 2.430806755017186e-10, 
    2.4171667421853078e-10, 2.4044205807270926e-10, 2.3927201946154807e-10, 
    2.3821864186854731e-10, 2.3729057304501109e-10, 2.3649280811962174e-10, 
    2.358266584104593e-10, 2.3528982209281327e-10, 2.34876588424318e-10, 
    2.3457809255127074e-10, 2.3438266637070848e-10, 2.3427617820952846e-10, 
    2.342424247152909e-10, 2.3426351468428172e-10, 2.3432028866534095e-10, 
    2.343927490753998e-10, 2.3446056228103806e-10, 2.3450358344362836e-10, 
    2.3450247683810883e-10, 2.3443935335492511e-10, 2.3429847805564188e-10, 
    2.3406692631943182e-10, 2.3373523607164912e-10, 2.332979215421229e-10, 
    2.3275386838188316e-10, 2.3210650252087286e-10, 2.3136376944248407e-10, 
    2.3053783224320997e-10, 2.2964456673144033e-10, 2.2870281167223246e-10, 
    2.2773346352820739e-10, 2.26758412182835e-10, 2.2579944488991872e-10, 
    2.2487711000094252e-10, 2.2400967788114967e-10, 2.2321220568183262e-10, 
    2.2249580675443566e-10, 2.2186711028295882e-10, 2.2132801437183713e-10, 
    2.2087567964009923e-10, 2.2050280977267378e-10, 2.2019816629448769e-10, 
    2.199473244784156e-10, 2.1973356978291416e-10, 2.1953895180434804e-10, 
    2.1934535621269435e-10, 2.1913560212634107e-10, 2.1889443446590004e-10, 
    2.1860940555569719e-10, 2.1827155108587128e-10, 2.1787585470496806e-10, 
    2.1742143007335693e-10, 2.1691146183558915e-10, 2.1635284685166801e-10, 
    2.157556309037861e-10, 2.1513220740816907e-10, 2.1449639620757852e-10, 
    2.1386242692308881e-10, 2.1324394054240216e-10, 2.1265302827328533e-10, 
    2.1209944333261164e-10, 2.11589986837933e-10, 2.1112814843412963e-10, 
    2.1071397668415329e-10, 2.1034422843530437e-10, 2.1001271554547335e-10, 
    2.0971085412662326e-10, 2.0942832908935865e-10, 2.0915384985661078e-10, 
    2.0887588242175163e-10, 2.0858336702782468e-10, 2.0826632905776506e-10, 
    2.0791638805545874e-10, 2.0752709512094618e-10, 2.0709415354202226e-10, 
    2.0661547106142272e-10, 2.0609109189332378e-10, 2.0552299517193314e-10, 
    2.0491481580653479e-10, 2.0427146807162961e-10, 2.0359874797434662e-10, 
    2.0290288720491594e-10, 2.0219012891422806e-10, 2.0146631565830029e-10, 
    2.007365420860493e-10, 2.0000484779749814e-10, 1.9927403129908613e-10, 
    1.9854553184144683e-10, 1.9781944385535228e-10, 1.9709463094220412e-10, 
    1.9636896694800365e-10, 1.9563966266455598e-10, 1.9490369954702239e-10, 
    1.9415830395512649e-10, 1.9340147704252625e-10, 1.9263246153823692e-10, 
    1.91852182771114e-10, 1.9106356347724408e-10, 1.9027169333009089e-10, 
    1.894837883126884e-10, 1.8870897819217063e-10, 1.879578848800948e-10, 
    1.872420428067136e-10, 1.8657318004896972e-10, 1.8596247044447593e-10, 
    1.8541978440274196e-10, 1.84953051295241e-10, 1.8456777325705091e-10, 
    1.8426675734285544e-10, 1.8405006415230968e-10, 1.839151985517106e-10, 
    1.8385747376283434e-10, 1.8387052540720281e-10, 1.8394685956588754e-10, 
    1.8407841158874246e-10, 1.8425698904400599e-10, 1.8447459261769441e-10, 
    1.8472355011120684e-10, 1.8499648980198039e-10, 1.8528614757316228e-10, 
    1.8558509765448172e-10, 1.8588540584280724e-10, 1.861783431349941e-10, 
    1.8645415902518748e-10, 1.8670201555021264e-10, 1.8691005989206494e-10, 
    1.8706569557539925e-10, 1.8715600906504477e-10, 1.8716833407463446e-10, 
    1.8709089194718485e-10, 1.8691349361757477e-10, 1.8662819239780777e-10, 
    1.8622989785133576e-10, 1.8571684695320102e-10, 1.8509095408674346e-10, 
    1.8435795777791973e-10, 1.8352741173839161e-10, 1.8261245936205347e-10, 
    1.8162945818554949e-10, 1.8059740508995242e-10, 1.7953724628729617e-10, 
    1.7847105164044107e-10, 1.7742112611503721e-10, 1.7640904986475718e-10, 
    1.7545474838605887e-10, 1.7457558595120855e-10, 1.7378558089572401e-10, 
    1.7309473269189477e-10, 1.7250856983872661e-10, 1.7202790127057388e-10, 
    1.7164882364870155e-10, 1.7136298674404454e-10, 1.7115811266464575e-10, 
    1.7101870848331824e-10, 1.7092698185720629e-10, 1.7086384869804628e-10, 
    1.7080999852554653e-10, 1.7074690448278125e-10, 1.706577596225524e-10, 
    1.7052823384025651e-10, 1.7034703924505842e-10, 1.7010625710212798e-10, 
    1.6980145383630804e-10, 1.694315718649819e-10, 1.6899866591621951e-10, 
    1.6850749913007054e-10, 1.6796508402064707e-10, 1.673802004977767e-10, 
    1.6676294630854489e-10, 1.6612432277224573e-10, 1.6547591295666036e-10, 
    1.6482960144706528e-10, 1.6419734920912302e-10, 1.6359096351705224e-10, 
    1.6302187110481017e-10, 1.6250079632404754e-10, 1.6203740056905103e-10, 
    1.6163982167658917e-10, 1.6131416605936714e-10, 1.6106394194273627e-10, 
    1.6088955065540685e-10, 1.6078784878690187e-10, 1.6075189111170761e-10, 
    1.6077087295272062e-10, 1.6083037765437822e-10, 1.6091291385630819e-10, 
    1.609987638002631e-10, 1.6106707243171793e-10, 1.6109715846498735e-10, 
    1.610698917200162e-10, 1.6096907365889756e-10, 1.6078264646733634e-10, 
    1.6050366323460583e-10, 1.6013088036835928e-10, 1.5966893403842496e-10, 
    1.5912805488362677e-10, 1.5852336287281909e-10, 1.5787374880529529e-10, 
    1.5720050852069742e-10, 1.565257756853415e-10, 1.5587094246521337e-10, 
    1.5525515887345193e-10, 1.5469405452615758e-10, 1.5419874914336885e-10, 
    1.5377524639736109e-10, 1.5342417686316424e-10, 1.5314095089320921e-10, 
    1.5291620885967158e-10, 1.5273657580809893e-10, 1.5258556385338866e-10, 
    1.5244462449681202e-10, 1.5229420858000839e-10, 1.5211481258252557e-10, 
    1.5188791507978674e-10, 1.5159681550177497e-10, 1.5122730321143923e-10, 
    1.5076819362913147e-10, 1.5021169053774213e-10, 1.4955362110669697e-10, 
    1.4879352454790193e-10, 1.4793463467603866e-10, 1.4698373913900924e-10, 
    1.4595095419745206e-10, 1.448493983474341e-10, 1.4369478674788895e-10, 
    1.4250492626069818e-10, 1.4129915284091168e-10, 1.400976690173792e-10, 
    1.3892084747379223e-10, 1.3778847624334888e-10, 1.3671901103172695e-10, 
    1.3572882470862268e-10, 1.3483154459795643e-10, 1.3403747951922317e-10, 
    1.3335320436191189e-10, 1.3278130147044776e-10, 1.3232032642455837e-10, 
    1.3196496574464339e-10, 1.3170641274189185e-10, 1.3153290889819966e-10, 
    1.3143045612192915e-10, 1.3138359041841939e-10, 1.313762293459707e-10, 
    1.3139249611836424e-10, 1.3141747581570715e-10, 1.3143785327292559e-10, 
    1.3144241141801509e-10, 1.3142234108392187e-10, 1.3137137825311191e-10, 
    1.3128575084188756e-10, 1.311639756022126e-10, 1.3100649492603255e-10, 
    1.3081524408064144e-10, 1.3059314328986269e-10, 1.3034359954110658e-10, 
    1.30070030597095e-10, 1.2977549621950202e-10, 1.2946241669272515e-10, 
    1.2913246219236115e-10, 1.2878656310552924e-10, 1.2842508216448965e-10, 
    1.280480853447409e-10, 1.2765570689106278e-10, 1.272485200320487e-10, 
    1.2682789697784165e-10, 1.2639626956974764e-10, 1.2595727160243673e-10, 
    1.2551569716145701e-10, 1.2507729360191312e-10, 1.2464837159015123e-10, 
    1.2423528498004015e-10, 1.2384380959529682e-10, 1.2347851368831085e-10, 
    1.2314217100860546e-10, 1.2283531277717661e-10, 1.2255595304963668e-10, 
    1.2229955934015331e-10, 1.2205927371819303e-10, 1.2182638718095072e-10, 
    1.2159100209478305e-10, 1.2134287903707742e-10, 1.2107232990002953e-10, 
    1.2077112923916952e-10, 1.204333042061968e-10, 1.2005577402782274e-10, 
    1.1963874319417283e-10, 1.191858346978946e-10, 1.1870393676305226e-10, 
    1.1820279034069614e-10, 1.176943535532594e-10, 1.171919976412575e-10, 
    1.1670961780558335e-10, 1.1626072956473952e-10, 1.1585760908219681e-10, 
    1.1551057653851687e-10, 1.152274332937657e-10, 1.1501311448801013e-10, 
    1.1486953721383925e-10, 1.1479566965387069e-10, 1.1478776787670632e-10, 
    1.1483976622233268e-10, 1.1494377183749995e-10, 1.1509061873954894e-10, 
    1.1527042902290461e-10, 1.154731663048773e-10, 1.1568910820435863e-10, 
    1.1590925918697085e-10, 1.1612564558872316e-10, 1.1633151823571685e-10, 
    1.1652143672208249e-10, 1.1669126755017429e-10, 1.1683809247267415e-10, 
    1.169600593329154e-10, 1.1705619914692647e-10, 1.1712623173143866e-10, 
    1.1717036719563985e-10, 1.171891633588333e-10, 1.1718341206340475e-10, 
    1.171540967600398e-10, 1.1710238653703805e-10, 1.1702969569186709e-10, 
    1.1693776882630493e-10, 1.1682877810927778e-10, 1.1670541050316311e-10, 
    1.1657092186924332e-10, 1.1642914376316307e-10, 1.162844173712044e-10, 
    1.1614146077772377e-10, 1.1600516981052531e-10, 1.1588036430857525e-10, 
    1.1577150103388946e-10, 1.1568236790467925e-10, 1.1561580789203073e-10, 
    1.1557346899125973e-10, 1.1555563053180267e-10, 1.1556109144069611e-10, 
    1.1558715240314367e-10, 1.156296848010596e-10, 1.1568326468837074e-10, 
    1.1574139028831925e-10, 1.157967421098512e-10, 1.1584147501076254e-10, 
    1.1586754374633811e-10, 1.1586703027642639e-10, 1.1583247884831694e-10, 
    1.1575722047132107e-10, 1.1563569679371631e-10, 1.1546375458863561e-10, 
    1.1523892956211491e-10, 1.1496068123870371e-10, 1.1463058268083242e-10, 
    1.1425242966322244e-10, 1.1383225859794126e-10, 1.1337824465717692e-10, 
    1.1290046645224708e-10, 1.1241053850052114e-10, 1.1192111237244179e-10, 
    1.1144526072677648e-10, 1.1099578845886347e-10, 1.1058452253263966e-10, 
    1.1022161990851755e-10, 1.0991494873274987e-10, 1.0966961110404818e-10, 
    1.0948764387099031e-10, 1.0936790702436075e-10, 1.0930619256643552e-10, 
    1.0929553113364898e-10, 1.0932665419848719e-10, 1.0938859406059393e-10, 
    1.094693503241514e-10, 1.0955656032275128e-10, 1.0963813777644877e-10, 
    1.0970281801199666e-10, 1.0974057216983457e-10, 1.0974288690469033e-10, 
    1.0970290400824754e-10, 1.0961543278854658e-10, 1.09476840574654e-10, 
    1.0928489310294768e-10, 1.0903855386784357e-10, 1.0873778140408725e-10, 
    1.0838335519602159e-10, 1.0797674637739569e-10, 1.0752004188453487e-10, 
    1.0701591745847014e-10, 1.0646763606006184e-10, 1.0587906876038476e-10, 
    1.0525470169067011e-10, 1.045996107037337e-10, 1.0391938554338295e-10, 
    1.0321999682048737e-10, 1.0250760029441641e-10, 1.0178830009001728e-10, 
    1.0106786429304994e-10, 1.0035145373266206e-10, 9.9643362380460514e-11, 
    9.8946824501983208e-11, 9.8263903349865013e-11, 9.7595481776979784e-11, 
    9.6941385810133953e-11, 9.6300612783726473e-11, 9.5671670180492023e-11, 
    9.5052991864070424e-11, 9.444337914263625e-11, 9.3842442384995173e-11, 
    9.325097216981839e-11, 9.2671190655339776e-11, 9.2106866781919247e-11, 
    9.1563242422370689e-11, 9.1046762550166088e-11, 9.0564647783519625e-11, 
    9.0124316599050085e-11, 8.9732723160094214e-11, 8.9395659730619339e-11, 
    8.9117119274175408e-11, 8.8898752920042339e-11, 8.8739509090534494e-11, 
    8.8635495615518426e-11, 8.8580066263351125e-11, 8.8564156452777597e-11, 
    8.8576832509391081e-11, 8.8606009681369345e-11, 8.8639289058790841e-11, 
    8.8664837456661705e-11, 8.8672234031066073e-11, 8.8653232225333334e-11, 
    8.860235701487654e-11, 8.851730412468789e-11, 8.8399116364340457e-11, 
    8.8252105376759042e-11, 8.8083557717779397e-11, 8.7903210147810099e-11, 
    8.7722562442973546e-11, 8.7554067906536055e-11, 8.7410249800592785e-11, 
    8.7302819373977367e-11, 8.7241854374058076e-11, 8.7235094695276465e-11, 
    8.728740782415874e-11, 8.7400460150253388e-11, 8.7572617255949294e-11, 
    8.7799064008364269e-11, 8.8072145493712833e-11, 8.8381873599354817e-11, 
    8.871657590991205e-11, 8.906360156409382e-11, 8.9410053729547893e-11, 
    8.9743472076115033e-11, 9.0052426659343178e-11, 9.0326978110043598e-11, 
    9.0558982685585208e-11, 9.0742247265714155e-11, 9.0872519104804332e-11, 
    9.094733806768874e-11, 9.0965788490744294e-11, 9.0928185150662362e-11, 
    9.0835733107230763e-11, 9.0690208155642281e-11, 9.0493706908769362e-11, 
    9.0248488117287055e-11, 8.9956941618739231e-11, 8.9621680369155531e-11, 
    8.9245752015851901e-11, 8.883294132258342e-11, 8.8388108948351688e-11, 
    8.7917524393584708e-11, 8.7429111036245891e-11, 8.6932562972084907e-11, 
    8.6439271261352019e-11, 8.5962039022464261e-11, 8.5514583543245723e-11, 
    8.5110854307140904e-11, 8.476421145058037e-11, 8.4486552603795794e-11, 
    8.4287454115562629e-11, 8.417343827298126e-11, 8.4147420692046363e-11, 
    8.4208400467367095e-11, 8.4351441117242405e-11, 8.4567912165019697e-11, 
    8.4845995174781627e-11, 8.5171383470285645e-11, 8.5528116738081925e-11, 
    8.5899466804529484e-11, 8.6268812616042983e-11, 8.6620421643039866e-11, 
    8.694011192490486e-11, 8.7215734388008521e-11, 8.743749720011777e-11, 
    8.7598102040353298e-11, 8.7692742488950198e-11, 8.771897535717048e-11, 
    8.7676502108768433e-11, 8.7566892295958506e-11, 8.7393284150893141e-11, 
    8.7160075372001343e-11, 8.6872633244356153e-11, 8.6537028693764234e-11, 
    8.6159813458793185e-11, 8.5747818661070023e-11, 8.5308002766729605e-11, 
    8.4847337370175438e-11, 8.4372726097057158e-11, 8.3890940191137975e-11, 
    8.3408592869128118e-11, 8.2932120339437404e-11, 8.2467761290408205e-11, 
    8.2021541486588694e-11, 8.1599225728685186e-11, 8.1206251099157213e-11, 
    8.0847621961374796e-11, 8.0527770055202451e-11, 8.0250393548589615e-11, 
    8.0018266689418599e-11, 7.983307096216112e-11, 7.9695233377918169e-11, 
    7.9603825892912138e-11, 7.9556528826073981e-11, 7.9549681624397197e-11, 
    7.9578408369971273e-11, 7.9636847096199081e-11, 7.9718431289703675e-11, 
    7.9816232740632652e-11, 7.9923299302923084e-11, 8.0032998697763378e-11, 
    8.0139294282794724e-11, 8.0236956069395503e-11, 8.0321692748176652e-11, 
    8.0390187477986502e-11, 8.0440037073498291e-11, 8.0469651275042303e-11, 
    8.047809143705899e-11, 8.0464916409514019e-11, 8.0430032446095654e-11, 
    8.03735977299353e-11, 8.0295969210409638e-11, 8.0197724299777152e-11, 
    8.0079723810116482e-11, 7.994322312188579e-11, 7.9789981707033416e-11, 
    7.9622374051647806e-11, 7.9443455562540781e-11, 7.9256970094444343e-11, 
    7.9067300183877956e-11, 7.8879361734035438e-11, 7.8698422458972114e-11, 
    7.852991624467067e-11, 7.8379249395852676e-11, 7.8251622611865842e-11, 
    7.8151900479707778e-11, 7.8084534615995596e-11, 7.8053538169249391e-11, 
    7.8062505646052349e-11, 7.8114649019286457e-11, 7.8212830810898311e-11, 
    7.8359549456560458e-11, 7.8556886904537998e-11, 7.8806355151432077e-11, 
    7.9108697456351101e-11, 7.9463625806887373e-11, 7.9869540581215805e-11, 
    8.0323264820231336e-11, 8.0819859561794836e-11, 8.1352532537875289e-11, 
    8.1912705567628651e-11, 8.2490236530748056e-11, 8.3073818118483578e-11, 
    8.3651489699442022e-11, 8.4211273288106972e-11, 8.4741846692506951e-11, 
    8.523319748401405e-11, 8.567719069822485e-11, 8.6068014850082423e-11, 
    8.6402434114083499e-11, 8.6679852468206997e-11, 8.690216676976743e-11, 
    8.7073439440759807e-11, 8.7199404054854571e-11, 8.7286876089076659e-11, 
    8.7343093975565739e-11, 8.7375070420322054e-11, 8.7388969283845283e-11, 
    8.7389588490956447e-11, 8.737994746771417e-11, 8.7361024006116166e-11, 
    8.7331629670600209e-11, 8.7288451621045259e-11, 8.7226228169327451e-11, 
    8.7138068751954603e-11, 8.7015885190030473e-11, 8.68509271182928e-11, 
    8.6634384869838265e-11, 8.6358043565096605e-11, 8.6014935700398118e-11, 
    8.5599971606849976e-11, 8.5110493026500861e-11, 8.4546718377595452e-11, 
    8.3912015958856203e-11, 8.3213005390087493e-11, 8.2459430755868816e-11, 
    8.1663823745768329e-11, 8.0840945937639634e-11, 8.0007056156869178e-11, 
    7.9179060223794379e-11, 7.8373585518644834e-11, 7.7606082201301605e-11, 
    7.6890023500723185e-11, 7.6236264114901748e-11, 7.5652648178892369e-11, 
    7.5143862599927918e-11, 7.4711570978861027e-11, 7.4354798203427479e-11, 
    7.4070509535524999e-11, 7.385432329924112e-11, 7.370127351060411e-11, 
    7.3606524179360689e-11, 7.3565976879381139e-11, 7.3576702745617918e-11, 
    7.3637158805840999e-11, 7.3747182121825344e-11, 7.3907776342921955e-11, 
    7.412073444724408e-11, 7.4388149665727066e-11, 7.4711854155384318e-11, 
    7.5092884129262086e-11, 7.553099200322585e-11, 7.6024260270896574e-11, 
    7.6568839375571957e-11, 7.7158819956871526e-11, 7.7786231417061104e-11, 
    7.8441168094234281e-11, 7.9112004295519688e-11, 7.9785693890802801e-11, 
    8.044813641550059e-11, 8.1084590442614296e-11, 8.1680110909622507e-11, 
    8.2220022587668219e-11, 8.2690417205960556e-11, 8.3078655483661104e-11, 
    8.3373853001440768e-11, 8.356735777769538e-11, 8.3653173641281999e-11, 
    8.36283079141019e-11, 8.3493000079853522e-11, 8.3250829620443921e-11, 
    8.2908643167106859e-11, 8.2476316120065759e-11, 8.1966336977177325e-11, 
    8.1393227554619312e-11, 8.0772827420758039e-11, 8.0121498300913562e-11, 
    7.945529819332607e-11, 7.8789184921134463e-11, 7.8136303475275213e-11, 
    7.7507429655213778e-11, 7.6910583617481348e-11, 7.6350861459109124e-11, 
    7.5830466887367084e-11, 7.5348958755829664e-11, 7.4903650472793233e-11, 
    7.4490144748127012e-11, 7.4102957950554164e-11, 7.3736154664967481e-11, 
    7.3383968627498785e-11, 7.3041353457871779e-11, 7.2704413212526584e-11, 
    7.23707186557707e-11, 7.2039450016294162e-11, 7.1711401112893382e-11, 
    7.1388823913098219e-11, 7.1075152379250841e-11, 7.0774622428486211e-11, 
    7.0491836135713475e-11, 7.0231300661544248e-11, 6.9996991932949346e-11, 
    6.9791984660731627e-11, 6.9618179018833898e-11, 6.9476139785137868e-11, 
    6.9365075161451757e-11, 6.9282938628329814e-11, 6.9226643062143078e-11, 
    6.9192366057709061e-11, 6.9175909079679476e-11, 6.9173078784012368e-11, 
    6.9180061752249736e-11, 6.9193746315190335e-11, 6.9211991701934991e-11, 
    6.9233813352289373e-11, 6.9259478030983392e-11, 6.929050926181894e-11, 
    6.9329604538196276e-11, 6.9380462754330692e-11, 6.9447542208106796e-11, 
    6.9535740643731284e-11, 6.9650030694985471e-11, 6.9795039097231339e-11, 
    6.9974610304203377e-11, 7.0191373140810002e-11, 7.0446328026517704e-11, 
    7.0738489986405946e-11, 7.1064622120957061e-11, 7.1419087059359987e-11, 
    7.1793833421412683e-11, 7.2178528656207e-11, 7.2560857938934345e-11, 
    7.2926960656127562e-11, 7.3261998178760714e-11, 7.3550816601965944e-11, 
    7.377867352230233e-11, 7.393197845214972e-11, 7.3999016849656238e-11, 
    7.3970605039128058e-11, 7.3840654262948532e-11, 7.3606602745635902e-11, 
    7.3269702469562056e-11, 7.2835137723376097e-11, 7.231197860656588e-11, 
    7.1712950385255067e-11, 7.1054055990265058e-11, 7.0354014299004813e-11, 
    6.9633585554702024e-11, 6.8914754021961156e-11, 6.8219843999159958e-11, 
    6.7570563585561312e-11, 6.6987050229667469e-11, 6.6486938533271345e-11, 
    6.6084526947512419e-11, 6.5790057033567933e-11, 6.5609192162380394e-11, 
    6.5542700285838589e-11, 6.558638311199837e-11, 6.573126205066195e-11, 
    6.5964014825004793e-11, 6.6267629187860759e-11, 6.6622260698425489e-11, 
    6.7006212118290066e-11, 6.7397009731500224e-11, 6.7772489647759242e-11, 
    6.8111857356632165e-11, 6.8396653543301213e-11, 6.8611598802071611e-11, 
    6.8745276152507698e-11, 6.8790630631890292e-11,
  // Sqw-total(8, 0-1999)
    0.020924657801382866, 0.020921578802110482, 0.020912419328806341, 
    0.020897406400730657, 0.020876900313328353, 0.020851369054497974, 
    0.020821355409662574, 0.020787439401983913, 0.020750199089240751, 
    0.020710172855287555, 0.020667826169496008, 0.020623525345387712, 
    0.020577520142438768, 0.02052993618528973, 0.02048077721069114, 
    0.020429936199842676, 0.020377213622058563, 0.020322340404125554, 
    0.020265002922431337, 0.020204867329177843, 0.020141600863363501, 
    0.020074888411313219, 0.020004443382307922, 0.01993001283891432, 
    0.019851377646517662, 0.019768349068699717, 0.019680763646169976, 
    0.01958847830653487, 0.019491367454467192, 0.01938932332553242, 
    0.019282260228601442, 0.019170122553636423, 0.01905289569613677, 
    0.018930618452844151, 0.018803395060563673, 0.018671404933949656, 
    0.018534908323118864, 0.018394246533116269, 0.018249835965249872, 
    0.018102155970385132, 0.017951731248306416, 0.017799110186960711, 
    0.017644841025321933, 0.017489447982029119, 0.017333409488601362, 
    0.017177140405691006, 0.017020979622279629, 0.016865183808078523, 
    0.016709927394630373, 0.016555308193256409, 0.016401357503887208, 
    0.016248053194836649, 0.016095334078218362, 0.015943113974222104, 
    0.015791294122317074, 0.015639773004025404, 0.015488453118600183, 
    0.015337244723580145, 0.015186066948712476, 0.015034846964710592, 
    0.014883518013520015, 0.014732017086840321, 0.014580282900785049, 
    0.014428254599269403, 0.014275871376344069, 0.014123072984688255, 
    0.013969800929343598, 0.013816000052071566, 0.013661620194795427, 
    0.013506617677830537, 0.013350956417358829, 0.013194608610448647, 
    0.013037555010783223, 0.01287978488714633, 0.01272129579213703, 
    0.012562093272490247, 0.012402190633800355, 0.012241608843741524, 
    0.012080376630557757, 0.011918530814888879, 0.01175611690392845, 
    0.011593189972454948, 0.011429815846366449, 0.011266072581279481, 
    0.01110205218492195, 0.010937862467083795, 0.010773628822118733, 
    0.010609495670853855, 0.010445627230080277, 0.010282207257556596, 
    0.010119437453052304, 0.0099575342871496188, 0.0097967241740419386, 
    0.00963723708617663, 0.0094792989025224515, 0.0093231229596351453, 
    0.0091689014079603531, 0.0090167970437864467, 0.0088669362790066101, 
    0.008719403827375613, 0.008574239539511485, 0.0084314376303125764, 
    0.0082909483369824569, 0.008152681848712609, 0.0080165141815343646, 
    0.0078822945485509856, 0.00774985370362174, 0.0076190127152693772, 
    0.0074895916511482008, 0.0073614177124239517, 0.0072343324411514543, 
    0.0071081977218530228, 0.0069829004019829046, 0.0068583554573961739, 
    0.0067345077222440292, 0.0066113322827800348, 0.0064888336969510605, 
    0.0063670442427443338, 0.0062460214157149876, 0.0061258448896096551, 
    0.0060066131259149756, 0.0058884397739799059, 0.0057714499513744537, 
    0.0056557764444810522, 0.0055415558322477552, 0.0054289245199965171, 
    0.005318014679763082, 0.0052089501282213705, 0.005101842226527608, 
    0.00499678594728078, 0.004893856308228986, 0.0047931054062850089, 
    0.0046945602877811708, 0.0045982218562644296, 0.0045040649492702331, 
    0.0044120396194212144, 0.0043220735475517176, 0.0042340754138374421, 
    0.0041479389737923917, 0.0040635475418918515, 0.0039807785820265206, 
    0.0038995081385949505, 0.003819614905126929, 0.0037409838042519765, 
    0.0036635090272648628, 0.003587096539131209, 0.003511666086152099, 
    0.0034371527461293599, 0.0033635080392527294, 0.0032907005822738929, 
    0.0032187162321640557, 0.0031475576416731504, 0.0030772431482683506, 
    0.003007804944807368, 0.0029392865336721574, 0.0028717395386616816, 
    0.0028052200289747438, 0.0027397845832497639, 0.0026754863755208661, 
    0.0026123715886772229, 0.0025504764488366921, 0.0024898251257860658, 
    0.0024304286655549854, 0.0023722850210139085, 0.0023153801377081614, 
    0.0022596899484943369, 0.0022051830444582473, 0.0021518237309458826, 
    0.002099575152372953, 0.0020484021794373031, 0.0019982737947182028, 
    0.00194916478092834, 0.001901056601086884, 0.0018539374509973976, 
    0.0018078015510122293, 0.001762647816803386, 0.0017184781007196402, 
    0.0016752952222929183, 0.0016331010078231873, 0.0015918945370699932, 
    0.0015516707547662803, 0.0015124195524693093, 0.0014741253693498599, 
    0.0014367673057385853, 0.0014003196962479869, 0.0013647530539548161, 
    0.0013300352753076164, 0.0012961329870180267, 0.0012630129195045129, 
    0.0012306432037536524, 0.0011989945065927498, 0.0011680409403371135, 
    0.001137760704165211, 0.0011081364347718871, 0.0010791552620416469, 
    0.0010508085815036795, 0.0010230915693705549, 0.0009960024782857482, 
    0.00096954176258613441, 0.00094371109068701786, 0.00091851230854986189, 
    0.00089394642133231903, 0.00087001265947411657, 0.00084670769011161557, 
    0.00082402502474087725, 0.00080195465993513997, 0.00078048297070726195, 
    0.00075959285730589307, 0.00073926412762395904, 0.0007194740807762764, 
    0.00070019824430916553, 0.00068141120901918622, 0.000663087501956041, 
    0.00064520243972602295, 0.00062773291001048536, 0.00061065803820866489, 
    0.00059395970707016232, 0.00057762290890437577, 0.00056163592143939115, 
    0.000545990308947543, 0.00053068075945381338, 0.00051570477654776605, 
    0.00050106225052455307, 0.00048675493832696164, 0.0004727858850400337, 
    0.00045915882141459101, 0.00044587757190636348, 0.00043294550585177606, 
    0.00042036506057453298, 0.000408137359512162, 0.00039626194116291563, 
    0.00038473660630360384, 0.00037355738221171828, 0.00036271859432907602, 
    0.00035221302869261608, 0.00034203216317095915, 0.00033216644250654454, 
    0.00032260557154319017, 0.0003133388027209035, 0.0003043551976220907, 
    0.00029564384755420396, 0.00028719404424824228, 0.00027899539808592418, 
    0.00027103790720313332, 0.00026331198577197161, 0.00025580846326421724, 
    0.00024851856821068497, 0.000241433909745207, 0.00023454646812052357, 
    0.00022784860170256909, 0.00022133307320399391, 0.00021499309280231883, 
    0.00020882237108946273, 0.00020281517129024454, 0.00019696634849053618, 
    0.00019127136409454772, 0.00018572626639585483, 0.00018032763264027741, 
    0.00017507247358494328, 0.00016995810740326695, 0.00016498201486529672, 
    0.00016014169116739685, 0.00015543451099211568, 0.00015085762213267294, 
    0.00014640787951835938, 0.00014208182631164404, 0.00013787572275895764, 
    0.00013378561761555842, 0.00012980745210375318, 0.00012593718315526226, 
    0.00012217091145580577, 0.00011850500052551342, 0.00011493617538722408, 
    0.00011146159273904797, 0.00010807887831113915, 0.00010478613065299288, 
    0.00010158189351826327, 9.846510105762135e-05, 9.5435001180656915e-05, 
    9.2491062871825997e-05, 8.9632873208672577e-05, 8.6860029617817332e-05, 
    8.4172032732089818e-05, 8.156818518458452e-05, 7.9047501758195096e-05, 
    7.6608636358850267e-05, 7.4249831085253771e-05, 7.1968892019648901e-05, 
    6.9763195115361764e-05, 6.7629723677023823e-05, 6.5565136519445556e-05, 
    6.3565863184639101e-05, 6.1628219917376681e-05, 5.9748537814522813e-05, 
    5.7923293011400104e-05, 5.6149228208838851e-05, 5.4423455404183504e-05, 
    5.2743531346362308e-05, 5.1107499813678561e-05, 4.9513898016038448e-05, 
    4.7961727869435484e-05, 4.6450396176149122e-05, 4.4979630492270003e-05, 
    4.3549379382147001e-05, 4.2159706666450035e-05, 4.0810689123107683e-05, 
    3.950232598281461e-05, 3.8234466672251935e-05, 3.700676087284529e-05, 
    3.5818632395241948e-05, 3.4669275924905818e-05, 3.3557673637433274e-05, 
    3.2482627202111928e-05, 3.1442799891882346e-05, 3.0436763403919304e-05, 
    2.9463044493376105e-05, 2.8520167489901781e-05, 2.760669002109048e-05, 
    2.6721230610481937e-05, 2.5862488067392647e-05, 2.5029253590444529e-05, 
    2.4220417168624811e-05, 2.3434970140887271e-05, 2.2672005686748231e-05, 
    2.1930718632370769e-05, 2.1210405374717296e-05, 2.0510464071063257e-05, 
    1.9830394635133581e-05, 1.9169797625051567e-05, 1.8528370873864279e-05, 
    1.7905902728925261e-05, 1.7302261022412968e-05, 1.6717377342743263e-05, 
    1.6151226744177967e-05, 1.560380363162597e-05, 1.5075095105581942e-05, 
    1.4565053473333192e-05, 1.4073569876379969e-05, 1.360045102211279e-05, 
    1.3145400841079454e-05, 1.270800854080034e-05, 1.2287744035548588e-05, 
    1.1883961150315927e-05, 1.1495908386548374e-05, 1.1122746454107692e-05, 
    1.0763571272711368e-05, 1.0417440768177589e-05, 1.0083403565548915e-05, 
    9.760527624637855e-06, 9.4479269726136159e-06, 9.14478494211748e-06, 
    8.8503726905898846e-06, 8.5640622124288778e-06, 8.2853335146141645e-06, 
    8.0137760609988867e-06, 7.74908496380518e-06, 7.4910526846748397e-06, 
    7.2395571910484151e-06, 6.9945475966181858e-06, 6.7560283121311126e-06, 
    6.5240426641902405e-06, 6.2986568299320009e-06, 6.0799448045278323e-06, 
    5.867974983764404e-06, 5.6627988125886571e-06, 5.4644418261322198e-06, 
    5.2728972875617437e-06, 5.0881225042776607e-06, 4.9100377754313802e-06, 
    4.7385277914662291e-06, 4.5734451742433245e-06, 4.4146157256219503e-06, 
    4.261844854215286e-06, 4.1149245884785745e-06, 3.9736405677442462e-06, 
    3.8377784374910965e-06, 3.707129157911384e-06, 3.5814928593966574e-06, 
    3.4606810304948593e-06, 3.3445169888923921e-06, 3.2328347463317712e-06, 
    3.125476521152401e-06, 3.0222892645477939e-06, 2.923120643101843e-06, 
    2.8278149556481572e-06, 2.7362094584719133e-06, 2.6481315298853866e-06, 
    2.5633970286485521e-06, 2.4818100943999966e-06, 2.4031645103694312e-06, 
    2.3272466064236031e-06, 2.2538395359707488e-06, 2.1827286243564522e-06, 
    2.1137073741424189e-06, 2.046583635233137e-06, 1.9811854172162163e-06, 
    1.9173658418163302e-06, 1.8550068063406851e-06, 1.7940210461273398e-06, 
    1.7343524334773632e-06, 1.6759745133690528e-06, 1.6188874338832418e-06, 
    1.5631135619138726e-06, 1.5086921690180559e-06, 1.4556736184512605e-06, 
    1.4041134829935419e-06, 1.3540669785780421e-06, 1.3055840238774131e-06, 
    1.2587051440243369e-06, 1.2134583434441228e-06, 1.1698569891699774e-06, 
    1.1278986812895841e-06, 1.08756504254398e-06, 1.0488223338864746e-06, 
    1.0116227903473547e-06, 9.7590656598583543e-07, 9.4160417077832926e-07, 
    9.0863927306792339e-07, 8.7693172686793096e-07, 8.4640066774576893e-07, 
    8.1696750775837808e-07, 7.8855865640085856e-07, 7.6110780429044531e-07, 
    7.3455763351478308e-07, 7.0886086142611931e-07, 6.8398058026120093e-07, 
    6.5988991546017381e-07, 6.3657108380297898e-07, 6.1401397908291983e-07, 
    5.9221444296698668e-07, 5.7117238721176705e-07, 5.5088992211626233e-07, 
    5.3136961735085038e-07, 5.1261298257609522e-07, 4.9461921306609072e-07, 
    4.7738420825027502e-07, 4.6089984340236719e-07, 4.4515346080469071e-07, 
    4.3012754584414598e-07, 4.1579956377077405e-07, 4.0214194889663869e-07, 
    3.8912225508017051e-07, 3.7670348802885241e-07, 3.6484464377298023e-07, 
    3.535014704166685e-07, 3.4262745401653537e-07, 3.3217500570612985e-07, 
    3.2209680136546448e-07, 3.1234720098303835e-07, 3.0288365776635211e-07, 
    2.9366801913722667e-07, 2.8466762541143994e-07, 2.7585612576829224e-07, 
    2.6721395393403992e-07, 2.5872843379205232e-07, 2.5039351523253077e-07, 
    2.4220916871552944e-07, 2.3418049146464549e-07, 2.2631659625679706e-07, 
    2.1862936561139663e-07, 2.1113215865683718e-07, 2.0383855658475648e-07, 
    1.9676122515601743e-07, 1.8991096079380786e-07, 1.8329597049890849e-07, 
    1.7692141693777429e-07, 1.7078923876632902e-07, 1.6489823511147595e-07, 
    1.592443826273648e-07, 1.5382133674369213e-07, 1.4862105612019383e-07, 
    1.4363448343079789e-07, 1.3885221597489608e-07, 1.3426510715360226e-07, 
    1.2986475232815624e-07, 1.2564382939535263e-07, 1.2159628201794436e-07, 
    1.1771735065532176e-07, 1.1400347019422311e-07, 1.104520627848588e-07, 
    1.0706125874107356e-07, 1.0382957861455369e-07, 1.0075560557055997e-07, 
    9.7837671677696493e-08, 9.5073575002656072e-08, 9.2460338941653255e-08, 
    8.9994020714390974e-08, 8.7669573706482523e-08, 8.5480767065656288e-08, 
    8.3420165904789283e-08, 8.1479174895981334e-08, 7.9648147126120456e-08, 
    7.7916557441111376e-08, 7.6273236109348863e-08, 7.4706653768587618e-08, 
    7.3205244013177475e-08, 7.175774544495521e-08, 7.0353542300163743e-08, 
    6.8982981439372229e-08, 6.7637644812453892e-08, 6.631055938481516e-08, 
    6.4996331527381736e-08, 6.3691198339990305e-08, 6.2392994720559003e-08, 
    6.1101040396908057e-08, 5.9815956346328264e-08, 5.8539423490243908e-08, 
    5.7273899449235906e-08, 5.6022310445590731e-08, 5.4787736392437666e-08, 
    5.3573106906172172e-08, 5.238092565232417e-08, 5.1213038952174441e-08, 
    5.007046288285665e-08, 4.895328008643621e-08, 4.7860613871110051e-08, 
    4.6790682166199904e-08, 4.5740928415131121e-08, 4.4708220130861293e-08, 
    4.3689100083519851e-08, 4.2680069690786803e-08, 4.1677880884197708e-08, 
    4.0679811073096323e-08, 3.9683897242614612e-08, 3.8689108660126688e-08, 
    3.7695443777458826e-08, 3.6703944105087365e-08, 3.5716626017777727e-08, 
    3.47363388453251e-08, 3.3766564129313146e-08, 3.2811175042246385e-08, 
    3.1874177208712536e-08, 3.0959451650532733e-08, 3.0070518597363968e-08, 
    2.9210337004363996e-08, 2.8381150565683998e-08, 2.7584386350430806e-08, 
    2.6820608478604823e-08, 2.6089525732948774e-08, 2.5390049734516356e-08, 
    2.472039817524537e-08, 2.4078236263251164e-08, 2.3460847954612684e-08, 
    2.286532734596188e-08, 2.2288779057491978e-08, 2.1728515402044751e-08, 
    2.1182237272440481e-08, 2.0648186024029617e-08, 2.0125254609375098e-08, 
    1.9613048941289302e-08, 1.9111893872101263e-08, 1.862278293341807e-08, 
    1.8147275698055471e-08, 1.7687351508732304e-08, 1.7245232105608572e-08, 
    1.6823188430282329e-08, 1.6423347693407047e-08, 1.6047516275171365e-08, 
    1.5697031535484824e-08, 1.5372652383072261e-08, 1.507449408969648e-08, 
    1.4802008791494899e-08, 1.4554008956371188e-08, 1.4328728093226798e-08, 
    1.4123910465673326e-08, 1.39369206469224e-08, 1.3764863187539729e-08, 
    1.3604703550276269e-08, 1.345338246241304e-08, 1.3307917758242908e-08, 
    1.3165489486075876e-08, 1.302350625879427e-08, 1.2879652478607793e-08, 
    1.2731917957910443e-08, 1.257861243318536e-08, 1.241836853071889e-08, 
    1.2250136737517186e-08, 1.2073175866033572e-08, 1.1887041539401236e-08, 
    1.1691574340747499e-08, 1.1486887847939728e-08, 1.1273355848341921e-08, 
    1.1051597013557944e-08, 1.0822455202441861e-08, 1.0586973551703391e-08, 
    1.0346361512548747e-08, 1.0101954861175355e-08, 9.8551702680787702e-09, 
    9.6074569239708749e-09, 9.3602487979437273e-09, 9.1149211454840138e-09, 
    8.8727547781934965e-09, 8.6349105103645835e-09, 8.4024150744446749e-09, 
    8.1761581292627639e-09, 7.956898782572746e-09, 7.7452787939235746e-09, 
    7.5418392072547981e-09, 7.3470369914330035e-09, 7.1612589450083201e-09, 
    6.9848308240865838e-09, 6.8180209832445148e-09, 6.6610387121151627e-09, 
    6.5140285789810508e-09, 6.3770625138208189e-09, 6.2501317758825702e-09, 
    6.1331406062407348e-09, 6.0259031048635434e-09, 5.9281440307920041e-09, 
    5.8395037399105756e-09, 5.7595466240912939e-09, 5.6877721596980586e-09, 
    5.6236272198980611e-09, 5.5665185122935283e-09, 5.5158239888266293e-09, 
    5.4709026070808391e-09, 5.4311020571483636e-09, 5.3957646760682134e-09, 
    5.3642318942588375e-09, 5.3358479815098425e-09, 5.3099637298860265e-09, 
    5.2859408302028948e-09, 5.2631573013871507e-09, 5.2410142742582328e-09, 
    5.2189438984120322e-09, 5.1964180573202812e-09, 5.1729571118024626e-09, 
    5.1481379756036331e-09, 5.1216005254812156e-09, 5.093051696849511e-09, 
    5.0622665469823292e-09, 5.0290861392787459e-09, 4.9934122236322526e-09, 
    4.9551993202311985e-09, 4.9144449600750447e-09, 4.8711793322253796e-09, 
    4.8254554978753244e-09, 4.7773415412155065e-09, 4.7269155494256574e-09, 
    4.6742642119588827e-09, 4.6194850694348399e-09, 4.5626921611989059e-09, 
    4.5040240947053381e-09, 4.4436533655289779e-09, 4.3817953764959169e-09, 
    4.3187157369888957e-09, 4.2547344696031255e-09, 4.1902262489700402e-09, 
    4.1256161074123631e-09, 4.0613707313089068e-09, 3.9979857686211666e-09, 
    3.9359701257838376e-09, 3.8758282987725476e-09, 3.8180421107565922e-09, 
    3.7630529576654363e-09, 3.7112457315509518e-09, 3.6629351505895365e-09, 
    3.6183552070979512e-09, 3.5776519554204973e-09, 3.5408798578200272e-09, 
    3.5080015370613264e-09, 3.4788908642149086e-09, 3.453339017409129e-09, 
    3.4310632641278442e-09, 3.4117180066137909e-09, 3.3949077448355031e-09, 
    3.3802013572142714e-09, 3.3671472698720703e-09, 3.3552888232060317e-09, 
    3.3441793327741818e-09, 3.333396143594689e-09, 3.3225532460886902e-09, 
    3.3113118859873871e-09, 3.2993889142139426e-09, 3.2865625574741888e-09, 
    3.2726756109327421e-09, 3.2576359869336291e-09, 3.2414148491558541e-09, 
    3.224042429478321e-09, 3.2056019263078164e-09, 3.1862216787226291e-09, 
    3.166066079790461e-09, 3.1453254910118267e-09, 3.1242056804738199e-09, 
    3.102917107105839e-09, 3.0816645832592815e-09, 3.0606376614811688e-09, 
    3.0400022560331544e-09, 3.0198937484776712e-09, 3.0004119635550209e-09, 
    2.9816180625059341e-09, 2.9635334973587944e-09, 2.946140820816631e-09, 
    2.9293862474939058e-09, 2.913183559310383e-09, 2.8974190858196049e-09, 
    2.8819572995410329e-09, 2.8666467793527989e-09, 2.8513261612004022e-09, 
    2.8358299646059943e-09, 2.819994089907925e-09, 2.8036610124019952e-09, 
    2.7866845827931588e-09, 2.7689345232552735e-09, 2.750300510216756e-09, 
    2.7306959004425495e-09, 2.7100608916647664e-09, 2.6883650766016003e-09, 
    2.6656091241596676e-09, 2.6418255081774695e-09, 2.6170780545724067e-09, 
    2.5914603134863595e-09, 2.5650926678356703e-09, 2.5381183511887076e-09, 
    2.5106984645144865e-09, 2.4830063194642321e-09, 2.4552213328266607e-09, 
    2.4275228524411841e-09, 2.4000841652348193e-09, 2.3730670456448976e-09, 
    2.3466170226654256e-09, 2.3208596244406395e-09, 2.2958976508619391e-09, 
    2.2718096480492274e-09, 2.2486495062695889e-09, 2.2264472385687617e-09, 
    2.2052107712438687e-09, 2.1849287084705328e-09, 2.1655738066487412e-09, 
    2.1471070316365556e-09, 2.129481860563078e-09, 2.1126486373642798e-09, 
    2.0965585854850912e-09, 2.081167301446636e-09, 2.0664373527788224e-09, 
    2.0523398898958758e-09, 2.0388550319303564e-09, 2.025971103714398e-09, 
    2.0136827159058474e-09, 2.0019879516695642e-09, 1.9908848674122776e-09, 
    1.9803677422156791e-09, 1.9704233700498077e-09, 1.9610278642571514e-09, 
    1.952144209217326e-09, 1.9437209110957274e-09, 1.9356918071636779e-09, 
    1.9279771522769806e-09, 1.9204858330664364e-09, 1.9131186153620084e-09, 
    1.9057720905455865e-09, 1.8983431006008028e-09, 1.8907332385947853e-09, 
    1.8828531762741668e-09, 1.8746264494397686e-09, 1.8659925398780407e-09, 
    1.8569089860162448e-09, 1.8473525061759966e-09, 1.837319011109536e-09, 
    1.8268226429221558e-09, 1.8158938714421e-09, 1.8045768852576575e-09, 
    1.7929264203039925e-09, 1.7810043135807769e-09, 1.7688759427945008e-09, 
    1.7566068361511985e-09, 1.7442595503655435e-09, 1.7318910397506718e-09, 
    1.7195505407893485e-09, 1.7072781105793482e-09, 1.6951037390805798e-09, 
    1.6830471405805428e-09, 1.6711180926999573e-09, 1.6593173393188103e-09, 
    1.6476379486404663e-09, 1.6360670794003279e-09, 1.624588020928322e-09, 
    1.6131824537640361e-09, 1.6018327381941428e-09, 1.5905241793674052e-09, 
    1.5792470547534887e-09, 1.5679983393243258e-09, 1.5567829507092164e-09, 
    1.5456144699224254e-09, 1.5345152301607992e-09, 1.523515798525648e-09, 
    1.5126538314246739e-09, 1.501972432395137e-09, 1.4915180420773286e-09, 
    1.4813381109059653e-09, 1.4714786094157425e-09, 1.461981635598725e-09, 
    1.4528832072840843e-09, 1.4442114233793461e-09, 1.4359850563087793e-09, 
    1.4282126803881441e-09, 1.420892283902546e-09, 1.4140114309544929e-09, 
    1.4075478272105512e-09, 1.4014702917359262e-09, 1.3957399722257251e-09, 
    1.3903117794502326e-09, 1.3851358995289721e-09, 1.3801593713206741e-09, 
    1.3753276260075613e-09, 1.3705860169224089e-09, 1.3658812489774977e-09, 
    1.3611627704145782e-09, 1.3563840362026752e-09, 1.3515036905922283e-09, 
    1.3464865852712428e-09, 1.3413046343639587e-09, 1.3359374264404398e-09, 
    1.3303725805171061e-09, 1.3246057659277975e-09, 1.3186404065438873e-09, 
    1.3124870033674717e-09, 1.3061621628373847e-09, 1.2996873140046102e-09, 
    1.2930872485096613e-09, 1.2863885264862488e-09, 1.2796179140677537e-09, 
    1.2728009150225328e-09, 1.265960565917269e-09, 1.2591165069939732e-09, 
    1.2522844813746322e-09, 1.2454762053688136e-09, 1.2386996620609933e-09, 
    1.2319597222664825e-09, 1.2252590493035638e-09, 1.2185991377240239e-09, 
    1.2119814159186591e-09, 1.2054082310445393e-09, 1.1988836711540507e-09, 
    1.1924140634747377e-09, 1.1860081637601451e-09, 1.1796769460043362e-09, 
    1.1734330658290164e-09, 1.1672900038827118e-09, 1.1612610172807535e-09, 
    1.155357948794882e-09, 1.149590079365491e-09, 1.1439630767285233e-09, 
    1.1384782174844306e-09, 1.1331319002553221e-09, 1.1279155803757248e-09, 
    1.12281608747961e-09, 1.1178163751098083e-09, 1.1128965720380675e-09, 
    1.1080353449709981e-09, 1.103211376478131e-09, 1.098404917151615e-09, 
    1.0935992088611469e-09, 1.0887817540222672e-09, 1.0839452389503211e-09, 
    1.0790881378990051e-09, 1.0742148681440893e-09, 1.0693355651656933e-09, 
    1.0644654223389994e-09, 1.0596237104608468e-09, 1.0548324841441327e-09, 
    1.0501151037704931e-09, 1.0454946169795866e-09, 1.040992154982521e-09, 
    1.0366253736022963e-09, 1.0324071096295892e-09, 1.0283442491881436e-09, 
    1.0244369778026183e-09, 1.0206783634049215e-09, 1.0170544040128863e-09, 
    1.0135444557580356e-09, 1.0101221000110719e-09, 1.0067563393714225e-09, 
    1.0034131098200743e-09, 1.0000569568914024e-09, 9.9665283330423051e-10, 
    9.9316784801809235e-10, 9.8957290557963683e-10, 9.8584406822613197e-10, 
    9.8196361945669183e-10, 9.7792069140010001e-10, 9.7371148101130907e-10, 
    9.6933897742400126e-10, 9.6481228155091187e-10, 9.6014552884986738e-10, 
    9.5535653558872726e-10, 9.5046521664847068e-10, 9.4549197387653096e-10, 
    9.4045610880107172e-10, 9.3537445045277883e-10, 9.3026023500344093e-10, 
    9.2512241892658378e-10, 9.1996537312045876e-10, 9.1478908251483321e-10, 
    9.0958973737723335e-10, 9.0436074711165622e-10, 8.990939796202058e-10, 
    8.9378123548975401e-10, 8.8841570940878851e-10, 8.8299340672389872e-10, 
    8.7751430029987585e-10, 8.7198321523268681e-10, 8.6641027515434476e-10, 
    8.6081095986691955e-10, 8.5520566933289097e-10, 8.4961892590336547e-10, 
    8.4407818005166767e-10, 8.3861240301935565e-10, 8.332504716008592e-10, 
    8.2801956863762169e-10, 8.2294361302284491e-10, 8.1804191688240763e-10, 
    8.1332807615223812e-10, 8.0880924510495626e-10, 8.0448575941999968e-10, 
    8.0035120503613841e-10, 7.9639284488507611e-10, 7.9259245634986015e-10, 
    7.8892743274865077e-10, 7.8537218266171319e-10, 7.8189963603711428e-10, 
    7.7848285837169332e-10, 7.7509658694520292e-10, 7.717186757638075e-10, 
    7.6833125361239757e-10, 7.6492162205176388e-10, 7.6148273230232634e-10, 
    7.5801329293961401e-10, 7.5451741398286052e-10, 7.510039147603555e-10, 
    7.4748525175457292e-10, 7.4397624607666704e-10, 7.4049265049017225e-10, 
    7.3704973504263466e-10, 7.3366094026269693e-10, 7.3033678869351057e-10, 
    7.2708405291029755e-10, 7.2390531715443011e-10, 7.2079886957163745e-10, 
    7.1775898788951035e-10, 7.1477650744335177e-10, 7.1183965818662957e-10, 
    7.0893501535742883e-10, 7.060485499043861e-10, 7.0316660102619087e-10, 
    7.0027676522072327e-10, 6.9736856283293699e-10, 6.9443390215403813e-10, 
    6.9146725720953349e-10, 6.8846562308834244e-10, 6.8542819643758966e-10, 
    6.8235592836244747e-10, 6.7925088615279035e-10, 6.7611563024425331e-10, 
    6.7295257167395042e-10, 6.6976347861584711e-10, 6.665491135661208e-10, 
    6.6330914031718649e-10, 6.6004222987630924e-10, 6.567464623823123e-10, 
    6.5341988571476564e-10, 6.5006126851713317e-10, 6.4667087325235345e-10, 
    6.4325122839566896e-10, 6.3980771656985029e-10, 6.3634897310306658e-10, 
    6.3288693217713952e-10, 6.2943657876303837e-10, 6.2601530564750369e-10, 
    6.2264201337417218e-10, 6.1933593597032819e-10, 6.1611539010343602e-10, 
    6.1299646603398499e-10, 6.0999187666097387e-10, 6.0711000237364128e-10, 
    6.0435427647225752e-10, 6.0172289066959456e-10, 5.9920893217622165e-10, 
    5.9680082625940895e-10, 5.9448314008294339e-10, 5.9223757135648247e-10, 
    5.9004413154975323e-10, 5.8788233238126819e-10, 5.8573238886455854e-10, 
    5.8357626453642035e-10, 5.8139859215969269e-10, 5.7918733679577764e-10, 
    5.7693426675676088e-10, 5.7463512821538586e-10, 5.722896243429699e-10, 
    5.6990113172517661e-10, 5.6747626867996493e-10, 5.6502426095586379e-10, 
    5.6255625552916185e-10, 5.6008453763350208e-10, 5.5762179330052964e-10, 
    5.5518038931583728e-10, 5.5277179641548157e-10, 5.5040611721407322e-10, 
    5.4809181214858366e-10, 5.4583556213396615e-10, 5.436423230812304e-10, 
    5.4151547750874131e-10, 5.3945711132940484e-10, 5.3746829369646847e-10, 
    5.3554939908565853e-10, 5.3370030917984532e-10, 5.3192058842068918e-10, 
    5.3020949315742592e-10, 5.2856589444017479e-10, 5.2698808449701309e-10, 
    5.2547352692884367e-10, 5.2401855629420657e-10, 5.2261814200035049e-10, 
    5.2126569439074762e-10, 5.1995304095423353e-10, 5.1867051796913508e-10, 
    5.1740728299941972e-10, 5.1615175059356688e-10, 5.1489220689678787e-10, 
    5.1361747463491696e-10, 5.1231763985609981e-10, 5.109847032530145e-10, 
    5.0961314780994465e-10, 5.0820029976634211e-10, 5.0674650880363999e-10, 
    5.0525503671301741e-10, 5.0373174624962681e-10, 5.0218453346318213e-10, 
    5.0062261248928468e-10, 4.9905566111745156e-10, 4.9749296725203321e-10, 
    4.9594257270179534e-10, 4.9441058270606228e-10, 4.9290061326320286e-10, 
    4.9141350122738511e-10, 4.8994722117664226e-10, 4.8849709024199487e-10, 
    4.8705615240214417e-10, 4.8561577901154124e-10, 4.8416634621943126e-10, 
    4.8269800173498712e-10, 4.8120137703281649e-10, 4.7966825213093298e-10, 
    4.7809205466202848e-10, 4.7646821991789947e-10, 4.7479432458468813e-10, 
    4.7307005970078557e-10, 4.7129698644333083e-10, 4.6947817567924231e-10, 
    4.6761768913779618e-10, 4.6572003884148702e-10, 4.6378959033345625e-10, 
    4.6183004062209149e-10, 4.5984396170160854e-10, 4.5783250823538596e-10, 
    4.5579527320480901e-10, 4.5373036783092211e-10, 4.5163468569932207e-10, 
    4.4950437937595082e-10, 4.4733546904942747e-10, 4.4512459556644636e-10, 
    4.4286977472364612e-10, 4.4057115251894169e-10, 4.3823160900590544e-10, 
    4.358572020840885e-10, 4.3345731552738358e-10, 4.3104454471741031e-10, 
    4.2863424191611293e-10, 4.2624379613196174e-10, 4.2389164816798698e-10, 
    4.2159617179587008e-10, 4.1937447749811027e-10, 4.1724128745596679e-10, 
    4.1520795689345659e-10, 4.1328177800482921e-10, 4.1146558643551354e-10, 
    4.0975775825710702e-10, 4.0815253755568886e-10, 4.0664070149509977e-10, 
    4.0521043521212107e-10, 4.0384836461774496e-10, 4.0254058137637083e-10, 
    4.0127359585236344e-10, 4.0003508332073932e-10, 3.9881438956689894e-10, 
    3.9760273557310292e-10, 3.9639316692734897e-10, 3.9518022674873048e-10, 
    3.9395951342448683e-10, 3.9272711895151987e-10, 3.9147912817913665e-10, 
    3.9021118542687756e-10, 3.8891826832655849e-10, 3.875946446532031e-10, 
    3.8623407429137523e-10, 3.8483018018345825e-10, 3.8337699841186926e-10, 
    3.8186957302313927e-10, 3.8030458968408478e-10, 3.7868091184373094e-10, 
    3.7700000919959324e-10, 3.7526618607760091e-10, 3.7348663001752713e-10, 
    3.7167122996391907e-10, 3.698322291530322e-10, 3.6798370010728604e-10, 
    3.6614092628792401e-10, 3.6431970934009225e-10, 3.6253567722989839e-10, 
    3.6080361030003458e-10, 3.5913685519017943e-10, 3.5754681646923665e-10, 
    3.5604257934542604e-10, 3.5463063513960423e-10, 3.5331474973222541e-10, 
    3.520959074073286e-10, 3.5097239580536693e-10, 3.4993995191558374e-10, 
    3.4899200888796409e-10, 3.4811999758416079e-10, 3.4731371426201103e-10, 
    3.4656173512930784e-10, 3.4585186267905666e-10, 3.4517158001949945e-10, 
    3.4450851659709746e-10, 3.4385086222561051e-10, 3.4318776045984364e-10, 
    3.4250960331475204e-10, 3.418082726444584e-10, 3.410772669278019e-10, 
    3.4031176898146275e-10, 3.3950861504273032e-10, 3.3866622900886566e-10, 
    3.3778450998889203e-10, 3.3686471294800833e-10, 3.3590931100101382e-10, 
    3.3492188844227287e-10, 3.3390699137539433e-10, 3.3287000354620152e-10, 
    3.3181695417960018e-10, 3.3075429299314142e-10, 3.2968857909018214e-10, 
    3.2862612273657466e-10, 3.2757253891680025e-10, 3.2653230282511024e-10, 
    3.2550829606008722e-10, 3.2450144859583864e-10, 3.2351047808856585e-10, 
    3.2253183448007891e-10, 3.215598326031168e-10, 3.205870326198977e-10, 
    3.196048055665371e-10, 3.1860409470372325e-10, 3.175762596128989e-10, 
    3.1651396429763645e-10, 3.1541198937676741e-10, 3.1426790280547176e-10, 
    3.1308250469694063e-10, 3.1186001780779863e-10, 3.1060797124002959e-10, 
    3.0933681504101096e-10, 3.0805926802784144e-10, 3.067894811075316e-10, 
    3.0554206224962928e-10, 3.043310649650309e-10, 3.0316898874777811e-10, 
    3.020659040746688e-10, 3.0102872468573041e-10, 3.0006071299773367e-10, 
    2.9916121358497719e-10, 2.9832566499842052e-10, 2.975458350005988e-10, 
    2.968103118569507e-10, 2.961051641659116e-10, 2.9541474831944872e-10, 
    2.9472258451986258e-10, 2.9401225685275105e-10, 2.9326824828755345e-10, 
    2.9247669506686816e-10, 2.9162596832810264e-10, 2.9070710772386491e-10, 
    2.8971405230781553e-10, 2.8864370399868578e-10, 2.8749581730925894e-10, 
    2.8627278421175957e-10, 2.849792949923173e-10, 2.8362198138647111e-10, 
    2.8220900086627373e-10, 2.807496531175264e-10, 2.7925400037026768e-10, 
    2.7773252553723443e-10, 2.7619579368253643e-10, 2.7465416368737337e-10, 
    2.7311746870586294e-10, 2.7159474299326767e-10, 2.7009391967342298e-10, 
    2.6862158055840265e-10, 2.6718270738943999e-10, 2.6578052979580423e-10, 
    2.6441643700634771e-10, 2.6309003833104177e-10, 2.6179932950350074e-10, 
    2.6054103902760824e-10, 2.5931108365824267e-10, 2.581051527002348e-10, 
    2.5691932975383606e-10, 2.5575073423514035e-10, 2.5459806344930187e-10, 
    2.534620198234133e-10, 2.5234549807845119e-10, 2.5125355718922092e-10, 
    2.501930999031296e-10, 2.491723254201925e-10, 2.4819994557571563e-10, 
    2.4728429849587879e-10, 2.4643238598746668e-10, 2.4564899944860385e-10, 
    2.4493597936228207e-10, 2.4429174595901196e-10, 2.4371110597087588e-10, 
    2.4318543023827095e-10, 2.4270311564286634e-10, 2.4225036396142799e-10, 
    2.4181213434167679e-10, 2.413732279544608e-10, 2.4091933449093844e-10, 
    2.4043801484098647e-10, 2.399194363728667e-10, 2.3935688780480657e-10, 
    2.3874695460570188e-10, 2.3808943446819433e-10, 2.3738694038828722e-10, 
    2.3664433529157997e-10, 2.3586799418839359e-10, 2.350650520641793e-10, 
    2.3424263968436192e-10, 2.3340726404813281e-10, 2.3256429849263823e-10, 
    2.317176983224941e-10, 2.3086985908691637e-10, 2.3002169273493751e-10, 
    2.291727985994788e-10, 2.28321771331234e-10, 2.2746652394780077e-10, 
    2.2660464556401164e-10, 2.2573369232218307e-10, 2.248514609038322e-10, 
    2.2395614408126175e-10, 2.2304645980877533e-10, 2.221216886833628e-10, 
    2.2118169747348966e-10, 2.202269078193322e-10, 2.1925831047428887e-10, 
    2.1827744351353766e-10, 2.1728644145302375e-10, 2.1628806231794852e-10, 
    2.1528576301123614e-10, 2.142837326672648e-10, 2.1328693542591061e-10, 
    2.1230105758786562e-10, 2.1133243632713871e-10, 2.1038785522768112e-10, 
    2.0947430719515779e-10, 2.0859864628358123e-10, 2.0776723856643968e-10, 
    2.0698555216051873e-10, 2.0625783210379334e-10, 2.0558678996446402e-10, 
    2.0497344986669253e-10, 2.0441707515078316e-10, 2.039152755746723e-10, 
    2.0346419294786973e-10, 2.0305884230053533e-10, 2.0269345023431474e-10, 
    2.0236187122387634e-10, 2.0205791809950528e-10, 2.0177567032180076e-10, 
    2.0150964196558722e-10, 2.0125488692075668e-10, 2.0100697560301992e-10, 
    2.0076193639833065e-10, 2.00516127694871e-10, 2.0026615897599132e-10, 
    2.0000880515208811e-10, 1.9974103310719299e-10, 1.9946006108275762e-10, 
    1.9916352207745344e-10, 1.9884962304355549e-10, 1.9851735766385106e-10, 
    1.9816662500654435e-10, 1.9779831952930163e-10, 1.9741426645408006e-10, 
    1.9701707715227893e-10, 1.9660982884657656e-10, 1.9619570256171219e-10, 
    1.9577752507351051e-10, 1.9535735058278847e-10, 1.9493607186220449e-10, 
    1.9451320087623911e-10, 1.9408677162937162e-10, 1.9365349938477889e-10, 
    1.932090978950343e-10, 1.9274883150462762e-10, 1.922681544402527e-10, 
    1.91763471060013e-10, 1.9123284047261492e-10, 1.9067662705494855e-10, 
    1.9009793299940139e-10, 1.8950283364609084e-10, 1.8890028942334847e-10, 
    1.8830181054174344e-10, 1.877207967899948e-10, 1.8717168857351188e-10, 
    1.8666891853854046e-10, 1.8622582310977104e-10, 1.8585351610329981e-10, 
    1.8555991755731883e-10, 1.8534892810306152e-10, 1.8521989437209229e-10, 
    1.8516733438398067e-10, 1.8518102930209548e-10, 1.8524638949548849e-10, 
    1.8534514829595804e-10, 1.8545627106769478e-10, 1.8555707058376315e-10, 
    1.8562438552008362e-10, 1.8563581880619705e-10, 1.8557088268697657e-10, 
    1.854120570253938e-10, 1.8514560837400669e-10, 1.8476223552278331e-10, 
    1.8425742663604993e-10, 1.8363159916602369e-10, 1.8288996233827178e-10, 
    1.8204220209813068e-10, 1.8110194488047665e-10, 1.800861138568874e-10, 
    1.79014137522835e-10, 1.7790712034381455e-10, 1.7678694350156615e-10, 
    1.7567539138068332e-10, 1.7459326001624232e-10, 1.735595622015459e-10, 
    1.7259077331880611e-10, 1.7170023102449907e-10, 1.708976398190552e-10, 
    1.7018879032014963e-10, 1.6957542026910407e-10, 1.6905532260924958e-10, 
    1.6862261397942655e-10, 1.6826822319837848e-10, 1.6798049026027466e-10, 
    1.6774591952759616e-10, 1.6754996960867419e-10, 1.673778964787551e-10, 
    1.6721551397626659e-10, 1.6704993209429964e-10, 1.6687015393243642e-10, 
    1.6666756908674614e-10, 1.6643626864756487e-10, 1.6617324876004174e-10, 
    1.6587843456224734e-10, 1.6555458807325245e-10, 1.6520707064387948e-10, 
    1.6484351314875396e-10, 1.6447335092162761e-10, 1.6410731950178622e-10, 
    1.6375685068436169e-10, 1.6343346205400749e-10, 1.6314809944061623e-10, 
    1.6291053331338932e-10, 1.6272875673777771e-10, 1.6260850291349983e-10, 
    1.6255282296808981e-10, 1.6256183220940426e-10, 1.6263256663622194e-10, 
    1.627590328838925e-10, 1.629323815951321e-10, 1.6314126835325924e-10, 
    1.6337232447469375e-10, 1.6361077211985157e-10, 1.6384108178406229e-10, 
    1.6404771130712474e-10, 1.6421582819644779e-10, 1.6433201361386475e-10, 
    1.6438487238602133e-10, 1.6436556149761282e-10, 1.6426815224297855e-10, 
    1.6408986416803551e-10, 1.6383109335431948e-10, 1.6349530712217441e-10, 
    1.6308872357626349e-10, 1.6261988602103453e-10, 1.6209907696885088e-10, 
    1.6153767282440593e-10, 1.6094743311874869e-10, 1.6033981166843978e-10, 
    1.597252995219699e-10, 1.5911289613814567e-10, 1.58509679218522e-10, 
    1.5792057938848963e-10, 1.5734831345415949e-10, 1.5679351938001531e-10, 
    1.5625503064172144e-10, 1.5573031407384994e-10, 1.5521597134209764e-10, 
    1.5470829374912621e-10, 1.5420378402307967e-10, 1.5369962975056679e-10, 
    1.5319402576267901e-10, 1.5268638770904186e-10, 1.5217738870102314e-10, 
    1.5166885842989748e-10, 1.511635277490647e-10, 1.5066470129211539e-10, 
    1.5017585671630111e-10, 1.4970025963604542e-10, 1.4924059778353933e-10, 
    1.487987263854475e-10, 1.4837549633576749e-10, 1.4797073727881266e-10, 
    1.4758334260497327e-10, 1.4721147922514681e-10, 1.4685287003262349e-10, 
    1.465051297125577e-10, 1.4616607459286823e-10, 1.4583402043952497e-10, 
    1.4550797754403419e-10, 1.4518776485679406e-10, 1.4487399201844596e-10, 
    1.4456795628595024e-10, 1.4427142211433804e-10, 1.4398636298299837e-10, 
    1.4371466595794193e-10, 1.4345786805079432e-10, 1.4321691144855642e-10, 
    1.4299200489235865e-10, 1.4278256390123495e-10, 1.4258726073379308e-10, 
    1.424041411766644e-10, 1.4223083604284299e-10, 1.4206480130309386e-10, 
    1.4190358848229621e-10, 1.4174508108919315e-10, 1.4158771479484706e-10, 
    1.4143062845514189e-10, 1.4127375671190433e-10, 1.4111783268717126e-10, 
    1.4096433958733554e-10, 1.4081537247746905e-10, 1.4067345539680126e-10, 
    1.4054130089159851e-10, 1.404215445566703e-10, 1.4031643106609486e-10, 
    1.4022753590717631e-10, 1.401554558987634e-10, 1.4009956981125753e-10, 
    1.4005783090412062e-10, 1.4002664593570102e-10, 1.4000083215203161e-10, 
    1.3997369588539314e-10, 1.3993718643951691e-10, 1.3988217660024622e-10, 
    1.3979880700249414e-10, 1.3967691208716258e-10, 1.3950645101583505e-10, 
    1.3927796495319418e-10, 1.3898299121204485e-10, 1.3861442532540819e-10, 
    1.3816679493965399e-10, 1.3763645734739615e-10, 1.370216923187708e-10, 
    1.3632271324264987e-10, 1.3554159954720655e-10, 1.3468217763166759e-10, 
    1.3374985109076756e-10, 1.3275142901089107e-10, 1.3169492602754354e-10, 
    1.3058938523856187e-10, 1.2944470414745554e-10, 1.2827147778946348e-10, 
    1.2708084215127564e-10, 1.258843348824145e-10, 1.2469373557314339e-10, 
    1.2352090476581413e-10, 1.2237759826268086e-10, 1.2127526948022717e-10, 
    1.2022482090412125e-10, 1.1923635725545114e-10, 1.1831891739313317e-10, 
    1.1748020123298834e-10, 1.1672630701761994e-10, 1.1606151069236364e-10, 
    1.1548809797172073e-10, 1.1500626628107672e-10, 1.1461412081427621e-10, 
    1.143077723093466e-10, 1.1408150801255178e-10, 1.1392806396587821e-10, 
    1.1383895243271941e-10, 1.13804817559962e-10, 1.1381578873891857e-10, 
    1.1386181694085773e-10, 1.139329446509296e-10, 1.1401952716512888e-10, 
    1.1411238037934472e-10, 1.1420288816434822e-10, 1.1428305793328857e-10, 
    1.1434558636676705e-10, 1.1438392754740261e-10, 1.1439239226852986e-10, 
    1.1436628422101679e-10, 1.1430206612193876e-10, 1.1419752492422848e-10, 
    1.1405193799555886e-10, 1.1386617091828242e-10, 1.1364270979363259e-10, 
    1.1338558481939136e-10, 1.1310018672435632e-10, 1.1279296818589332e-10, 
    1.1247106274076116e-10, 1.1214185028152036e-10, 1.1181251066807711e-10, 
    1.114896059336814e-10, 1.1117873720039948e-10, 1.1088431063345163e-10, 
    1.1060942995920052e-10, 1.1035590775800668e-10, 1.101243967121759e-10, 
    1.099146076948148e-10, 1.097255818199658e-10, 1.0955597458756855e-10, 
    1.0940430609161392e-10, 1.0926918290194259e-10, 1.091494263827212e-10, 
    1.0904412086713268e-10, 1.0895259559481044e-10, 1.0887433750199482e-10, 
    1.0880886686863763e-10, 1.0875559380174168e-10, 1.0871367789232007e-10, 
    1.0868192242739855e-10, 1.0865869339623101e-10, 1.0864189028402772e-10, 
    1.0862894175250375e-10, 1.0861684724864061e-10, 1.0860221902119688e-10, 
    1.0858134472109628e-10, 1.0855024723059407e-10, 1.0850473088230225e-10, 
    1.0844044027618484e-10, 1.0835292454666409e-10, 1.0823772306789687e-10, 
    1.0809048809639902e-10, 1.0790715700223185e-10, 1.0768417762895599e-10, 
    1.0741877382133873e-10, 1.0710925623144151e-10, 1.0675532737552401e-10, 
    1.0635836361919944e-10, 1.0592163545145759e-10, 1.0545041274176876e-10, 
    1.0495195073453411e-10, 1.0443531606621882e-10, 1.0391106619411762e-10, 
    1.033907798631136e-10, 1.0288648737215377e-10, 1.0241002861250729e-10, 
    1.0197239399880463e-10, 1.0158311164083504e-10, 1.0124972008667164e-10, 
    1.0097735348244991e-10, 1.0076849828790489e-10, 1.0062290635141502e-10, 
    1.0053767706231504e-10, 1.0050747845006892e-10, 1.0052490142809413e-10, 
    1.0058091657779366e-10, 1.0066539423266259e-10, 1.0076767164565162e-10, 
    1.0087713358470322e-10, 1.0098379802271208e-10, 1.0107886407201129e-10, 
    1.0115521074945534e-10, 1.012078194125329e-10, 1.0123408405876691e-10, 
    1.0123398330292207e-10, 1.0121007811874495e-10, 1.0116732214793329e-10, 
    1.0111266486757214e-10, 1.0105446460055896e-10, 1.0100172309315568e-10, 
    1.0096321213104989e-10, 1.009465502659451e-10, 1.0095731431517864e-10, 
    1.0099828771838672e-10, 1.0106892537920629e-10, 1.0116509921838396e-10, 
    1.0127919603346618e-10, 1.0140055090036382e-10, 1.015162177420654e-10, 
    1.0161199364931485e-10, 1.0167363031378087e-10, 1.0168808720691362e-10, 
    1.0164473453370328e-10, 1.0153636451995422e-10, 1.0135991693927544e-10, 
    1.0111685178760792e-10, 1.0081312623871774e-10, 1.0045878356238546e-10, 
    1.0006719922411747e-10, 9.9654058272611048e-11, 9.9236173837116324e-11, 
    9.8830234739651012e-11, 9.8451618755839332e-11, 9.8113365723326259e-11, 
    9.7825378148949192e-11, 9.7593900934726744e-11, 9.7421312703788238e-11, 
    9.7306220079989852e-11, 9.7243796357985661e-11, 9.7226342395494378e-11, 
    9.7243987418270287e-11, 9.7285444150521708e-11, 9.7338789255958325e-11, 
    9.7392176414082545e-11, 9.7434451705120378e-11, 9.7455651591669441e-11, 
    9.7447363829584974e-11, 9.7402949083782394e-11, 9.731764947293519e-11, 
    9.7188609476492578e-11, 9.7014815738428091e-11, 9.6796972769746504e-11, 
    9.6537352096642051e-11, 9.623959513714811e-11, 9.5908485950478622e-11, 
    9.55496821300709e-11, 9.5169398306815746e-11, 9.4774049905779887e-11, 
    9.4369857260951541e-11, 9.3962418508938308e-11, 9.3556291422574699e-11, 
    9.3154605804143954e-11, 9.2758748868578895e-11, 9.2368155038184158e-11, 
    9.1980234809741469e-11, 9.1590470971996897e-11, 9.1192672373502124e-11, 
    9.0779382134052128e-11, 9.0342417482687134e-11, 8.9873494919755858e-11, 
    8.9364894779428222e-11, 8.8810104758722237e-11, 8.8204398055938925e-11, 
    8.7545301006395495e-11, 8.6832912627035552e-11, 8.6070051423480792e-11, 
    8.5262251156567724e-11, 8.4417568225191336e-11, 8.3546277454640683e-11, 
    8.2660440376336454e-11, 8.1773401165866151e-11, 8.0899251338566886e-11, 
    8.0052278175365102e-11, 7.9246425898533841e-11, 7.8494805765535216e-11, 
    7.7809252064804943e-11, 7.7199938459809196e-11, 7.6675047422513806e-11, 
    7.6240520500287057e-11, 7.5899846743136147e-11, 7.5653931472250136e-11, 
    7.5501039409599027e-11, 7.5436805512365828e-11, 7.5454329151143559e-11, 
    7.5544370677769105e-11, 7.5695630025956907e-11, 7.5895124229430777e-11, 
    7.6128647661782257e-11, 7.6381295187011155e-11, 7.6638033417024878e-11, 
    7.6884282645301109e-11, 7.7106484341268553e-11, 7.7292626301558776e-11, 
    7.7432682859370251e-11, 7.751896568011374e-11, 7.7546344163196378e-11, 
    7.7512344833110329e-11, 7.7417118596553306e-11, 7.7263270802115218e-11, 
    7.7055578424392894e-11, 7.6800609132744709e-11, 7.6506256911017862e-11, 
    7.6181234539810769e-11, 7.583454461556872e-11, 7.5474966075280709e-11, 
    7.5110589741531253e-11, 7.4748434148828211e-11, 7.4394161326936848e-11, 
    7.4051918249990177e-11, 7.3724307443010746e-11, 7.341248488781124e-11, 
    7.3116379254740221e-11, 7.2835003308514349e-11, 7.2566821791077896e-11, 
    7.2310152389750009e-11, 7.2063555863886427e-11, 7.1826179269670441e-11, 
    7.1598005565463428e-11, 7.1380020802095212e-11, 7.1174247073985361e-11, 
    7.0983673394177221e-11, 7.0812061186453767e-11, 7.0663675605608989e-11, 
    7.0542950259702859e-11, 7.0454124885630153e-11, 7.0400889766220477e-11, 
    7.0386076164638603e-11, 7.0411408811856346e-11, 7.0477354255089598e-11, 
    7.0583063214919728e-11, 7.0726413518481204e-11, 7.0904144212582726e-11, 
    7.1112057891230699e-11, 7.1345257021018336e-11, 7.1598416435706176e-11, 
    7.1866022430505411e-11, 7.214259798412008e-11, 7.2422866296440988e-11, 
    7.2701859726537391e-11, 7.2974976834008237e-11, 7.3237991114222444e-11, 
    7.3487012864854118e-11, 7.3718462021201268e-11, 7.3929018856767841e-11, 
    7.4115614514465279e-11, 7.4275454206343746e-11, 7.4406081775559254e-11, 
    7.4505485382151169e-11, 7.4572248370158451e-11, 7.4605704504312687e-11, 
    7.4606115781637303e-11, 7.4574798584598458e-11, 7.4514231885415513e-11, 
    7.4428067794129885e-11, 7.4321073874369458e-11, 7.4198977031063137e-11, 
    7.4068216979018468e-11, 7.39356202713217e-11, 7.3808031013253174e-11, 
    7.3691903498020709e-11, 7.3592925664455901e-11, 7.3515665846160162e-11, 
    7.3463317593855108e-11, 7.3437512490710777e-11, 7.3438246733796163e-11, 
    7.3463902848894544e-11, 7.3511364958932841e-11, 7.3576170788381117e-11, 
    7.3652737398785036e-11, 7.3734579046646551e-11, 7.3814542665737058e-11, 
    7.3885024083698335e-11, 7.3938183992318611e-11, 7.396615598056611e-11, 
    7.3961274526882819e-11, 7.3916316774708392e-11, 7.3824800635674008e-11, 
    7.3681299921343213e-11, 7.34818165918951e-11, 7.3224144853535538e-11, 
    7.2908235721490937e-11, 7.2536496325778036e-11, 7.2114000917132671e-11, 
    7.1648544627727365e-11, 7.1150551028145049e-11, 7.0632768497090119e-11, 
    7.0109800302890565e-11, 6.9597438192238162e-11, 6.9111893148210146e-11, 
    6.866891534747599e-11, 6.8282919653611644e-11, 6.7966149868397193e-11, 
    6.772797098266349e-11, 6.7574302161638996e-11, 6.7507288729005227e-11, 
    6.7525185094661041e-11, 6.7622489324388212e-11, 6.7790281400428486e-11, 
    6.8016768509210844e-11, 6.8287968843573931e-11, 6.8588502106588239e-11, 
    6.8902412047708093e-11, 6.921400430154277e-11, 6.9508592171496115e-11, 
    6.9773175737962811e-11, 6.999696193032705e-11, 7.0171743683601749e-11, 
    7.0292107826849694e-11, 7.0355488478332824e-11, 7.0362047908602251e-11, 
    7.0314457810491541e-11, 7.0217569475902859e-11, 7.007803072940173e-11, 
    6.9903877459343974e-11, 6.9704142185166799e-11, 6.9488489513981234e-11, 
    6.9266919011183904e-11, 6.9049511579305517e-11, 6.8846251572230714e-11, 
    6.8666857320974055e-11, 6.852066723814379e-11, 6.8416486159163465e-11, 
    6.8362440587131232e-11, 6.83657819507929e-11, 6.8432668020434765e-11, 
    6.8567907886400517e-11, 6.8774706046808356e-11, 6.9054415193845905e-11, 
    6.9406338891060865e-11, 6.9827587290529731e-11, 7.0313043013824766e-11, 
    7.0855394328571008e-11, 7.1445298071195018e-11, 7.2071636063178275e-11, 
    7.2721866442036272e-11, 7.3382440708008556e-11, 7.4039304533234688e-11, 
    7.467842202799505e-11, 7.5286340326962576e-11, 7.5850740832631412e-11, 
    7.636098261368401e-11, 7.6808572928447301e-11, 7.7187570183000217e-11, 
    7.7494849375128304e-11, 7.7730237126387524e-11, 7.7896441747363801e-11, 
    7.7998821325412969e-11, 7.8044938942330865e-11, 7.8043964363456049e-11, 
    7.8005934262309961e-11, 7.794095126124414e-11, 7.7858370010476274e-11, 
    7.7766077822049337e-11, 7.7669903660089202e-11, 7.7573262857771761e-11, 
    7.7477046559629846e-11, 7.737979166398351e-11, 7.7278104777492372e-11, 
    7.7167305804490653e-11, 7.7042209668308648e-11, 7.6897971508973898e-11, 
    7.6730862840135265e-11, 7.6538929434857453e-11, 7.6322409870901195e-11, 
    7.6083888446318372e-11, 7.5828135879432411e-11, 7.5561681367957133e-11, 
    7.5292159214742632e-11, 7.5027504187406794e-11, 7.4775103963211081e-11, 
    7.4541024992721172e-11, 7.4329378558198221e-11, 7.4141942816217457e-11, 
    7.3978030921116522e-11, 7.3834660106490101e-11, 7.3706938793823158e-11, 
    7.3588648604116157e-11, 7.3472891573094808e-11, 7.3352760492672108e-11, 
    7.3221897975634895e-11, 7.3074919470780309e-11, 7.2907649969402625e-11, 
    7.2717169540610516e-11, 7.2501694073696433e-11, 7.2260354123950367e-11, 
    7.1992918870744757e-11, 7.1699546748731351e-11, 7.1380587846169848e-11, 
    7.1036510489965e-11, 7.0667933381249085e-11, 7.0275768201711329e-11, 
    6.9861428545210189e-11, 6.9427072602257411e-11, 6.8975811076364405e-11, 
    6.8511856002295894e-11, 6.8040547095363589e-11, 6.7568259230532576e-11, 
    6.7102180000190909e-11, 6.6649979591076568e-11, 6.6219385919247384e-11, 
    6.5817737777773041e-11, 6.5451543700434541e-11, 6.5126094135962391e-11, 
    6.4845155994930374e-11, 6.4610794939565316e-11, 6.4423325962880932e-11, 
    6.4281391428941413e-11, 6.4182149802750064e-11, 6.4121565738183216e-11, 
    6.4094744529351668e-11, 6.4096300052986489e-11, 6.4120706445046758e-11, 
    6.4162605701060229e-11, 6.4217043448611083e-11, 6.4279621401634552e-11, 
    6.4346562018637331e-11, 6.4414678985934046e-11, 6.4481276313926345e-11, 
    6.4543990139244593e-11, 6.4600599907619344e-11, 6.4648837350884004e-11, 
    6.4686213285833336e-11, 6.4709905054343872e-11, 6.4716695777188164e-11, 
    6.4703005271146473e-11, 6.4665003130404932e-11, 6.4598805242745382e-11, 
    6.4500731276044671e-11, 6.4367620685579262e-11, 6.4197160568486e-11, 
    6.3988207493600988e-11, 6.3741064395686226e-11, 6.3457686459232738e-11, 
    6.314178205741172e-11, 6.2798790259172299e-11, 6.2435738038518184e-11, 
    6.2060959848528342e-11, 6.1683713521156464e-11, 6.1313704487899339e-11, 
    6.0960569976721504e-11, 6.0633354950537501e-11, 6.0340027834963456e-11, 
    6.0087081653641659e-11, 5.9879256357689274e-11, 5.9719398756238117e-11, 
    5.9608477491191643e-11, 5.9545741151613115e-11, 5.9529007185866646e-11, 
    5.9555038260955725e-11, 5.9619973825026661e-11, 5.9719766190425012e-11, 
    5.9850583446810577e-11, 6.0009132105263125e-11, 6.0192868589827652e-11, 
    6.0400089465000783e-11, 6.0629875437075231e-11, 6.0881914439294705e-11, 
    6.1156215413056676e-11, 6.1452735150282355e-11, 6.1770971033383971e-11, 
    6.2109554879565787e-11, 6.2465900271637341e-11, 6.2835940756295986e-11, 
    6.321398711767575e-11, 6.359274149219915e-11, 6.3963468097537742e-11, 
    6.4316309441646243e-11, 6.4640730595140997e-11, 6.4926049629051265e-11, 
    6.5162021511475288e-11, 6.5339403607184886e-11, 6.5450476985561822e-11, 
    6.5489460398505165e-11, 6.5452806227289117e-11, 6.5339336449834461e-11, 
    6.515023669538724e-11, 6.4888901735842619e-11, 6.4560670075427854e-11, 
    6.4172456540482661e-11, 6.3732342898422774e-11, 6.3249150385784334e-11, 
    6.2732030523073678e-11, 6.2190108450787861e-11, 6.163220098193388e-11, 
    6.1066625948732075e-11, 6.0501094699004578e-11, 5.9942689475208706e-11, 
    5.9397907410440309e-11, 5.8872728375821482e-11, 5.8372701458040927e-11, 
    5.7902987112876175e-11, 5.7468353256007807e-11, 5.707309179697821e-11, 
    5.6720860071304175e-11, 5.64144539715619e-11, 5.6155548223438407e-11, 
    5.5944436325178022e-11, 5.5779829013100471e-11, 5.5658753359909298e-11, 
    5.557659469512627e-11, 5.5527308002534744e-11, 5.5503801982127923e-11, 
    5.5498461742059927e-11, 5.5503782067720289e-11, 5.5513029840014618e-11, 
    5.5520869722740333e-11, 5.5523876604801584e-11,
  // Sqw-total(9, 0-1999)
    0.018573087278200315, 0.018570966064277734, 0.018564665303538626, 
    0.01855436884812562, 0.018540367546982441, 0.018523037251051252, 
    0.018502810629165971, 0.018480145140671565, 0.018455489824965796, 
    0.01842925364899067, 0.018401777987213676, 0.018373315402899996, 
    0.018344016286367761, 0.018313924140633781, 0.018282979462465578, 
    0.01825103133579736, 0.018217855127227442, 0.018183174135211387, 
    0.018146682762059576, 0.018108068788056153, 0.01806703263036559, 
    0.018023302026942651, 0.017976641322045784, 0.017926855342304815, 
    0.017873788624026995, 0.017817321370386965, 0.017757363889293054, 
    0.01769385133356564, 0.017626740325911869, 0.017556008543114756, 
    0.017481657642352644, 0.017403719154328881, 0.017322262271735136, 
    0.01723740194668762, 0.017149305466164239, 0.017058195743453942, 
    0.016964349936374364, 0.016868092618600082, 0.016769783488143935, 
    0.016669800374541584, 0.016568518981494359, 0.016466291273608474, 
    0.016363424620774555, 0.016260163733964213, 0.016156677089810795, 
    0.016053049013671213, 0.015949277960250089, 0.015845280891573839, 
    0.015740903088152774, 0.015635932302096995, 0.015530115903176161, 
    0.015423179583278466, 0.015314846249711909, 0.015204853915194889, 
    0.015092971637142511, 0.014979012827539082, 0.014862845511759608, 
    0.014744399335955912, 0.014623669295847715, 0.014500716283467432, 
    0.014375664629387146, 0.014248696868498887, 0.014120045992599759, 
    0.013989985488199852, 0.013858817506356862, 0.013726859581707317, 
    0.013594430412307042, 0.013461835324193533, 0.013329352159622943, 
    0.013197218422837741, 0.01306562056442615, 0.012934686257577542, 
    0.012804480395905661, 0.012675005314507154, 0.012546205411951818, 
    0.012417975958048869, 0.012290175454281238, 0.012162640525635985, 
    0.012035202021551105, 0.011907700839709285, 0.011780001992282872, 
    0.011652005618805718, 0.01152365399492305, 0.011394934048433267, 
    0.011265875411002877, 0.0111365445344679, 0.011007035816102491, 
    0.01087746095283418, 0.0107479378478557, 0.010618580319473991, 
    0.010489489633646877, 0.010360748543307666, 0.010232418128133488, 
    0.010104537350205814, 0.009977124929090371, 0.0098501829330680107, 
    0.0097237013986192083, 0.009597663321766859, 0.0094720494864565935, 
    0.0093468427674121644, 0.0092220317239914817, 0.0090976134483953426, 
    0.0089735957195500749, 0.0088499985337201648, 0.008726855043055412, 
    0.0086042118574507203, 0.008482128585589695, 0.0083606764408986275, 
    0.0082399357432123184, 0.0081199922197838781, 0.0080009321459346763, 
    0.0078828365463289377, 0.007765774870774473, 0.0076497987263209151, 
    0.007534936354920199, 0.0074211885666662708, 0.0073085267602354103, 
    0.0071968934884155599, 0.0070862057767358336, 0.0069763611082896406, 
    0.006867245685663618, 0.0067587443100102854, 0.006650751011643103, 
    0.0065431794511667798, 0.0064359720987867105, 0.0063291072936208894, 
    0.0062226034745627608, 0.0061165201396485127, 0.0060109554045323201, 
    0.0059060403602920692, 0.005801930742177489, 0.0056987966811546196, 
    0.0055968114907932803, 0.005496140522567341, 0.0053969310929308503, 
    0.0052993043480376563, 0.0052033497021495212, 0.0051091221909021151, 
    0.0050166427566862406, 0.0049259011706030819, 0.0048368610324811302, 
    0.0047494661090079189, 0.0046636471901738792, 0.004579328671467626, 
    0.0044964341940269296, 0.0044148908744158569, 0.0043346318976708589, 
    0.0042555974953948916, 0.0041777345500933552, 0.004100995229298487, 
    0.0040253351402631289, 0.0039507115022745197, 0.0038770817652356991, 
    0.0038044029766558804, 0.0037326320381811271, 0.0036617268239380421, 
    0.0035916479818570361, 0.0035223611267540381, 0.0034538390739675389, 
    0.0033860637598170295, 0.0033190275464202003, 0.0032527337023485806, 
    0.0031871959707427842, 0.0031224372638037757, 0.0030584876382802172, 
    0.0029953817948900076, 0.0029331563946871043, 0.0028718474924656137, 
    0.0028114883529440854, 0.0027521078469044799, 0.0026937295331413303, 
    0.0026363714318906597, 0.002580046400642222, 0.0025247629466722751, 
    0.0024705262619587826, 0.0024173392508793881, 0.0023652033400785224, 
    0.0023141189093587857, 0.0022640852546614693, 0.0022151000785291803, 
    0.0021671585877913045, 0.0021202523505985172, 0.0020743681150434323, 
    0.0020294868121789396, 0.0019855829540425013, 0.001942624593585173, 
    0.0019005739438255956, 0.0018593886673990438, 0.0018190237566431335, 
    0.0017794338409545089, 0.0017405756939195126, 0.0017024106766619, 
    0.0016649068511150659, 0.0016280405281127732, 0.0015917970762591048, 
    0.0015561709004147965, 0.0015211645923857797, 0.0014867873488006238, 
    0.0014530528304388341, 0.0014199766937292963, 0.0013875740524512186, 
    0.0013558571236523276, 0.0013248332785223398, 0.001294503662271162, 
    0.0012648624755409305, 0.0012358969334801825, 0.0012075878471395306, 
    0.0011799107136223463, 0.0011528371621930102, 0.0011263365859378585, 
    0.0011003777920375285, 0.0010749305249622217, 0.0010499667507367328, 
    0.0010254616307337097, 0.0010013941542515884, 0.00097774743541997476, 
    0.00095450870831311559, 0.00093166907290664284, 0.00090922305374280385, 
    0.00088716803426712898, 0.00086550362495851961, 0.00084423101504059049, 
    0.00082335234793604712, 0.00080287015133821867, 0.00078278684472394753, 
    0.00076310434052511561, 0.00074382374968019781, 0.00072494519729126574, 
    0.00070646774897816411, 0.00068838944282121749, 0.00067070741543394277, 
    0.00065341810403132274, 0.00063651750003265186, 0.00062000142467290244, 
    0.00060386579425358486, 0.00058810684286458479, 0.00057272127413640682, 
    0.00055770632085725259, 0.00054305970158317559, 0.00052877947563917068, 
    0.0005148638106957351, 0.0005013106887390321, 0.00048811758509016137, 
    0.0004752811598267801, 0.00046279700069957021, 0.00045065945128870189, 
    0.00043886154831614181, 0.00042739507899093923, 0.00041625075476174611, 
    0.0004054184838420245, 0.00039488771321664212, 0.00038464780301981899, 
    0.00037468839308539239, 0.00036499972331367433, 0.00035557287579100272, 
    0.00034639991630072654, 0.00033747392457410757, 0.00032878891482269692, 
    0.00032033965933862645, 0.0003121214370969565, 0.00030412973557428501, 
    0.0002963599370639605, 0.00028880702065509588, 0.00028146530810039503, 
    0.0002743282765853016, 0.00026738845460875068, 0.00026063740950606125, 
    0.00025406582727956423, 0.00024766367797462795, 0.00024142045337937029, 
    0.00023532545874739515, 0.00022936813682641403, 0.00022353840085405173, 
    0.00021782695334263518, 0.00021222556926197788, 0.000206727325379495, 
    0.00020132676169109593, 0.00019601996571328475, 0.00019080457555956294, 
    0.00018567970289511517, 0.00018064578180640052, 0.00017570435413631004, 
    0.00017085780573425794, 0.00016610907116292698, 0.00016146132647195917, 
    0.00015691769046868257, 0.00015248095428027658, 0.00014815335678693465, 
    0.00014393641972301329, 0.00013983085109712148, 0.00013583651948006643, 
    0.00013195249524864484, 0.00012817714876597319, 0.00012450829046241558, 
    0.00012094333449163769, 0.00011747946650959352, 0.00011411379730503739, 
    0.00011084348732681047, 0.00010766583212764952, 0.00010457830467015598, 
    0.00010157855648329753, 9.8664384990270298e-05, 9.583367824761904e-05, 
    9.3084350372802201e-05, 9.0414280912843014e-05, 8.7821269453110579e-05, 
    8.5303013286966938e-05, 8.2857111574269324e-05, 8.048109481749819e-05, 
    7.8172474379406304e-05, 7.5928803737401295e-05, 7.3747741606405663e-05, 
    7.1627107104937682e-05, 6.9564918683289828e-05, 6.7559411250737154e-05, 
    6.5609029352971959e-05, 6.3712397809335917e-05, 6.1868274391159314e-05, 
    6.0075491469384507e-05, 5.8332894801035591e-05, 5.6639287658093388e-05, 
    5.4993387412016665e-05, 5.3393799704464503e-05, 5.1839012799991687e-05, 
    5.0327412012451e-05, 4.8857311598173875e-05, 4.7426999524464928e-05, 
    4.6034789266418762e-05, 4.46790723532746e-05, 4.3358365759639075e-05, 
    4.2071349292494597e-05, 4.0816889665971824e-05, 3.9594049739837785e-05, 
    3.8402083178347764e-05, 3.7240416340001587e-05, 3.6108620367815001e-05, 
    3.500637711266754e-05, 3.3933442667492778e-05, 3.2889611964168572e-05, 
    3.1874687196250886e-05, 3.0888451920041651e-05, 2.9930651711233681e-05, 
    2.9000981356168149e-05, 2.8099077849748752e-05, 2.7224518022790274e-05, 
    2.6376819451080437e-05, 2.5555443379001772e-05, 2.4759798662617118e-05, 
    2.3989246116103629e-05, 2.324310304528685e-05, 2.2520648091661586e-05, 
    2.1821126733027464e-05, 2.1143757859534081e-05, 2.0487741766284489e-05, 
    1.9852269698845111e-05, 1.923653480326369e-05, 1.8639744023383636e-05, 
    1.806113021671335e-05, 1.7499963576633953e-05, 1.6955561391860553e-05, 
    1.6427295258090205e-05, 1.5914595075950098e-05, 1.5416949492823595e-05, 
    1.493390282910663e-05, 1.4465048914390463e-05, 1.4010022591358027e-05, 
    1.356848987560704e-05, 1.3140137858488103e-05, 1.2724665395773869e-05, 
    1.2321775450591612e-05, 1.1931169684086751e-05, 1.1552545557098275e-05, 
    1.1185595868197553e-05, 1.0830010355601264e-05, 1.0485478767101914e-05, 
    1.015169467668265e-05, 9.8283593032042646e-06, 9.5151846582263789e-06, 
    9.2118954957463039e-06, 8.9182297319693335e-06, 8.6339372192436855e-06, 
    8.3587769713709749e-06, 8.0925131254167598e-06, 7.8349100743761937e-06, 
    7.5857273043623531e-06, 7.3447145159805503e-06, 7.1116075994895647e-06, 
    6.8861259708783088e-06, 6.6679716650061651e-06, 6.4568304321822959e-06, 
    6.2523749064997612e-06, 6.0542697240409613e-06, 5.8621782821779694e-06, 
    5.6757706671404613e-06, 5.4947321509230703e-06, 5.3187715857402885e-06, 
    5.1476290118133269e-06, 4.9810818461059503e-06, 4.8189491297022703e-06, 
    4.6610934702681863e-06, 4.5074205057232065e-06, 4.3578759179345416e-06, 
    4.2124402191461776e-06, 4.0711217020369408e-06, 3.9339480705478311e-06, 
    3.8009573452725048e-06, 3.6721886596734998e-06, 3.5476735360001517e-06, 
    3.4274281590489062e-06, 3.3114470642888152e-06, 3.1996985356386899e-06, 
    3.0921218809283792e-06, 2.9886266284384709e-06, 2.8890935749128861e-06, 
    2.7933775169556251e-06, 2.7013114172494831e-06, 2.6127116935849114e-06, 
    2.5273842735513453e-06, 2.4451310298869455e-06, 2.3657562031806665e-06, 
    2.2890724300679274e-06, 2.2149060291140931e-06, 2.1431012520382992e-06, 
    2.0735232846137451e-06, 2.0060598736018916e-06, 1.940621557675894e-06, 
    1.8771405809504532e-06, 1.8155686587019744e-06, 1.7558738355761733e-06, 
    1.6980367215030806e-06, 1.6420464052409927e-06, 1.5878963322754984e-06, 
    1.535580396628857e-06, 1.485089444165117e-06, 1.4364083264613933e-06, 
    1.3895135891968899e-06, 1.3443718326706827e-06, 1.3009387491431496e-06, 
    1.2591588205741213e-06, 1.2189656489779518e-06, 1.1802828836950744e-06, 
    1.1430257011117112e-06, 1.1071027776287402e-06, 1.0724186754512051e-06, 
    1.0388765333765453e-06, 1.0063809263365404e-06, 9.7484073267419875e-07, 
    9.4417183407865897e-07, 9.1429947365745424e-07, 8.8516011618433678e-07, 
    8.5670268955911353e-07, 8.2888913535236263e-07, 8.0169425204283688e-07, 
    7.7510487111838671e-07, 7.4911845576061429e-07, 7.2374124990858659e-07, 
    6.989861279583953e-07, 6.7487030266174337e-07, 6.51413041568051e-07, 
    6.2863352516835676e-07, 6.0654895555369788e-07, 5.8517299789042519e-07, 
    5.6451461010803271e-07, 5.4457729152430221e-07, 5.2535875796462407e-07, 
    5.068510300464714e-07, 4.8904090070260655e-07, 4.7191072871843915e-07, 
    4.5543948615868707e-07, 4.3960397162455376e-07, 4.2438008910100942e-07, 
    4.0974408712722627e-07, 3.9567365586792392e-07, 3.8214879253527588e-07, 
    3.6915236699477159e-07, 3.5667034855952532e-07, 3.4469168787388641e-07, 
    3.3320788143101493e-07, 3.2221227571933788e-07, 3.1169919065807339e-07, 
    3.0166295439753213e-07, 2.9209694386273038e-07, 2.8299271711053688e-07, 
    2.7433930765057184e-07, 2.6612272917691692e-07, 2.5832571599503441e-07, 
    2.5092770181238751e-07, 2.4390502091102391e-07, 2.3723130159140846e-07, 
    2.308780135792338e-07, 2.2481512740734519e-07, 2.1901184463143518e-07, 
    2.1343736064387523e-07, 2.0806162655090053e-07, 2.02856080904545e-07, 
    1.977943263557492e-07, 1.9285272924964505e-07, 1.8801092288333245e-07, 
    1.8325219703501055e-07, 1.7856375868758943e-07, 1.7393685139004435e-07, 
    1.6936672441360022e-07, 1.6485244731816512e-07, 1.6039657149042925e-07, 
    1.5600464682030314e-07, 1.5168460956387463e-07, 1.4744606522737856e-07, 
    1.4329949850835548e-07, 1.3925544930847219e-07, 1.3532369970665568e-07, 
    1.3151251979183898e-07, 1.2782802055526524e-07, 1.2427365803724051e-07, 
    1.2084992522656132e-07, 1.1755425612153633e-07, 1.1438115132364338e-07, 
    1.1132251707605889e-07, 1.0836819217512512e-07, 1.0550662080788834e-07, 
    1.0272561688791584e-07, 1.0001315761314137e-07, 9.7358142680130918e-08, 
    9.475106019118491e-08, 9.2184511086955397e-08, 8.9653558657459537e-08, 
    8.7155887184828389e-08, 8.4691770986484654e-08, 8.2263870785284185e-08, 
    7.987688596801702e-08, 7.7537098711873408e-08, 7.5251848390104461e-08, 
    7.3028973387520372e-08, 7.0876253083327909e-08, 6.8800877467880617e-08, 
    6.6808966211369007e-08, 6.4905154948934373e-08, 6.309226344797424e-08, 
    6.1371058981339338e-08, 5.9740126894368217e-08, 5.819585891838801e-08, 
    5.673256639293829e-08, 5.5342720265348732e-08, 5.4017311828690803e-08, 
    5.2746318741419384e-08, 5.1519250444219481e-08, 5.0325737872684826e-08, 
    4.9156125187623347e-08, 4.8002018342075997e-08, 4.6856746578721026e-08, 
    4.5715699454766593e-08, 4.4576512305416701e-08, 4.3439086723686187e-08, 
    4.2305447195177191e-08, 4.1179449468322288e-08, 4.0066368297621154e-08, 
    3.8972401187815195e-08, 3.790412949181158e-08, 3.6867979201970506e-08, 
    3.5869720692059091e-08, 3.4914041028419379e-08, 3.4004214408276922e-08, 
    3.3141887597780764e-08, 3.2326987771677662e-08, 3.1557751568232086e-08, 
    3.0830865977869706e-08, 3.0141705167061454e-08, 2.9484641834918563e-08, 
    2.8853408248088027e-08, 2.8241480113786534e-08, 2.7642456709290494e-08, 
    2.7050412403820188e-08, 2.6460198560373778e-08, 2.5867679585828097e-08, 
    2.5269893036245353e-08, 2.4665129718403097e-08, 2.4052935848426289e-08, 
    2.3434044337230379e-08, 2.2810246253904604e-08, 2.218421580995242e-08, 
    2.1559303309490915e-08, 2.0939310016558524e-08, 2.0328257839963965e-08, 
    1.9730164860278777e-08, 1.9148836084438371e-08, 1.8587677056625814e-08, 
    1.8049536861910413e-08, 1.7536585944764661e-08, 1.7050233516980136e-08, 
    1.659108814583141e-08, 1.6158963882456895e-08, 1.5752932048030342e-08, 
    1.5371416292121215e-08, 1.5012325149297108e-08, 1.4673213204741275e-08, 
    1.4351458846520973e-08, 1.4044444706158367e-08, 1.3749726014317965e-08, 
    1.3465173151613967e-08, 1.3189077068916119e-08, 1.2920210334062216e-08, 
    1.2657841169782365e-08, 1.2401703050455525e-08, 1.2151926767130443e-08, 
    1.1908945429021043e-08, 1.1673384600891122e-08, 1.1445950122573982e-08, 
    1.1227324570621052e-08, 1.1018080921398505e-08, 1.0818618452261509e-08, 
    1.0629122722991159e-08, 1.0449548275284906e-08, 1.0279620641898943e-08, 
    1.0118852856594641e-08, 9.9665716131017004e-09, 9.8219485830553478e-09, 
    9.6840336830865868e-09, 9.5517881971780026e-09, 9.4241170750838805e-09, 
    9.2999003866406479e-09, 9.1780245875964738e-09, 9.0574140599436739e-09, 
    8.9370632073015476e-09, 8.8160685543613996e-09, 8.6936598116915948e-09, 
    8.5692280175809567e-09, 8.4423485735132788e-09, 8.3127966804184489e-09, 
    8.1805530146942535e-09, 8.0457978259704551e-09, 7.9088926578586885e-09, 
    7.770349779177457e-09, 7.6307908051223657e-09, 7.4908969982306732e-09, 
    7.3513549676603919e-09, 7.2128020732837888e-09, 7.0757763326226176e-09, 
    6.9406753411221061e-09, 6.8077282116842221e-09, 6.6769832645869881e-09, 
    6.5483129191883177e-09, 6.4214354279417308e-09, 6.2959516185977673e-09, 
    6.1713932125771413e-09, 6.0472783741577044e-09, 5.923169358100725e-09, 
    5.7987272535892842e-09, 5.67375904947929e-09, 5.5482533351805374e-09, 
    5.4224019070683059e-09, 5.2966060960170017e-09, 5.1714677468860693e-09, 
    5.0477661197522374e-09, 4.9264227203038674e-09, 4.8084568767269302e-09, 
    4.6949349930835127e-09, 4.5869166287451755e-09, 4.485400246129317e-09, 
    4.3912713865085733e-09, 4.3052555435929037e-09, 4.2278779066895757e-09, 
    4.1594316731029755e-09, 4.0999565964471374e-09, 4.0492289306736915e-09, 
    4.0067637952655432e-09, 3.9718303321515637e-09, 3.9434796226282081e-09, 
    3.9205843967426172e-09, 3.9018889957144196e-09, 3.8860670064534215e-09, 
    3.8717834405103577e-09, 3.8577575953247497e-09, 3.8428226400805127e-09, 
    3.8259778371964297e-09, 3.8064299117223462e-09, 3.7836206719855607e-09, 
    3.7572392452198286e-09, 3.7272183052831821e-09, 3.6937152100323911e-09, 
    3.6570799262101168e-09, 3.6178128807786362e-09, 3.5765163435979567e-09, 
    3.5338434657803559e-09, 3.4904488545540839e-09, 3.4469443297218061e-09, 
    3.4038625967525727e-09, 3.3616308546412885e-09, 3.3205551736315836e-09, 
    3.2808157105853382e-09, 3.2424717649544693e-09, 3.205475232164558e-09, 
    3.1696903557761168e-09, 3.1349176641778999e-09, 3.1009197661551666e-09, 
    3.0674470547106923e-09, 3.0342614556860729e-09, 3.001156895200884e-09, 
    2.9679753821823941e-09, 2.9346181780030016e-09, 2.9010516800401051e-09, 
    2.8673082034184355e-09, 2.8334818997918617e-09, 2.7997205239915131e-09, 
    2.766213748841211e-09, 2.7331790805291635e-09, 2.7008463334318407e-09, 
    2.6694418566404951e-09, 2.6391735034710632e-09, 2.6102174251680216e-09, 
    2.5827074473959615e-09, 2.5567277834338457e-09, 2.5323093995616813e-09, 
    2.5094302800020292e-09, 2.4880193797390257e-09, 2.4679639715692699e-09, 
    2.449119654306707e-09, 2.4313222926699896e-09, 2.4144008166020204e-09, 
    2.3981899047884017e-09, 2.3825414214122939e-09, 2.3673337336335486e-09, 
    2.3524780645410505e-09, 2.3379214334189555e-09, 2.3236459217671084e-09, 
    2.3096644977035533e-09, 2.2960138016862157e-09, 2.2827447541471252e-09, 
    2.2699118856548806e-09, 2.2575625609491617e-09, 2.2457270915033316e-09, 
    2.2344107480233028e-09, 2.2235883366073814e-09, 2.2132018443331254e-09, 
    2.2031612016659794e-09, 2.1933480762898966e-09, 2.1836221704409914e-09, 
    2.1738294764358209e-09, 2.1638116463042777e-09, 2.1534157700590927e-09, 
    2.142503713565865e-09, 2.1309604229358034e-09, 2.1187005727922321e-09, 
    2.1056732665384718e-09, 2.0918644793829745e-09, 2.0772972918085175e-09, 
    2.0620299143517161e-09, 2.0461518199467753e-09, 2.0297782184521547e-09, 
    2.01304334718964e-09, 1.9960929088530742e-09, 1.9790761894997774e-09, 
    1.962138183717536e-09, 1.9454122157298155e-09, 1.9290133151501975e-09, 
    1.9130327535080209e-09, 1.8975339108987276e-09, 1.8825497616907762e-09, 
    1.8680820445890533e-09, 1.8541022602437629e-09, 1.840554406117864e-09, 
    1.8273594145701452e-09, 1.8144209919665289e-09, 1.801632610451087e-09, 
    1.7888851492312274e-09, 1.7760747650156667e-09, 1.7631103837813269e-09, 
    1.7499203525148241e-09, 1.7364577054954101e-09, 1.7227037447820297e-09, 
    1.7086696211673671e-09, 1.6943959106835831e-09, 1.6799501868058785e-09, 
    1.6654229151092214e-09, 1.6509219439103719e-09, 1.6365661148111628e-09, 
    1.6224784052797132e-09, 1.6087791426323855e-09, 1.5955796666742153e-09, 
    1.5829768423670069e-09, 1.5710486227355178e-09, 1.5598508929460312e-09, 
    1.5494155812268087e-09, 1.5397501026941217e-09, 1.5308379812177889e-09, 
    1.5226405913512748e-09, 1.5150998033103609e-09, 1.5081413905506445e-09, 
    1.501678958719455e-09, 1.4956182244380909e-09, 1.489861347331125e-09, 
    1.4843111792233313e-09, 1.4788751354970678e-09, 1.4734685631480737e-09, 
    1.468017390395961e-09, 1.4624600309918581e-09, 1.4567484165120297e-09, 
    1.4508482563781147e-09, 1.444738496343037e-09, 1.4384101810585511e-09, 
    1.4318647687151763e-09, 1.4251121145627555e-09, 1.4181682239227986e-09, 
    1.4110529703700395e-09, 1.4037878495987894e-09, 1.3963939617571808e-09, 
    1.3888902496318709e-09, 1.3812921562241544e-09, 1.3736106833778935e-09, 
    1.3658519928169532e-09, 1.3580174657064154e-09, 1.3501042863803139e-09, 
    1.3421064280932838e-09, 1.334016009596946e-09, 1.3258248476596812e-09, 
    1.317526126195687e-09, 1.3091159832300361e-09, 1.300594934875939e-09, 
    1.291968954060211e-09, 1.2832501842358706e-09, 1.2744571509693888e-09, 
    1.2656145220743223e-09, 1.2567523513785849e-09, 1.2479049169782722e-09, 
    1.2391091624444172e-09, 1.2304029060144264e-09, 1.2218228664472653e-09, 
    1.2134027370076449e-09, 1.2051713786791266e-09, 1.1971513604028866e-09, 
    1.1893579267682862e-09, 1.1817985537815585e-09, 1.1744730911745749e-09, 
    1.1673745641580532e-09, 1.1604904867970581e-09, 1.1538046410353372e-09, 
    1.1472990691927664e-09, 1.1409561488114459e-09, 1.1347604677430004e-09, 
    1.1287003853291759e-09, 1.1227690714367753e-09, 1.1169649964321524e-09, 
    1.1112917924123322e-09, 1.1057575987336812e-09, 1.1003739120087083e-09, 
    1.0951541471535253e-09, 1.0901119872899045e-09, 1.0852597353153334e-09, 
    1.0806067476809365e-09, 1.0761581215413578e-09, 1.0719136383853045e-09, 
    1.0678671068354869e-09, 1.0640060328012681e-09, 1.0603117071450227e-09, 
    1.0567595927039589e-09, 1.0533200722806769e-09, 1.0499594120087012e-09, 
    1.0466409714995974e-09, 1.0433265194821888e-09, 1.0399776622634498e-09, 
    1.0365572426503236e-09, 1.0330307193827051e-09, 1.0293674002558372e-09, 
    1.0255415326783204e-09, 1.0215331530520662e-09, 1.0173287205979982e-09, 
    1.0129214509612284e-09, 1.0083114130128324e-09, 1.0035053090924782e-09, 
    9.9851604399948621e-10, 9.9336201296326249e-10, 9.8806623411869382e-10, 
    9.8265529195327421e-10, 9.7715819939723246e-10, 9.7160519028671858e-10, 
    9.6602654292062742e-10, 9.6045142895020429e-10, 9.5490690406463546e-10, 
    9.4941701466374121e-10, 9.4400209286442105e-10, 9.3867820534301265e-10, 
    9.3345681054921304e-10, 9.2834454605052259e-10, 9.2334321242315929e-10, 
    9.1844987093785036e-10, 9.1365711092460602e-10, 9.0895344293479532e-10, 
    9.0432387454731831e-10, 8.9975061370672945e-10, 8.952139761783809e-10, 
    8.9069342436121154e-10, 8.8616875783271257e-10, 8.816213444624848e-10, 
    8.7703538412278087e-10, 8.7239903979457225e-10, 8.6770539851071143e-10, 
    8.6295311074565566e-10, 8.5814669110705667e-10, 8.5329634882191067e-10, 
    8.4841744336518324e-10, 8.4352950477175538e-10, 8.3865496905903336e-10, 
    8.3381765006945556e-10, 8.2904115984654234e-10, 8.2434731682619433e-10, 
    8.1975473435059134e-10, 8.1527762311647539e-10, 8.1092494806353126e-10, 
    8.0669992168557589e-10, 8.0259992383014025e-10, 7.9861675979071206e-10, 
    7.9473731698939462e-10, 7.9094449250143926e-10, 7.8721839730225373e-10, 
    7.8353769716702392e-10, 7.7988106677725637e-10, 7.7622859881435269e-10, 
    7.7256312566128006e-10, 7.6887129848577874e-10, 7.6514439857912587e-10, 
    7.6137874608009398e-10, 7.5757573694306143e-10, 7.5374142696192638e-10, 
    7.4988577483756683e-10, 7.4602153806989699e-10, 7.4216300394372944e-10, 
    7.383245818670754e-10, 7.3451950942372503e-10, 7.3075868704902109e-10, 
    7.2704984878718059e-10, 7.2339706429297147e-10, 7.1980069147337918e-10, 
    7.162576952169569e-10, 7.1276236296517283e-10, 7.0930726206317539e-10, 
    7.0588439644070397e-10, 7.0248635708629842e-10, 6.991074247791469e-10, 
    6.9574443732685919e-10, 6.9239738440205413e-10, 6.8906962481680272e-10, 
    6.8576776337452555e-10, 6.8250114039223352e-10, 6.7928107201767329e-10, 
    6.7611982779488445e-10, 6.7302955217574181e-10, 6.7002114698296034e-10, 
    6.6710329780980794e-10, 6.642816612659e-10, 6.6155834270217571e-10, 
    6.5893164866032881e-10, 6.5639616359007954e-10, 6.5394306603676887e-10, 
    6.5156072956569204e-10, 6.4923542385422934e-10, 6.4695216668680082e-10, 
    6.4469554859873162e-10, 6.4245054054621478e-10, 6.402031646231984e-10, 
    6.3794105398557342e-10, 6.3565381014966912e-10, 6.3333323402586523e-10, 
    6.3097336180785702e-10, 6.2857040679108619e-10, 6.2612257587407079e-10, 
    6.2362984944451792e-10, 6.2109369808012457e-10, 6.1851682383196563e-10, 
    6.1590287194850611e-10, 6.1325619396209897e-10, 6.105815739806565e-10, 
    6.0788399888898426e-10, 6.0516838220240841e-10, 6.0243931975930307e-10, 
    5.9970078728398969e-10, 5.9695589371426105e-10, 5.9420663689325653e-10, 
    5.9145374637180739e-10, 5.8869659792363128e-10, 5.8593330067264412e-10, 
    5.8316088863201875e-10, 5.8037571725237709e-10, 5.7757395387604833e-10, 
    5.7475220891230012e-10, 5.7190816472028199e-10, 5.6904121184954467e-10, 
    5.6615294334653931e-10, 5.6324749749018815e-10, 5.6033164895809827e-10, 
    5.5741466835325872e-10, 5.5450789221413667e-10, 5.5162411587866912e-10, 
    5.4877678735007222e-10, 5.4597916182452075e-10, 5.432434209596778e-10, 
    5.4057992620908255e-10, 5.3799659977656834e-10, 5.3549854432290965e-10, 
    5.3308786187789298e-10, 5.3076374040294413e-10, 5.2852270070883173e-10, 
    5.2635904432839677e-10, 5.2426537556316045e-10, 5.2223322024828533e-10, 
    5.2025362578419054e-10, 5.1831777646164421e-10, 5.1641751728165587e-10, 
    5.1454585530051202e-10, 5.1269731572436003e-10, 5.1086825188481868e-10, 
    5.0905698647815398e-10, 5.0726385363046019e-10, 5.0549107303203042e-10, 
    5.0374248937307856e-10, 5.020231296135505e-10, 5.0033866362879697e-10, 
    4.9869471644476893e-10, 4.9709617041571416e-10, 4.9554642567242526e-10, 
    4.9404677679192516e-10, 4.9259589175281239e-10, 4.9118952442961656e-10, 
    4.8982044415215258e-10, 4.8847864950058178e-10, 4.871518143465531e-10, 
    4.8582598129810989e-10, 4.8448638594496004e-10, 4.8311839543090244e-10, 
    4.8170841447005056e-10, 4.8024474270797241e-10, 4.7871823740439367e-10, 
    4.7712280306002581e-10, 4.7545560471337416e-10, 4.7371707494887485e-10, 
    4.7191066390008589e-10, 4.7004245253326691e-10, 4.6812061235487615e-10, 
    4.6615484613860952e-10, 4.6415580249664355e-10, 4.6213458336679163e-10, 
    4.6010230880689143e-10, 4.5806982588226743e-10, 4.5604748492707592e-10, 
    4.5404503544955339e-10, 4.5207154435548814e-10, 4.5013535435856455e-10, 
    4.4824400315970269e-10, 4.4640411834299043e-10, 4.446212342869887e-10, 
    4.4289957865456926e-10, 4.4124179405703132e-10, 4.3964868671976041e-10, 
    4.3811898149324199e-10, 4.3664918604589965e-10, 4.3523354004386912e-10, 
    4.3386413614734578e-10, 4.3253117051289034e-10, 4.3122336442395378e-10, 
    4.2992847291338336e-10, 4.2863390151066398e-10, 4.2732731542707795e-10, 
    4.2599723627192897e-10, 4.2463352085052766e-10, 4.2322773711249623e-10, 
    4.2177334715480073e-10, 4.2026576349724019e-10, 4.1870223216732613e-10, 
    4.1708163837118427e-10, 4.1540422518911565e-10, 4.1367133647927959e-10, 
    4.1188517837649287e-10, 4.1004868329794554e-10, 4.0816544325943996e-10, 
    4.0623975903312885e-10, 4.0427672333785326e-10, 4.0228235410371225e-10, 
    4.0026366663929761e-10, 3.9822870390382253e-10, 3.9618641999627591e-10, 
    3.94146463146503e-10, 3.921188074342669e-10, 3.901133110494726e-10, 
    3.8813920079327088e-10, 3.8620458987704265e-10, 3.8431604372339849e-10, 
    3.8247828944254018e-10, 3.8069406847721673e-10, 3.789641741699943e-10, 
    3.7728763100317082e-10, 3.7566202262869652e-10, 3.7408383893701972e-10, 
    3.7254887687396819e-10, 3.7105254325867334e-10, 3.6959008692976132e-10, 
    3.6815668288092092e-10, 3.6674741608606127e-10, 3.653571662762273e-10, 
    3.639804733856506e-10, 3.6261142340545121e-10, 3.6124366015154926e-10, 
    3.5987052522143111e-10, 3.5848541969628041e-10, 3.5708232506203517e-10, 
    3.5565649715977643e-10, 3.5420521516051506e-10, 3.5272853544214812e-10, 
    3.5122989707465163e-10, 3.4971651193856277e-10, 3.4819942023434363e-10, 
    3.4669318489351946e-10, 3.4521519106575511e-10, 3.4378460919763764e-10, 
    3.4242107398476243e-10, 3.4114323009497175e-10, 3.3996723411599301e-10, 
    3.3890541487447526e-10, 3.37965161726913e-10, 3.3714820312971748e-10, 
    3.3645027649310376e-10, 3.3586127804790083e-10, 3.3536580461591887e-10, 
    3.3494407389720404e-10, 3.3457307801460666e-10, 3.3422791708966808e-10, 
    3.3388313976048201e-10, 3.3351404296518423e-10, 3.3309780151662184e-10, 
    3.3261441793728162e-10, 3.3204740981163665e-10, 3.3138428870938419e-10, 
    3.3061679300102466e-10, 3.2974094056572763e-10, 3.2875690394661902e-10, 
    3.2766876224507796e-10, 3.2648413137111963e-10, 3.2521371830433246e-10, 
    3.2387078988205277e-10, 3.2247059815361129e-10, 3.2102973753099781e-10, 
    3.1956549961945166e-10, 3.180951868896155e-10, 3.1663546667702175e-10, 
    3.1520173564766317e-10, 3.1380755610950541e-10, 3.1246414784710705e-10, 
    3.1117998774477825e-10, 3.0996046803108795e-10, 3.0880768439737769e-10, 
    3.0772030002554012e-10, 3.0669353563806183e-10, 3.0571926469624805e-10, 
    3.0478625159616657e-10, 3.0388053586097605e-10, 3.0298599140864555e-10, 
    3.0208504288327939e-10, 3.011595680952186e-10, 3.0019192048754976e-10, 
    2.9916606103541608e-10, 2.9806868836711155e-10, 2.9689032565541857e-10, 
    2.9562621969878343e-10, 2.9427699962254034e-10, 2.9284898955096772e-10, 
    2.9135414035404992e-10, 2.89809531434302e-10, 2.8823650682961244e-10, 
    2.8665945650824202e-10, 2.8510437947705548e-10, 2.8359729666675506e-10, 
    2.821626978486997e-10, 2.8082209701562222e-10, 2.795928447104546e-10, 
    2.7848725114289838e-10, 2.7751210795135176e-10, 2.7666855831844411e-10, 
    2.7595237097663734e-10, 2.7535449536748569e-10, 2.7486186163636884e-10, 
    2.744583215414729e-10, 2.7412565119428267e-10, 2.7384450802185261e-10, 
    2.7359532242719013e-10, 2.7335900782565946e-10, 2.7311753548094769e-10, 
    2.7285430306827921e-10, 2.7255436222256972e-10, 2.7220448919336748e-10, 
    2.7179316678849951e-10, 2.7131049643888833e-10, 2.7074810278281144e-10, 
    2.7009903770448921e-10, 2.6935774398792076e-10, 2.6852006440806588e-10, 
    2.6758332843845342e-10, 2.6654646351906928e-10, 2.6541017362440027e-10, 
    2.6417707638716944e-10, 2.6285184610876161e-10, 2.614412546986097e-10, 
    2.5995415159980602e-10, 2.584012998692912e-10, 2.5679512702350203e-10, 
    2.5514934661941064e-10, 2.5347852347161852e-10, 2.5179756168053212e-10, 
    2.5012120643713129e-10, 2.4846354908127302e-10, 2.4683761065081227e-10, 
    2.4525497133725711e-10, 2.4372551970587504e-10, 2.4225725576167015e-10, 
    2.4085620895969982e-10, 2.395263853565111e-10, 2.3826980276397695e-10, 
    2.3708654817009693e-10, 2.3597489073998485e-10, 2.3493141749415188e-10, 
    2.3395122606130559e-10, 2.3302814589311257e-10, 2.3215501855072841e-10, 
    2.3132399795932407e-10, 2.3052691280671831e-10, 2.297556049070164e-10, 
    2.2900230782955662e-10, 2.2825996297726011e-10, 2.2752253592349409e-10, 
    2.2678523675107156e-10, 2.2604471414185638e-10, 2.2529913671074463e-10, 
    2.2454823462702875e-10, 2.2379322720309072e-10, 2.2303670329993378e-10, 
    2.2228239382740805e-10, 2.2153489766943901e-10, 2.2079930435221024e-10, 
    2.2008078789170432e-10, 2.1938413311279264e-10, 2.1871328032066703e-10, 
    2.1807085563467695e-10, 2.1745781218328892e-10, 2.1687313772615313e-10, 
    2.1631374491624712e-10, 2.1577449982732381e-10, 2.1524846425011432e-10, 
    2.147272695100822e-10, 2.1420166459741085e-10, 2.1366211403556725e-10, 
    2.130994575080515e-10, 2.1250549202118405e-10, 2.1187349952840155e-10, 
    2.1119857983419112e-10, 2.1047785673249059e-10, 2.0971047698444908e-10, 
    2.0889747856029368e-10, 2.0804150964515336e-10, 2.0714651143267356e-10, 
    2.0621733822972236e-10, 2.0525944884793883e-10, 2.0427861786397711e-10, 
    2.0328076786979577e-10, 2.0227184466125552e-10, 2.012578049005685e-10, 
    2.0024461011687288e-10, 1.9923827557579455e-10, 1.9824487477052041e-10, 
    1.9727054253734443e-10, 1.9632140405260901e-10, 1.9540349119283263e-10, 
    1.9452258146349391e-10, 1.9368405835468706e-10, 1.928927262534665e-10, 
    1.9215267444233368e-10, 1.9146713028935098e-10, 1.908383760253428e-10, 
    1.9026765673768031e-10, 1.8975514820023506e-10, 1.8929988886476059e-10, 
    1.8889976600983181e-10, 1.8855145491131003e-10, 1.8825040898116101e-10, 
    1.8799081973501054e-10, 1.8776565556875162e-10, 1.8756671302919021e-10, 
    1.8738478013787568e-10, 1.8720984973525921e-10, 1.8703146409531738e-10, 
    1.8683910022964542e-10, 1.8662266584300197e-10, 1.8637298751017925e-10, 
    1.8608233902933927e-10, 1.8574487764886776e-10, 1.8535704866227675e-10, 
    1.8491782315577707e-10, 1.8442883871500333e-10, 1.8389435575969791e-10, 
    1.8332110169062098e-10, 1.8271792525077767e-10, 1.8209538941721314e-10, 
    1.8146522149453285e-10, 1.8083973522472871e-10, 1.8023118705049519e-10, 
    1.7965115341247158e-10, 1.791098951506021e-10, 1.7861580336634828e-10, 
    1.78174888731372e-10, 1.7779040885824266e-10, 1.7746259213544056e-10, 
    1.7718855522855477e-10, 1.7696237436567594e-10, 1.7677538426251896e-10, 
    1.7661664140175307e-10, 1.7647361215333409e-10, 1.7633297570168505e-10, 
    1.76181574647259e-10, 1.760073591838929e-10, 1.7580032783054224e-10, 
    1.7555331052917369e-10, 1.7526258271013347e-10, 1.7492816428968807e-10, 
    1.7455384647370043e-10, 1.7414685584751043e-10, 1.7371723718314882e-10, 
    1.7327693991782531e-10, 1.7283876479949819e-10, 1.7241517756689292e-10, 
    1.7201719579122701e-10, 1.7165336742337178e-10, 1.7132901709564691e-10, 
    1.7104574374448191e-10, 1.7080130603473126e-10, 1.7058981669610431e-10, 
    1.7040230011021684e-10, 1.7022746717586029e-10, 1.70052729272565e-10, 
    1.6986526456530992e-10, 1.6965311357796075e-10, 1.694061421212085e-10, 
    1.6911685612621815e-10, 1.6878093178399249e-10, 1.6839750279855202e-10, 
    1.6796910552858734e-10, 1.6750137793037569e-10, 1.6700247139719515e-10, 
    1.6648231352542793e-10, 1.6595170092871339e-10, 1.6542140631612142e-10, 
    1.6490129270391244e-10, 1.6439958490310808e-10, 1.6392231066826104e-10, 
    1.6347301240433497e-10, 1.6305269642600926e-10, 1.6266007786385064e-10, 
    1.6229203585949329e-10, 1.6194428197424262e-10, 1.6161209085399846e-10, 
    1.6129109085860111e-10, 1.6097795412253483e-10, 1.6067096101318196e-10, 
    1.6037030976379718e-10, 1.6007821348310597e-10, 1.5979870758665915e-10, 
    1.5953724848833064e-10, 1.5930009534946989e-10, 1.5909362708941765e-10, 
    1.5892358706169311e-10, 1.5879442763048611e-10, 1.5870874557143938e-10, 
    1.5866693746538517e-10, 1.5866701690127029e-10, 1.5870468609841369e-10, 
    1.5877355056433534e-10, 1.5886551139223464e-10, 1.5897120674761189e-10, 
    1.5908052206739248e-10, 1.5918304319453822e-10, 1.592684822277953e-10, 
    1.5932698348102996e-10, 1.5934937154296813e-10, 1.5932728663259522e-10, 
    1.5925328763407513e-10, 1.5912088937541763e-10, 1.5892463192141941e-10, 
    1.5866015319557011e-10, 1.5832433350123233e-10, 1.5791546115620331e-10, 
    1.5743348290657093e-10, 1.5688025199789436e-10, 1.5625979360982274e-10, 
    1.5557849476433682e-10, 1.5484522930255629e-10, 1.5407131000549712e-10, 
    1.5327029459353764e-10, 1.5245757646158553e-10, 1.516498056128555e-10, 
    1.5086411428040548e-10, 1.5011725314622543e-10, 1.4942464058977381e-10, 
    1.4879947069911238e-10, 1.4825189230191605e-10, 1.4778840773548625e-10, 
    1.474114924408891e-10, 1.4711952893255385e-10, 1.4690701077703179e-10, 
    1.4676505830955312e-10, 1.4668214567144057e-10, 1.4664501604730772e-10, 
    1.4663964230572193e-10, 1.4665221162340632e-10, 1.4666998363402641e-10, 
    1.4668199325980421e-10, 1.4667951389290864e-10, 1.4665629216559519e-10, 
    1.466084896903676e-10, 1.4653443501609992e-10, 1.4643416358929855e-10, 
    1.463088592525749e-10, 1.4616021426060097e-10, 1.4598983511359678e-10, 
    1.4579871326657046e-10, 1.4558684907392288e-10, 1.4535302496972729e-10, 
    1.4509480221519414e-10, 1.44808667432517e-10, 1.4449038327942056e-10, 
    1.441354377114816e-10, 1.4373959381183032e-10, 1.4329945442619589e-10, 
    1.4281301778835803e-10, 1.4228012193743336e-10, 1.4170279904084828e-10, 
    1.4108545655984601e-10, 1.4043490058481438e-10, 1.3976016858911799e-10, 
    1.3907222088553945e-10, 1.3838345333012932e-10, 1.3770711945121162e-10, 
    1.3705666046836564e-10, 1.3644500612847325e-10, 1.3588385290240232e-10, 
    1.3538301752818908e-10, 1.3494985865989074e-10, 1.3458883918278216e-10, 
    1.3430121894428293e-10, 1.3408495495419701e-10, 1.3393477438858489e-10, 
    1.3384246871290859e-10, 1.3379734162123958e-10, 1.3378685695455273e-10, 
    1.3379738876348353e-10, 1.3381507742991071e-10, 1.3382668825048228e-10, 
    1.3382045730565361e-10, 1.3378682485542677e-10, 1.3371902151858408e-10, 
    1.3361344074730951e-10, 1.3346978428362693e-10, 1.3329092148145525e-10, 
    1.3308252154022023e-10, 1.3285242344381003e-10, 1.3260984113670755e-10, 
    1.3236442280322471e-10, 1.3212527738639689e-10, 1.3190001317345508e-10, 
    1.3169392127253277e-10, 1.3150931062160728e-10, 1.3134512581830472e-10, 
    1.3119682819235188e-10, 1.3105660103931037e-10, 1.3091381055222801e-10, 
    1.3075574967824932e-10, 1.3056854125594661e-10, 1.3033817534292985e-10, 
    1.3005153881652847e-10, 1.2969740504313423e-10, 1.2926724178445915e-10, 
    1.2875581688678316e-10, 1.2816151832483453e-10, 1.2748639169670839e-10, 
    1.2673586774277021e-10, 1.259182565956658e-10, 1.2504401108882771e-10, 
    1.2412488504439039e-10, 1.2317303130002616e-10, 1.2220016060702726e-10, 
    1.2121680795904444e-10, 1.2023181321168998e-10, 1.192520172256946e-10, 
    1.182822356649088e-10, 1.1732546098509077e-10, 1.1638330131716539e-10, 
    1.1545654464043438e-10, 1.145458291427159e-10, 1.1365231506584054e-10, 
    1.127782802581643e-10, 1.119275656282398e-10, 1.1110584954229691e-10, 
    1.1032067628767567e-10, 1.0958127397846633e-10, 1.0889814259827127e-10, 
    1.0828248849620055e-10, 1.0774550140922652e-10, 1.0729760202675903e-10, 
    1.0694767525627348e-10, 1.0670238194656605e-10, 1.0656557588347571e-10, 
    1.0653790163394406e-10, 1.0661655103800845e-10, 1.0679523252523492e-10, 
    1.0706429774484784e-10, 1.0741103872626566e-10, 1.0782008200726604e-10, 
    1.0827388624172704e-10, 1.0875326422769959e-10, 1.092379340525556e-10, 
    1.0970705621091001e-10, 1.1013976979374531e-10, 1.1051570215389235e-10, 
    1.1081550190706509e-10, 1.1102136712782924e-10, 1.1111761200748837e-10, 
    1.1109124378681699e-10, 1.1093255755801835e-10, 1.1063569955535926e-10, 
    1.101991699722867e-10, 1.0962620545155918e-10, 1.08924992594803e-10, 
    1.0810863652474696e-10, 1.0719488644335315e-10, 1.0620556834739221e-10, 
    1.051657656581224e-10, 1.0410274900804711e-10, 1.0304476426797017e-10, 
    1.0201971246645139e-10, 1.0105385791590796e-10, 1.0017062010319402e-10, 
    9.938955777152515e-11, 9.8725604856940038e-11, 9.8188606767239637e-11, 
    9.7783148837414302e-11, 9.7508713475182906e-11, 9.7360090414585948e-11, 
    9.7328021604462791e-11, 9.7399991350291146e-11, 9.7561124705929712e-11, 
    9.7795098615563774e-11, 9.8085031990859895e-11, 9.8414282486805887e-11, 
    9.8767133089911435e-11, 9.9129323481485641e-11, 9.9488429127847951e-11, 
    9.9834069751987202e-11, 1.0015797295130462e-10, 1.0045387991632318e-10, 
    1.0071735170844906e-10, 1.0094547430676764e-10, 1.0113652413319753e-10, 
    1.0128960605691571e-10, 1.0140433001238802e-10, 1.0148054089729546e-10, 
    1.0151814283906882e-10, 1.0151703788344425e-10, 1.0147717420873793e-10, 
    1.0139869842547995e-10, 1.012821941685338e-10, 1.0112893746284251e-10, 
    1.0094115932080055e-10, 1.0072223015742678e-10, 1.0047674483035657e-10, 
    1.0021044883820133e-10, 9.9930023127988123e-11, 9.9642700595088117e-11, 
    9.9355759512797742e-11, 9.9075945815603755e-11, 9.8808874000040508e-11, 
    9.855845895776005e-11, 9.8326480805068881e-11, 9.8112296392098194e-11, 
    9.7912771512316837e-11, 9.7722408296814977e-11, 9.7533710348410847e-11, 
    9.7337734273462273e-11, 9.7124798736307481e-11, 9.6885289546590689e-11, 
    9.6610514441894594e-11, 9.6293541507094266e-11, 9.5929955879588791e-11, 
    9.5518477252054162e-11, 9.5061402909818076e-11, 9.45648156253955e-11, 
    9.4038552218542459e-11, 9.349589085414902e-11, 9.2952986564994684e-11, 
    9.2428052417138159e-11, 9.1940344800209251e-11, 9.1508979270329721e-11, 
    9.1151690378544496e-11, 9.0883587623723207e-11, 9.0716017405501765e-11, 
    9.065562240730785e-11, 9.0703684085341699e-11, 9.0855804509676671e-11, 
    9.1101991717673835e-11, 9.1427139498704332e-11, 9.1811891747899684e-11, 
    9.2233826311190774e-11, 9.2668882595430909e-11, 9.3092902076161421e-11, 
    9.3483181442314442e-11, 9.3819890994196618e-11, 9.4087260215481057e-11, 
    9.4274425003610349e-11, 9.437589131353582e-11, 9.4391572946801514e-11, 
    9.4326440843028035e-11, 9.4189817175957851e-11, 9.3994412304721076e-11, 
    9.3755178875693492e-11, 9.3488110562645163e-11, 9.3209081811732846e-11, 
    9.2932809688715162e-11, 9.2671996972054567e-11, 9.2436715568947844e-11, 
    9.2234033679674906e-11, 9.2067875284486276e-11, 9.1939089905450309e-11, 
    9.1845706193484991e-11, 9.1783292267349277e-11, 9.1745424156366256e-11, 
    9.1724186075217996e-11, 9.1710686716495905e-11, 9.1695559037217976e-11, 
    9.1669434033187198e-11, 9.1623351879266164e-11, 9.1549132742402005e-11, 
    9.1439686168266976e-11, 9.1289272290844673e-11, 9.1093678074114694e-11, 
    9.0850371434426355e-11, 9.0558580071517341e-11, 9.0219328747845513e-11, 
    8.9835419707283777e-11, 8.9411357366847421e-11, 8.8953216080580596e-11, 
    8.8468446628034851e-11, 8.7965601155522552e-11, 8.7453998059537966e-11, 
    8.6943308251210366e-11, 8.6443084884257119e-11, 8.5962237114982201e-11, 
    8.5508488754695024e-11, 8.5087853501001023e-11, 8.4704156598591794e-11, 
    8.4358650025814164e-11, 8.4049771883084826e-11, 8.3773062720143127e-11, 
    8.3521281360780546e-11, 8.3284708895048597e-11, 8.3051636134189764e-11, 
    8.2809014933477414e-11, 8.2543208375392964e-11, 8.2240807076701149e-11, 
    8.1889444524278346e-11, 8.1478538490403108e-11, 8.0999939640661946e-11, 
    8.0448416903194576e-11, 7.9821969709307228e-11, 7.912197056816019e-11, 
    7.8353125277036649e-11, 7.7523277105650615e-11, 7.6643096069964355e-11, 
    7.5725666048120507e-11, 7.4786014461545851e-11, 7.3840580404234001e-11, 
    7.2906682576712243e-11, 7.2001940564979408e-11, 7.1143699835344713e-11, 
    7.0348444320124327e-11, 6.9631198220401295e-11, 6.900492858719893e-11, 
    6.8479980180245829e-11, 6.8063553456087523e-11, 6.7759275641656844e-11, 
    6.7566901900965311e-11, 6.7482176018842759e-11, 6.7496907737711611e-11, 
    6.7599262391516299e-11, 6.7774279882485091e-11, 6.800460436437631e-11, 
    6.8271376421940882e-11, 6.855524744739605e-11, 6.8837419901618978e-11, 
    6.9100659208599478e-11, 6.9330189654541951e-11, 6.9514416831308467e-11, 
    6.9645412083470835e-11, 6.9719159945294164e-11, 6.9735536669727046e-11, 
    6.9698062857699242e-11, 6.9613439580704889e-11, 6.949094166302086e-11, 
    6.9341695540930735e-11, 6.9177908943858995e-11, 6.9012082548814978e-11, 
    6.8856258914048077e-11, 6.8721309446686018e-11, 6.86163114057331e-11, 
    6.8548006484743993e-11, 6.8520379285751655e-11, 6.8534352517243236e-11, 
    6.858763730271899e-11, 6.8674754310158878e-11, 6.8787246116750859e-11, 
    6.8914079105882007e-11, 6.9042258821983695e-11, 6.9157621436213515e-11, 
    6.924577346103536e-11, 6.9293112006778319e-11, 6.9287866375566956e-11, 
    6.9221057821421126e-11, 6.9087308255771122e-11, 6.8885401693231464e-11, 
    6.8618556253949228e-11, 6.829435757081129e-11, 6.7924367859972253e-11, 
    6.7523425105041413e-11, 6.7108702573517795e-11, 6.669861085575784e-11, 
    6.6311630886796035e-11, 6.5965171169109015e-11, 6.5674552077671376e-11, 
    6.5452159368331394e-11, 6.5306841366407288e-11, 6.5243551107017138e-11, 
    6.5263234903955713e-11, 6.5362958865875135e-11, 6.5536219619217424e-11, 
    6.5773399449848593e-11, 6.6062342596932327e-11, 6.638897923321838e-11, 
    6.6737994026943017e-11, 6.7093498996580741e-11, 6.7439691997410787e-11, 
    6.7761486179396216e-11, 6.8045104842589234e-11, 6.8278617602221302e-11, 
    6.8452413672506663e-11, 6.8559581807648181e-11, 6.8596192747663882e-11, 
    6.8561447959879016e-11, 6.845768970579269e-11, 6.8290258419684648e-11, 
    6.8067194824731498e-11, 6.7798791673863017e-11, 6.7497033091792219e-11, 
    6.717492506298217e-11, 6.6845790486412877e-11, 6.6522552836880242e-11, 
    6.6217073404781274e-11, 6.5939571710719087e-11, 6.5698180274553665e-11, 
    6.5498666395304728e-11, 6.5344316621439314e-11, 6.5235986713814006e-11, 
    6.517232206803796e-11, 6.5150083077172441e-11, 6.5164569958622112e-11, 
    6.521008509192023e-11, 6.5280391580923793e-11, 6.5369138590656778e-11, 
    6.5470215806302919e-11, 6.5578019788493797e-11, 6.5687647932585459e-11, 
    6.5794998070555885e-11, 6.5896832972889751e-11, 6.599080397905343e-11, 
    6.6075474057202826e-11, 6.6150363726729462e-11, 6.6216025899975354e-11, 
    6.6274129009479199e-11, 6.6327563876386189e-11, 6.6380510874807984e-11, 
    6.6438452900140285e-11, 6.6508071146744907e-11, 6.6597022740755769e-11, 
    6.6713546487381318e-11, 6.6865926642041951e-11, 6.7061829089416054e-11, 
    6.7307564476883505e-11, 6.7607319633876255e-11, 6.7962479387588162e-11, 
    6.8371081525637261e-11, 6.8827500884847109e-11, 6.9322396811950899e-11, 
    6.984296985706055e-11, 7.0373507148565722e-11, 7.0896187503319238e-11, 
    7.139207306787521e-11, 7.1842212087296782e-11, 7.2228735161924113e-11, 
    7.2535869585680207e-11, 7.2750774286781879e-11, 7.2864131754159558e-11, 
    7.2870476413249604e-11, 7.2768248513624613e-11, 7.2559583467790351e-11, 
    7.2249925275991756e-11, 7.1847493925913249e-11, 7.1362696329503861e-11, 
    7.0807539613717149e-11, 7.0195105747698933e-11, 6.953912061224057e-11, 
    6.8853630676765433e-11, 6.8152778516721808e-11, 6.7450662000383235e-11, 
    6.6761217995201295e-11, 6.6098121597675103e-11, 6.5474632033708094e-11, 
    6.4903376101794307e-11, 6.4396054281197066e-11, 6.3963061542115815e-11, 
    6.3613057897728431e-11, 6.3352515614572271e-11, 6.3185293975628145e-11, 
    6.3112294168620931e-11, 6.3131240191349905e-11, 6.3236639927657916e-11, 
    6.3419933003950982e-11, 6.3669857269114514e-11, 6.397301889185286e-11, 
    6.4314624596185543e-11, 6.4679328917182157e-11, 6.505214081370812e-11, 
    6.5419302147293883e-11, 6.5769070441713454e-11, 6.6092335365693911e-11, 
    6.6383014165163492e-11, 6.6638190195213698e-11, 6.6857989489882426e-11, 
    6.7045204720433964e-11, 6.7204713172324467e-11, 6.7342739488577765e-11, 
    6.7466043919371014e-11, 6.7581106232895383e-11, 6.7693387069098621e-11, 
    6.7806727112901831e-11, 6.792293093037537e-11, 6.804157323477463e-11, 
    6.8160031209068774e-11, 6.8273725297557803e-11, 6.837654788898268e-11, 
    6.8461430464729779e-11, 6.8520990661868324e-11, 6.8548208208760636e-11, 
    6.853706273427537e-11, 6.8483085144110899e-11, 6.8383783476186547e-11, 
    6.8238892221393309e-11, 6.8050454996538376e-11, 6.782272307985327e-11, 
    6.75618918555638e-11, 6.7275695884597573e-11, 6.6972910019605061e-11, 
    6.6662807378635906e-11, 6.6354606176003929e-11, 6.6056962215581847e-11, 
    6.5777544782055411e-11, 6.5522714848066018e-11, 6.5297334143787819e-11, 
    6.5104692580165309e-11, 6.494655257972884e-11, 6.4823294412991909e-11, 
    6.473412717824662e-11, 6.4677341844907325e-11, 6.4650585782612482e-11, 
    6.465112033582299e-11, 6.4676051223184514e-11, 6.4722526911894927e-11, 
    6.4787874671928121e-11, 6.4869695905752382e-11, 6.4965907724251432e-11, 
    6.5074753435731629e-11, 6.519477294428868e-11, 6.5324747783180556e-11, 
    6.5463635828504616e-11, 6.5610499200809148e-11, 6.5764424452383922e-11, 
    6.5924454769792168e-11, 6.6089525136034613e-11, 6.6258410858924146e-11, 
    6.6429692492503557e-11, 6.6601736317166859e-11, 6.6772693537469382e-11, 
    6.6940527744659398e-11, 6.7103065846850462e-11, 6.7258065834484743e-11, 
    6.7403305839520166e-11, 6.753669936628728e-11, 6.7656400342257137e-11, 
    6.7760894438602315e-11, 6.7849069476546185e-11, 6.7920240996025979e-11, 
    6.7974119301107552e-11, 6.8010707084171114e-11, 6.8030150205881848e-11, 
    6.8032522767131932e-11, 6.8017596138394163e-11, 6.798460738260943e-11, 
    6.7932066969495184e-11, 6.7857630181423418e-11, 6.77580696326314e-11, 
    6.7629365710424591e-11, 6.7466907431155156e-11, 6.7265806115242312e-11, 
    6.7021281508938887e-11, 6.6729097634454355e-11, 6.6385990321521655e-11, 
    6.5990055805631403e-11, 6.5541049129720511e-11, 6.5040573092147497e-11, 
    6.4492125216751804e-11, 6.39010216461782e-11, 6.32741835336573e-11, 
    6.2619817170161744e-11, 6.1947017213677794e-11, 6.1265312847909184e-11, 
    6.0584205764078639e-11, 5.9912718192597175e-11, 5.9258988147718361e-11, 
    5.862993555552561e-11, 5.8031013856740793e-11, 5.7466079952910471e-11, 
    5.6937369509372482e-11, 5.6445598159457359e-11, 5.5990166264258742e-11, 
    5.5569469651147174e-11, 5.5181271907065296e-11, 5.4823117260500954e-11, 
    5.4492742646038512e-11, 5.4188443535797106e-11, 5.390936492516221e-11, 
    5.365567353508776e-11, 5.3428593450035896e-11, 5.3230314922173588e-11, 
    5.3063750641489908e-11, 5.2932188189620403e-11, 5.2838862604466579e-11, 
    5.2786492125958175e-11, 5.2776816052980971e-11, 5.2810196263411078e-11, 
    5.2885304265791401e-11, 5.2998943737040662e-11, 5.3146014892283473e-11, 
    5.331964439415357e-11, 5.3511461161774021e-11, 5.3712013386942515e-11, 
    5.3911282413179063e-11, 5.4099276480672355e-11, 5.4266636215064969e-11, 
    5.4405218138577085e-11, 5.4508597156337064e-11, 5.457246900706669e-11, 
    5.4594890190937372e-11, 5.4576353908751331e-11, 5.4519688790268315e-11, 
    5.4429790957318193e-11, 5.4313213846658458e-11, 5.4177642197047117e-11, 
    5.4031314156689039e-11, 5.388241675734484e-11, 5.3738524068630356e-11, 
    5.3606114009872028e-11, 5.349019602170808e-11, 5.3394082425266032e-11, 
    5.3319298204925407e-11, 5.3265636880727499e-11, 5.3231342894007816e-11, 
    5.3213382910308507e-11, 5.3207794692035401e-11, 5.3210060995871877e-11, 
    5.3215488359419409e-11, 5.321956020613197e-11, 5.3218240798461493e-11, 
    5.3208219219279004e-11, 5.3187085289112655e-11, 5.315342596586062e-11, 
    5.3106852510518028e-11, 5.3047957797137726e-11, 5.2978209275464619e-11, 
    5.2899787364452688e-11, 5.2815385369702678e-11, 5.2727982677707796e-11, 
    5.264060684454566e-11, 5.2556114308973611e-11, 5.2477002514643941e-11, 
    5.2405273034660129e-11, 5.2342361867211297e-11, 5.228914055147857e-11, 
    5.2245977074850014e-11, 5.2212861627307692e-11, 5.2189552696814883e-11, 
    5.21757366867926e-11, 5.217116277874156e-11 ;

 Sqw-F =
  // Sqw-F(0, 0-1999)
    0.16136447708711191, 0.16037292987799107, 0.15743758240836772, 
    0.15267366194698462, 0.14626461674834162, 0.13845007624525399, 
    0.12951059957609859, 0.1197505818031073, 0.10948078212393837, 
    0.099001872351916514, 0.088590195873806357, 0.078486613399132682, 
    0.068888938935655231, 0.059948087312207132, 0.051767708484442933, 
    0.044406808717272157, 0.037884675584239365, 0.032187338811470657, 
    0.02727480524190963, 0.023088386418068808, 0.019557568357179003, 
    0.016606030239174917, 0.014156579174830158, 0.012134913820324724, 
    0.010472248194183641, 0.0091069126441880935, 0.0079851009460679117, 
    0.0070609545341737681, 0.0062961729505271822, 0.0056593208881653674, 
    0.0051249736697229278, 0.0046728106156180074, 0.0042867340468010435, 
    0.0039540636122580479, 0.0036648327968791068, 0.0034111972899171779, 
    0.0031869530310231768, 0.0029871543937593859, 0.0028078191210180584, 
    0.002645705304856747, 0.0024981460421825063, 0.0023629287146176535, 
    0.0022382076398340832, 0.0021224407916349149, 0.0020143431851043871, 
    0.0019128512604043666, 0.0018170941215630274, 0.0017263687757338873, 
    0.0016401175723422044, 0.0015579068677794507, 0.0014794065529060226, 
    0.0014043704955547724, 0.0013326181916380974, 0.0012640180146259762, 
    0.0011984724364384749, 0.0011359054977128258, 0.0010762526659752868, 
    0.0010194530673028406, 0.00096544393580859681, 0.00091415701378992403, 
    0.0008655165638766938, 0.00081943862582878259, 0.00077583116129583654, 
    0.00073459477187573204, 0.00069562373858272084, 0.0006588072030338846, 
    0.00062403038178922125, 0.00059117576683592765, 0.00056012431132877966, 
    0.00053075662740480222, 0.00050295423192587099, 0.00047660086847678597, 
    0.0004515839137548922, 0.00042779584872311747, 0.00040513574514960163, 
    0.00038351069189540527, 0.00036283706723651239, 0.00034304155704582042, 
    0.00032406182553360014, 0.00030584676527013342, 0.00028835628429608784, 
    0.00027156062655376434, 0.00025543926280023317, 0.00023997942733695041, 
    0.00022517440638810716, 0.00021102170295608037, 0.00019752120828506035, 
    0.00018467350144119952, 0.0001724783776563048, 0.00016093367628554711, 
    0.00015003444481798318, 0.00013977244100566837, 0.00013013594508049669, 
    0.00012110983145390462, 0.00011267583607603376, 0.00010481295208069522, 
    9.7497891353455718e-05, 9.0705561067516564e-05, 8.4409519257951779e-05, 
    7.8582389286041446e-05, 7.3196227071572247e-05, 6.8222845433853037e-05, 
    6.3634105843712763e-05, 5.9402189308582331e-05, 5.5499855705377214e-05, 
    5.1900695899081613e-05, 4.8579374939383642e-05, 4.5511858996487031e-05, 
    4.2675614685540709e-05, 4.0049767817071732e-05, 3.7615209657781104e-05, 
    3.5354642257871934e-05, 3.3252559641144292e-05, 3.1295167748731272e-05, 
    2.9470251957166283e-05, 2.776700582900188e-05, 2.6175837787725817e-05, 
    2.4688173264258197e-05, 2.3296268518929726e-05, 2.1993049131381276e-05, 
    2.0771981655448323e-05, 1.9626981896212759e-05, 1.8552358432117501e-05, 
    1.7542786026936579e-05, 1.6593300901688354e-05, 1.5699308667886993e-05, 
    1.4856596004754862e-05, 1.4061338630056416e-05, 1.3310100355892577e-05, 
    1.2599820575056706e-05, 1.1927789954358523e-05, 1.129161608435732e-05, 
    1.0689182148298833e-05, 1.0118602276947607e-05, 9.578177220754841e-06, 
    9.0663534600597907e-06, 8.5816880819838006e-06, 8.122820870812585e-06, 
    7.6884542278882854e-06, 7.2773408420163091e-06, 6.8882784918521886e-06, 
    6.5201109564450811e-06, 6.1717336956123265e-06, 5.8421027043167243e-06, 
    5.5302447311574683e-06, 5.2352669063324889e-06, 4.9563637946536751e-06, 
    4.6928200380841225e-06, 4.4440071255641219e-06, 4.2093734425906487e-06, 
    3.9884275734743018e-06, 3.780715771031033e-06, 3.585795440539632e-06, 
    3.403207260633526e-06, 3.2324490379068547e-06, 3.0729544635837795e-06, 
    2.9240795626464435e-06, 2.7850988318957601e-06, 2.6552119513130963e-06, 
    2.5335606829809443e-06, 2.4192543258544509e-06, 2.3114010568363599e-06, 
    2.2091418036712743e-06, 2.1116830539947067e-06, 2.0183252230348528e-06, 
    1.9284838320788537e-06, 1.8417016797362022e-06, 1.7576512788572321e-06, 
    1.6761279279288573e-06, 1.597034750494343e-06, 1.520361761780076e-06, 
    1.4461614465196197e-06, 1.3745234373857137e-06, 1.3055506958704289e-06, 
    1.2393391693160471e-06, 1.1759623081058551e-06, 1.1154611552553416e-06, 
    1.0578400518221568e-06, 1.0030674030910795e-06, 9.5108048257067258e-07, 
    9.0179294702591352e-07, 8.5510361802964739e-07, 8.1090514652263486e-07, 
    7.6909139834782794e-07, 7.2956273778116682e-07, 6.9222879455666599e-07, 
    6.570087174751933e-07, 6.2382929119151999e-07, 5.9262157212325299e-07, 
    5.6331685586501399e-07, 5.3584280662702967e-07, 5.101204701697755e-07, 
    4.8606267967016286e-07, 4.6357409109048268e-07, 4.4255279543824609e-07, 
    4.2289319704212067e-07, 4.0448965452854089e-07, 3.8724028163254322e-07, 
    3.7105030412880467e-07, 3.5583446293241611e-07, 3.4151812013010883e-07, 
    3.2803693721052059e-07, 3.1533521785403101e-07, 3.0336321114561713e-07, 
    2.9207382443875041e-07, 2.8141928098669473e-07, 2.7134826351682711e-07, 
    2.6180401508008176e-07, 2.5272373077808794e-07, 2.4403939148438465e-07, 
    2.3567998580990967e-07, 2.2757487019442008e-07, 2.1965785340521976e-07, 
    2.1187148479531466e-07, 2.0417098783852049e-07, 1.9652731776659037e-07, 
    1.8892892729319639e-07, 1.8138198408754728e-07, 1.739089737586101e-07, 
    1.6654581918139631e-07, 1.5933782284262322e-07, 1.5233487285227622e-07, 
    1.4558642867692613e-07, 1.3913681281112631e-07, 1.3302128044942586e-07, 
    1.2726323144309218e-07, 1.2187278324823457e-07, 1.1684676044450451e-07, 
    1.1216999668129313e-07, 1.0781770801765389e-07, 1.037585965296863e-07, 
    9.995829031046171e-08, 9.6382721592865892e-08, 9.3001086762405377e-08, 
    8.9788110367711083e-08, 8.6725438787155121e-08, 8.3802102263049653e-08, 
    8.1014093850879635e-08, 7.8363206743237402e-08, 7.5855339492080772e-08, 
    7.3498514987231021e-08, 7.1300864070236059e-08, 6.9268799542319537e-08, 
    6.7405558294762449e-08, 6.5710225175947755e-08, 6.4177282434869147e-08, 
    6.2796660992824907e-08, 6.1554214018194921e-08, 6.043249382988864e-08, 
    5.9411695097839904e-08, 5.8470630035686758e-08, 5.7587623525217637e-08, 
    5.6741251813752383e-08, 5.5910892136341172e-08, 5.5077092876706881e-08, 
    5.4221809298216898e-08, 5.3328570736526384e-08, 5.238264983699927e-08, 
    5.1371291379295577e-08, 5.0284032076316146e-08, 4.91131073392122e-08, 
    4.7853905746236065e-08, 4.6505401989982381e-08, 4.5070482846113765e-08, 
    4.3556079576864124e-08, 4.1973037166180668e-08, 4.0335681099705445e-08, 
    3.8661082371481702e-08, 3.6968063801300878e-08, 3.5276028404188631e-08, 
    3.360371775333681e-08, 3.1968020965006232e-08, 3.0382951581286295e-08, 
    2.885889152425237e-08, 2.7402171077576764e-08, 2.6015017420582782e-08, 
    2.4695864536728659e-08, 2.343998173835152e-08, 2.224034767026777e-08, 
    2.1088676570230121e-08, 1.9976492702934575e-08, 1.8896149402200043e-08, 
    1.7841698145050145e-08, 1.6809531237041018e-08, 1.5798744738071813e-08, 
    1.4811196677867788e-08, 1.3851264523180295e-08, 1.2925335005682829e-08, 
    1.2041084653372991e-08, 1.1206629486187485e-08, 1.0429634111537183e-08, 
    9.7164736642320845e-09, 9.0715346046410794e-09, 8.4967245041696866e-09, 
    7.9912362363041144e-09, 7.5515837121199149e-09, 7.1718950743893071e-09, 
    6.8444217036921384e-09, 6.5601984595986444e-09, 6.3097772741094611e-09, 
    6.0839520157571625e-09, 5.8743994795917397e-09, 5.6741762329790094e-09, 
    5.4780333337050095e-09, 5.2825351574402629e-09, 5.0859934064620346e-09, 
    4.8882473880805167e-09, 4.6903363784996087e-09, 4.494115960407259e-09, 
    4.3018695563597939e-09, 4.1159578151669497e-09, 3.9385364537402684e-09, 
    3.7713576452352959e-09, 3.6156560341293479e-09, 3.4721083121161307e-09, 
    3.3408480410026046e-09, 3.2215143826984667e-09, 3.113315663617649e-09, 
    3.0150936780655166e-09, 2.9253819633987455e-09, 2.8424579775850369e-09, 
    2.7643949920582296e-09, 2.6891216426524305e-09, 2.6144969412430742e-09, 
    2.5384050651766684e-09, 2.4588692008630666e-09, 2.3741779598017419e-09, 
    2.2830128289652516e-09, 2.1845620916340603e-09, 2.0786063020397461e-09, 
    1.9655625713683566e-09, 1.8464797062868937e-09, 1.7229822356021876e-09, 
    1.597168056587881e-09, 1.4714700914020919e-09, 1.3484964166779167e-09, 
    1.2308652029756683e-09, 1.1210501310467395e-09, 1.0212489873558684e-09, 
    9.3328399156715912e-10, 8.5853707284314146e-10, 7.9791869701552508e-10, 
    7.518647419633671e-10, 7.2035385488562864e-10, 7.0293713583720481e-10, 
    6.9877323129015378e-10, 7.0666435892336767e-10, 7.2509192074177276e-10, 
    7.5225305241818797e-10, 7.8610174656815507e-10, 8.2439871232356348e-10, 
    8.6477352404974235e-10, 9.0480049261651541e-10, 9.4208667848704643e-10, 
    9.7436732993857182e-10, 9.9960124096023187e-10, 1.0160569078282615e-09, 
    1.0223804328457215e-09, 1.0176374202408619e-09, 1.0013244435568799e-09, 
    9.7334930080233535e-10, 9.3398356103898564e-10, 8.8379439169065028e-10, 
    8.2356530693308878e-10, 7.5421609211997547e-10, 6.7673177533416313e-10, 
    5.9210785809445806e-10, 5.0131623945027343e-10, 4.0529209803835291e-10, 
    3.049390961837339e-10, 2.0114721393490929e-10, 9.4816393210914468e-11, 
    -1.312118789757855e-11, -1.2168600256649056e-10, -2.2984741626263447e-10, 
    -3.3653233614393561e-10, -4.4064554335010656e-10, 
    -5.4109824208987382e-10, -6.3684059727907791e-10, 
    -7.2689345821513993e-10, -8.1037523828118242e-10, -8.865213105582918e-10, 
    -9.5469523971553829e-10, -1.0143928895852122e-09, 
    -1.0652423729714043e-09, -1.1070032466194471e-09, 
    -1.1395687323064353e-09, -1.1629734902168533e-09, 
    -1.1774079157328486e-09, -1.1832375588513342e-09, 
    -1.1810244420825093e-09, -1.1715447023524373e-09, 
    -1.1557967367280997e-09, -1.1349937156361591e-09, 
    -1.1105361343962878e-09, -1.0839621053444173e-09, 
    -1.0568766404622605e-09, -1.0308639725848257e-09, 
    -1.0073902490218445e-09, -9.8770585940199749e-10, 
    -9.7275761391989101e-10, -9.6312045757852167e-10, -9.589567620319394e-10, 
    -9.6000828764250786e-10, -9.6562259044561024e-10, 
    -9.7481179672931196e-10, -9.8633844609831401e-10, 
    -9.9882020734742117e-10, -1.0108436042924088e-09, 
    -1.0210761742116106e-09, -1.0283670630726436e-09, 
    -1.0318273239123176e-09, -1.0308837251253173e-09, 
    -1.0253025490834534e-09, -1.0151828563352647e-09, 
    -1.0009217160269127e-09, -9.8315625820044338e-10, 
    -9.6268941519087305e-10, -9.4040727898809852e-10, 
    -9.1719607485187303e-10, -8.9386641864093151e-10, 
    -8.7109096649532086e-10, -8.4935991642461148e-10, 
    -8.2895664562805388e-10, -8.0995372637143147e-10, 
    -7.9222756653801917e-10, -7.7548855241945349e-10, 
    -7.5932234682491369e-10, -7.4323775218067641e-10, 
    -7.2671626144793141e-10, -7.0925914528928058e-10, 
    -6.9042839341441465e-10, -6.6987897502142599e-10, 
    -6.4738072664057245e-10, -6.2282945284335926e-10, -5.962473883471355e-10, 
    -5.6777449717874354e-10, -5.3765214121981049e-10, 
    -5.0620160047180951e-10, -4.7379972172646765e-10, 
    -4.4085416276555162e-10, -4.0778021156621972e-10, -3.749809710289324e-10, 
    -3.4283175085720586e-10, -3.116692088246429e-10, -2.8178490800658549e-10, 
    -2.5342266987745215e-10, -2.2677861125168573e-10, 
    -2.0200279880949216e-10, -1.7920143609219725e-10, 
    -1.5843897440303813e-10, -1.3973964979783085e-10, -1.230887376999774e-10, 
    -1.0843382220672532e-10, -9.5686910303983067e-11, 
    -8.4728003251773724e-11, -7.5410855320272659e-11, 
    -6.7571000575371119e-11, -6.1036007140742447e-11, 
    -5.5637083063983736e-11, -5.122107503382039e-11, -4.7661277487111793e-11, 
    -4.4865662361955061e-11, -4.2781091502505297e-11, 
    -4.1392665262170312e-11, -4.0717733052875187e-11, 
    -4.0795048915375626e-11, -4.1669986919432197e-11, 
    -4.3377580263888214e-11, -4.5925368807733704e-11, 
    -4.9278313978102751e-11, -5.3347780942342901e-11, 
    -5.7986234439804845e-11, -6.298863795684959e-11, -6.8100677533867614e-11, 
    -7.3033269536815905e-11, -7.74819976759528e-11, -8.1149506234801031e-11, 
    -8.3768853611805776e-11, -8.5125335214778735e-11, 
    -8.5074992950278487e-11, -8.3557968777304165e-11, 
    -8.0605808472974989e-11, -7.6342137149932138e-11, 
    -7.0976952155010889e-11, -6.4795111149468629e-11, 
    -5.8140230390848729e-11, -5.1395199346314672e-11, -4.496089248255838e-11, 
    -3.9234429917742718e-11, -3.4588405101336589e-11, -3.135204476405966e-11, 
    -2.9795318452990064e-11, -3.0116479759278886e-11, -3.243354319866762e-11, 
    -3.677977413525342e-11, -4.3103289095252649e-11, -5.1270578188207027e-11, 
    -6.1073751533399743e-11, -7.224110211335509e-11, -8.4450536513783e-11, 
    -9.7345173113073138e-11, -1.1055042641929599e-10, 
    -1.2369158978821725e-10, -1.3641105696154557e-10, 
    -1.4838409786327352e-10, -1.5933239938520855e-10, 
    -1.6903451682356346e-10, -1.7733283589042308e-10, 
    -1.8413672082816722e-10, -1.8942196219049648e-10, 
    -1.9322678925370163e-10, -1.9564497812739127e-10, 
    -1.9681662007720879e-10, -1.9691725100221659e-10, 
    -1.9614591338705963e-10, -1.9471280800184232e-10, 
    -1.9282702984380576e-10, -1.9068495860501984e-10, 
    -1.8845980160998412e-10, -1.8629288801693988e-10, 
    -1.8428724097948287e-10, -1.8250390782737586e-10, 
    -1.8096151100290001e-10, -1.7963910496279764e-10, 
    -1.7848231281709881e-10, -1.7741223140435834e-10, 
    -1.7633637469893055e-10, -1.7516067766137398e-10, 
    -1.7380125810426767e-10, -1.7219482934775672e-10, 
    -1.7030667098406985e-10, -1.6813539805292035e-10, 
    -1.6571411149991052e-10, -1.6310798713802387e-10, 
    -1.6040866099293333e-10, -1.5772626703463718e-10, 
    -1.5517998826284449e-10, -1.528882213068693e-10, -1.5095934824346203e-10, 
    -1.494839669529538e-10, -1.4852915428845292e-10, -1.4813512841551438e-10, 
    -1.4831434793767409e-10, -1.4905289545726396e-10, 
    -1.5031368990766218e-10, -1.5204116382535984e-10, 
    -1.5416666014486616e-10, -1.5661412321115083e-10, -1.593054823644214e-10, 
    -1.6216538098330763e-10, -1.6512485835754388e-10, 
    -1.6812392100791557e-10, -1.7111284661145746e-10, 
    -1.7405242456404561e-10, -1.7691317274997013e-10, 
    -1.7967389369949203e-10, -1.8231971381091706e-10, 
    -1.8483998610223312e-10, -1.8722618988472436e-10, -1.894701148066938e-10, 
    -1.9156233215212501e-10, -1.9349113827338127e-10, 
    -1.9524181832088013e-10, -1.9679638061140756e-10, -1.981334779337647e-10, 
    -1.9922863674940799e-10, -2.0005461584063916e-10, 
    -2.0058201218696398e-10, -2.0077995253133151e-10, 
    -2.0061713755342317e-10, -2.000630345960067e-10, -1.9908947644955264e-10, 
    -1.9767253349476191e-10, -1.9579464888279884e-10, 
    -1.9344695026564996e-10, -1.9063156822033751e-10, -1.873637274478962e-10, 
    -1.8367346002881877e-10, -1.7960656153500076e-10, 
    -1.7522476219437451e-10, -1.7060478051585953e-10, 
    -1.6583635269368114e-10, -1.6101908769086303e-10, 
    -1.5625843835050584e-10, -1.5166081979013953e-10, -1.473283372652622e-10, 
    -1.4335330994679638e-10, -1.3981315190428237e-10, 
    -1.3676582598787991e-10, -1.3424637996933296e-10, -1.322647172251195e-10, 
    -1.3080493967784111e-10, -1.298261898720869e-10, -1.2926512860369093e-10, 
    -1.2903971733798746e-10, -1.2905413836286607e-10, 
    -1.2920443450246411e-10, -1.2938452598989091e-10, 
    -1.2949204506166701e-10, -1.2943374094869952e-10, 
    -1.2912998413715488e-10, -1.2851817844575301e-10, 
    -1.2755488840775252e-10, -1.2621667491092322e-10, 
    -1.2449961682735354e-10, -1.2241779238111969e-10, 
    -1.2000079677361937e-10, -1.1729066506053916e-10, -1.143384194635165e-10, 
    -1.1120057135714788e-10, -1.0793575599493653e-10, 
    -1.0460181190500436e-10, -1.0125333232501419e-10, 
    -9.7939888454114207e-11, -9.4704861160408585e-11, -9.158491901079751e-11, 
    -8.8609991427191553e-11, -8.5803665209999592e-11, 
    -8.3183843569524714e-11, -8.0763560363805589e-11, 
    -7.8551829472157465e-11, -7.6554410794443036e-11, 
    -7.4774471440099357e-11, -7.3213132692002831e-11, 
    -7.1869838591066782e-11, -7.0742606950428984e-11, 
    -6.9828159044892937e-11, -6.9121973542838671e-11, 
    -6.8618206790696819e-11, -6.8309535672102023e-11, 
    -6.8186898295076255e-11, -6.8239140194589828e-11, -6.845259688154466e-11, 
    -6.8810625047680524e-11, -6.9293161682588158e-11, 
    -6.9876421064508214e-11, -7.0532717160792213e-11, 
    -7.1230630466722338e-11, -7.1935424380254715e-11, -7.260989815842158e-11, 
    -7.3215537445601055e-11, -7.3714034345635802e-11, 
    -7.4068962440871244e-11, -7.4247643431287647e-11, -7.422291599802762e-11, 
    -7.397477810878575e-11, -7.3491676970406271e-11, -7.2771430393369511e-11, 
    -7.1821592997553974e-11, -7.0659313389426256e-11, 
    -6.9310619093718962e-11, -6.780926224688504e-11, -6.6195105992604663e-11, 
    -6.4512262055308171e-11, -6.2807027456308314e-11, 
    -6.1125843380796884e-11, -5.9513307112134632e-11, 
    -5.8010412839686143e-11, -5.6653050471520656e-11, 
    -5.5470863933363084e-11, -5.4486419376693461e-11, -5.371473578482379e-11, 
    -5.3163125314909948e-11, -5.2831336257927674e-11, 
    -5.2711958805785487e-11, -5.2791045391882219e-11, 
    -5.3048956738778178e-11, -5.3461414018931551e-11, 
    -5.4000719219823153e-11, -5.463707635762672e-11, -5.5340025811231428e-11, 
    -5.607990145365486e-11, -5.682920001748421e-11, -5.7563827041009377e-11, 
    -5.8264038995923835e-11, -5.8915120601251844e-11, 
    -5.9507603961424364e-11, -6.0037131244572865e-11, 
    -6.0503868254602077e-11, -6.0911639256561669e-11, 
    -6.1266769300725481e-11, -6.1576884444568317e-11, 
    -6.1849668896503932e-11, -6.209181871977495e-11, -6.2308252031014208e-11, 
    -6.2501649427002244e-11, -6.2672349679495716e-11, -6.281862361528462e-11, 
    -6.2937188033748462e-11, -6.3023969471799616e-11, 
    -6.3074907195605639e-11, -6.3086810420098478e-11, 
    -6.3058032834925894e-11, -6.2989018825834941e-11, 
    -6.2882574507165494e-11, -6.2743931852067474e-11, 
    -6.2580539921988487e-11, -6.2401669153523481e-11, 
    -6.2217857004470397e-11, -6.2040243893616003e-11, 
    -6.1879868512602726e-11, -6.174697205149453e-11, -6.1650317630014382e-11, 
    -6.1596672122414075e-11, -6.1590324673464434e-11, 
    -6.1632830871601275e-11, -6.172286795789649e-11, -6.1856312786114311e-11, 
    -6.2026424896600745e-11, -6.2224268058423212e-11, 
    -6.2439189894016493e-11, -6.2659445250131226e-11, -6.287278620336904e-11, 
    -6.3067157249783809e-11, -6.3231228508621942e-11, -6.335488069761159e-11, 
    -6.3429542633635731e-11, -6.3448412704130025e-11, 
    -6.3406512444789808e-11, -6.3300643003629442e-11, 
    -6.3129234348702191e-11, -6.2892160726080151e-11, 
    -6.2590530806503019e-11, -6.2226481317779468e-11, 
    -6.1803024562996764e-11, -6.1323939380687123e-11, 
    -6.0793686780891132e-11, -6.0217363402579701e-11, 
    -5.9600669923159553e-11, -5.8949831628772722e-11, 
    -5.8271515490323882e-11, -5.7572676128423171e-11, 
    -5.6860358939839398e-11, -5.6141499149613694e-11, -5.542266598177318e-11, 
    -5.4709851004773577e-11, -5.4008285371961752e-11, 
    -5.3322339066729096e-11, -5.2655484403431281e-11, -5.201035160422211e-11, 
    -5.1388858164506626e-11, -5.0792377384292605e-11, 
    -5.0221928761479321e-11, -4.9678384203668321e-11, 
    -4.9162587764291643e-11, -4.8675470586730863e-11, 
    -4.8218069611946291e-11, -4.7791495076068687e-11, 
    -4.7396811484043405e-11, -4.7034991147980463e-11, 
    -4.6706765043682787e-11, -4.641254192010135e-11, -4.6152345108816579e-11, 
    -4.592583006620561e-11, -4.5732269120101104e-11, -4.5570652402260277e-11, 
    -4.5439699663594603e-11, -4.5337910861696078e-11, -4.526353662609192e-11, 
    -4.5214527691198337e-11, -4.5188379219333424e-11, 
    -4.5181983728053434e-11, -4.5191414133192044e-11, 
    -4.5211764134006079e-11, -4.5236984254543799e-11, 
    -4.5259904931651343e-11, -4.5272302521525259e-11, 
    -4.5265149607861545e-11, -4.5228976809413799e-11, 
    -4.5154407249071642e-11, -4.503270598164851e-11, -4.4856404468277355e-11, 
    -4.4619861431961911e-11, -4.4319725350428609e-11, 
    -4.3955232934646338e-11, -4.3528371897600295e-11, 
    -4.3043751948217403e-11, -4.2508370237338351e-11, 
    -4.1931139302444202e-11, -4.1322325037172014e-11, 
    -4.0692899722561087e-11, -4.0053886909027705e-11, 
    -3.9415753847156535e-11, -3.8787875343596329e-11, 
    -3.8178116160598721e-11, -3.7592544177567803e-11, -3.703526707760013e-11, 
    -3.6508398545435262e-11, -3.6012125322759386e-11, 
    -3.5544886568055562e-11, -3.5103649174262728e-11, 
    -3.4684205572841523e-11, -3.4281591388035748e-11, 
    -3.3890528865747282e-11, -3.3505912114880531e-11, 
    -3.3123303989574654e-11, -3.273939940347908e-11, -3.2352470681633267e-11, 
    -3.1962657916022332e-11, -3.157216838007568e-11, -3.1185252191055099e-11, 
    -3.0808033199118274e-11, -3.0448060048939353e-11, 
    -3.0113747586640418e-11, -2.9813641887828797e-11, 
    -2.9555625384507897e-11, -2.9346097496818405e-11, 
    -2.9189313898215525e-11, -2.9086828263264555e-11, 
    -2.9037197461376141e-11, -2.9035974620167061e-11, 
    -2.9075964280838912e-11, -2.9147759085474779e-11, 
    -2.9240506128756629e-11, -2.9342787891052506e-11, 
    -2.9443587329971038e-11, -2.9533175432680541e-11, -2.960391738036195e-11, 
    -2.9650845127719167e-11, -2.9671996504749437e-11, 
    -2.9668475509653057e-11, -2.9644253494484647e-11, 
    -2.9605733401994915e-11, -2.9561120059977793e-11, 
    -2.9519660590307088e-11, -2.9490833726992958e-11, 
    -2.9483525692503987e-11, -2.9505289027972959e-11, 
    -2.9561687716896974e-11, -2.9655823458437018e-11, 
    -2.9787980685993437e-11, -2.995551002866235e-11, -3.0152838319026363e-11, 
    -3.037168898311113e-11, -3.0601419968364292e-11, -3.0829537567596921e-11, 
    -3.1042289370376575e-11, -3.122536724242135e-11, -3.136464755040162e-11, 
    -3.1446982395941795e-11, -3.1460938420779759e-11, 
    -3.1397528031760036e-11, -3.1250788473737657e-11, 
    -3.1018289570412959e-11, -3.0701406257743422e-11, 
    -3.0305428018738543e-11, -2.9839423861935181e-11, 
    -2.9315917100553119e-11, -2.8750323922754679e-11, 
    -2.8160240263198847e-11, -2.7564597041021025e-11, -2.698274836816937e-11, 
    -2.64335502380222e-11, -2.593448781308676e-11, -2.5500909940896673e-11, 
    -2.5145394435854996e-11, -2.487729354045542e-11, -2.4702418157970003e-11, 
    -2.4622954114447647e-11, -2.4637455251782624e-11, 
    -2.4741037275403084e-11, -2.4925652481285597e-11, 
    -2.5180490067685164e-11, -2.5492421263464191e-11, 
    -2.5846548655101242e-11, -2.6226796693218442e-11, 
    -2.6616549682755161e-11, -2.6999328695529923e-11, 
    -2.7359463074136702e-11, -2.7682752462855119e-11, 
    -2.7957059025888638e-11, -2.8172827326019873e-11, 
    -2.8323436897026162e-11, -2.8405429999550337e-11, 
    -2.8418528061675673e-11, -2.8365467808081754e-11, 
    -2.8251659371360701e-11, -2.8084697132370911e-11, 
    -2.7873768213761016e-11, -2.7628994771950891e-11, 
    -2.7360780775921507e-11, -2.7079228699314951e-11, 
    -2.6793626761790804e-11, -2.6512084470292175e-11, 
    -2.6241270379433348e-11, -2.598635048864733e-11, -2.5750983608053195e-11, 
    -2.5537463781126145e-11, -2.5346891107722171e-11, 
    -2.5179413131446384e-11, -2.5034452970341541e-11, 
    -2.4910906070794486e-11, -2.4807307351960112e-11, 
    -2.4721955550289671e-11, -2.4652977188210763e-11, 
    -2.4598344779611218e-11, -2.4555860937731002e-11, 
    -2.4523128402864943e-11, -2.4497527967400102e-11, 
    -2.4476179034007234e-11, -2.4455982916552604e-11, 
    -2.4433665432107474e-11, -2.4405910058941443e-11, 
    -2.4369495272024408e-11, -2.4321506478931855e-11, 
    -2.4259524177450244e-11, -2.4181834393129056e-11, 
    -2.4087569716786367e-11, -2.3976813969224306e-11, 
    -2.3850600845386348e-11, -2.3710840220834455e-11, 
    -2.3560133393755135e-11, -2.3401521310350499e-11, 
    -2.3238177969805898e-11, -2.3073078941458019e-11, -2.2908692920707e-11, 
    -2.2746711424076575e-11, -2.2587879226189595e-11, 
    -2.2431910759970661e-11, -2.227753041744486e-11, -2.2122620870516172e-11, 
    -2.1964453923601305e-11, -2.1799991865731856e-11, 
    -2.1626234027186126e-11, -2.144057227760665e-11, -2.1241076054388747e-11, 
    -2.1026767082022802e-11, -2.0797803072931239e-11, 
    -2.0555553356570924e-11, -2.0302631573097447e-11, 
    -2.0042800921805541e-11, -1.9780832156763257e-11, 
    -1.9522274724914805e-11, -1.9273224461423746e-11, 
    -1.9040010856402705e-11, -1.8828894503553881e-11, 
    -1.8645726917631132e-11, -1.8495646182022006e-11, 
    -1.8382737149629462e-11, -1.8309768728104994e-11, 
    -1.8277894363188873e-11, -1.8286514688382426e-11, 
    -1.8333129885294903e-11, -1.8413339898752902e-11, 
    -1.8520945648043963e-11, -1.8648193504190341e-11, 
    -1.8786116331798753e-11, -1.8925032520373612e-11, 
    -1.9055090696961982e-11, -1.916688707531252e-11, -1.9252037663783427e-11, 
    -1.9303771690223465e-11, -1.9317316528875382e-11, 
    -1.9290215825908848e-11, -1.9222391673611779e-11, 
    -1.9116083757531037e-11, -1.89755493457031e-11, -1.8806650940587332e-11, 
    -1.8616320683697735e-11, -1.8411998819143012e-11, -1.820104859413791e-11, 
    -1.7990280050244108e-11, -1.7785527384173072e-11, 
    -1.7591402626679447e-11, -1.7411135972004784e-11, 
    -1.7246582675858834e-11, -1.7098286178339139e-11, 
    -1.6965640701018151e-11, -1.6847061509085728e-11, 
    -1.6740197010808132e-11, -1.6642080098861543e-11, 
    -1.6549328105528142e-11, -1.6458272697336387e-11, 
    -1.6365096624190749e-11, -1.6265973797890982e-11, 
    -1.6157249936506273e-11, -1.6035607206752926e-11, 
    -1.5898281323263225e-11, -1.5743240984554698e-11, 
    -1.5569421570274505e-11, -1.5376838310709821e-11, 
    -1.5166733026431508e-11, -1.4941547467922272e-11, 
    -1.4704864285396525e-11, -1.4461221612175062e-11, 
    -1.4215862085950621e-11, -1.3974388517453367e-11, -1.374242646536685e-11, 
    -1.3525251892136532e-11, -1.3327467067111692e-11, 
    -1.3152721002119191e-11, -1.3003554298784538e-11, 
    -1.2881288355877767e-11, -1.2786041054211922e-11, 
    -1.2716803729491959e-11, -1.2671614607655623e-11, 
    -1.2647747319064754e-11, -1.2641954600524828e-11, -1.265069905109743e-11, 
    -1.2670386839615106e-11, -1.269757679222775e-11, -1.2729183507874467e-11, 
    -1.2762613570011313e-11, -1.2795904435909923e-11, 
    -1.2827812153829778e-11, -1.2857888754038965e-11, 
    -1.2886505016579926e-11, -1.291483700434183e-11, -1.2944818685448251e-11, 
    -1.2979012069374562e-11, -1.3020461255053402e-11, -1.307245606832188e-11, 
    -1.3138272782971901e-11, -1.3220860338658525e-11, -1.332253297322418e-11, 
    -1.3444644987878415e-11, -1.358732725605039e-11, -1.3749286354268936e-11, 
    -1.3927692734868343e-11, -1.411817778653061e-11, -1.431497360203142e-11, 
    -1.4511132983818977e-11, -1.4698913461657353e-11, 
    -1.4870181706367918e-11, -1.5016913693709025e-11, 
    -1.5131685938611264e-11, -1.5208148265974487e-11, 
    -1.5241420680963514e-11, -1.5228412881053632e-11, 
    -1.5168037295468148e-11, -1.5061266288344174e-11, 
    -1.4911109315376164e-11, -1.4722424372455599e-11, 
    -1.4501667436664321e-11, -1.4256522368754784e-11, 
    -1.3995510172935831e-11, -1.3727535037725101e-11, 
    -1.3461450496064884e-11, -1.3205634659341032e-11, 
    -1.2967624960848458e-11, -1.2753805537608239e-11, 
    -1.2569187562754569e-11, -1.2417270974672978e-11, 
    -1.2300002944725501e-11, -1.2217807228589986e-11, 
    -1.2169706578160304e-11, -1.2153485683207124e-11, 
    -1.2165901689298371e-11, -1.2202944627489078e-11, 
    -1.2260050551927037e-11, -1.2332341845460682e-11, -1.241488557360181e-11, 
    -1.2502868806132341e-11, -1.2591779603031098e-11, -1.267756037382742e-11, 
    -1.275672265436199e-11, -1.2826433130467739e-11, -1.2884580634371609e-11, 
    -1.2929794884609895e-11, -1.2961449277337052e-11, 
    -1.2979614569253928e-11, -1.2985014211712517e-11, 
    -1.2978923313797709e-11, -1.2963062170694963e-11, 
    -1.2939462416556368e-11, -1.2910341818140073e-11, -1.2877936002214e-11, 
    -1.2844364321986357e-11, -1.2811467676868884e-11, 
    -1.2780676356046204e-11, -1.2752883049430418e-11, 
    -1.2728329482200486e-11, -1.2706545241270147e-11, 
    -1.2686321101321307e-11, -1.2665721264830274e-11, 
    -1.2642200455380357e-11, -1.2612741222866606e-11, 
    -1.2574071089271997e-11, -1.2522931174809083e-11, 
    -1.2456379364017744e-11, -1.2372083299737303e-11, 
    -1.2268610251858926e-11, -1.2145636519886325e-11, 
    -1.2004076950650996e-11, -1.1846120817542368e-11, 
    -1.1675113140432592e-11, -1.1495335848730581e-11, 
    -1.1311711952235356e-11, -1.1129382888677622e-11, -1.095330470895381e-11, 
    -1.0787829173936526e-11, -1.0636344717470859e-11, 
    -1.0501048811656827e-11, -1.0382782986495115e-11, -1.028107729726407e-11, 
    -1.0194270975897393e-11, -1.011979231361635e-11, -1.0054506019196672e-11, 
    -9.9951091052266377e-12, -9.9385187335614135e-12, 
    -9.8822378956404691e-12, -9.8246051987711268e-12, 
    -9.7649777337055531e-12, -9.7037624125338446e-12, 
    -9.6423617494718063e-12, -9.5829907642264388e-12, 
    -9.5284287994121922e-12, -9.4817172050168489e-12, 
    -9.4458228147912893e-12, -9.42333915344512e-12, -9.4162206703346691e-12, 
    -9.4255402577522034e-12, -9.4513761995323294e-12, 
    -9.4927226702940611e-12, -9.5475059426394255e-12, 
    -9.6126701702064857e-12, -9.6843229630116287e-12, 
    -9.7579151509894604e-12, -9.8284682782929012e-12, 
    -9.8908270081908426e-12, -9.9399230626336499e-12, 
    -9.9710275782309448e-12, -9.9799941605191271e-12, 
    -9.9634976775163294e-12, -9.9192484144429924e-12, -9.846124284103607e-12, 
    -9.7443236230698248e-12, -9.6154123445572625e-12, 
    -9.4623505075677157e-12, -9.2894222100633552e-12, -9.102132942492578e-12, 
    -8.9070044143767618e-12, -8.7113351808511598e-12, -8.522866196448468e-12, 
    -8.3494308749806671e-12, -8.1985544722129068e-12, 
    -8.0770273564023707e-12, -7.9905161609194048e-12, 
    -7.9432009601735154e-12, -7.9374420297345844e-12, -7.973582217404091e-12, 
    -8.049829292822548e-12, -8.1622803162556956e-12, -8.3050613929646017e-12, 
    -8.4706585060762375e-12, -8.6502765515110007e-12, 
    -8.8343516139264418e-12, -9.0131227692352348e-12, 
    -9.1772055611010806e-12, -9.3181362111758902e-12, 
    -9.4288690263570809e-12, -9.5041479097595095e-12, 
    -9.5407698441680991e-12, -9.5377067678680572e-12, 
    -9.4960674404161345e-12, -9.4189423439344752e-12, 
    -9.3111396814535315e-12, -9.1788319892610214e-12, 
    -9.0291596793117263e-12, -8.8697864713326393e-12, 
    -8.7084720100646118e-12, -8.5526894105165082e-12, 
    -8.4092336817054825e-12, -8.2839105736295547e-12, 
    -8.1812782229419066e-12, -8.1044590596472381e-12, 
    -8.0550153324893868e-12, -8.0329051267179568e-12, 
    -8.0365423504418111e-12, -8.0629091200174056e-12, 
    -8.1077645332051595e-12, -8.1659430931443255e-12, 
    -8.2316900951677079e-12, -8.2990338587203604e-12, 
    -8.3621866222647629e-12, -8.4158947387940101e-12, 
    -8.4557620940618533e-12, -8.4784833980742617e-12, 
    -8.4819803404259745e-12, -8.4654437270121007e-12, 
    -8.4292758768836791e-12, -8.3749225822511088e-12, 
    -8.3046615338677509e-12, -8.2213424325518993e-12, 
    -8.1281259955742971e-12, -8.0282198965821077e-12, 
    -7.9246897477576778e-12, -7.8202975872030788e-12, 
    -7.7174593908198209e-12, -7.6182027176641705e-12, 
    -7.5242506161569973e-12, -7.4371017123898146e-12, 
    -7.3581461814152068e-12, -7.2887848794898042e-12, 
    -7.2305217291495002e-12, -7.1849826688030111e-12, 
    -7.1539149721297218e-12, -7.1390894820629715e-12, 
    -7.1421656959310255e-12, -7.1644759494879064e-12, 
    -7.2068238348401652e-12, -7.2692420856304961e-12, -7.350796432966222e-12, 
    -7.4494460795265295e-12, -7.5619983169202308e-12, 
    -7.6841442093227318e-12, -7.8106379386482385e-12, -7.935550209256457e-12, 
    -8.0526354337930181e-12, -8.155745640838098e-12, -8.2392859193975277e-12, 
    -8.2986049613950307e-12, -8.3303630363809896e-12, 
    -8.3327767558506506e-12, -8.3057413842731273e-12, 
    -8.2507905846568221e-12, -8.1709528096979899e-12, 
    -8.0704295342539225e-12, -7.9542422592123011e-12, 
    -7.8277737204184651e-12, -7.6963425735393842e-12, 
    -7.5647738939544605e-12, -7.4370887324654822e-12, 
    -7.3162494882850612e-12, -7.2040512974374269e-12, 
    -7.1011042591245818e-12, -7.0069432876005238e-12, 
    -6.9201990813781956e-12, -6.8388426988054348e-12, 
    -6.7604546500442091e-12, -6.6824700855969809e-12, 
    -6.6024481957554444e-12, -6.5182706460330258e-12, -6.428300830927277e-12, 
    -6.3314782619800934e-12, -6.2274297183709214e-12, 
    -6.1164497889618157e-12, -5.9995459060701889e-12, 
    -5.8783586536658545e-12, -5.7551619601303115e-12, 
    -5.6327311851283628e-12, -5.5143022736552605e-12, 
    -5.4033833079662576e-12, -5.3036637307598951e-12, 
    -5.2187550872325612e-12, -5.1520736239485528e-12, 
    -5.1065478966111799e-12, -5.0844706508100716e-12, 
    -5.0872623887991199e-12, -5.1153641488108157e-12, 
    -5.1681140981916348e-12, -5.2437795682763564e-12, 
    -5.3395686846221438e-12, -5.4518406226954125e-12, 
    -5.5762785737947055e-12, -5.7081807837005253e-12, 
    -5.8427554473485309e-12, -5.9754100149970429e-12, 
    -6.1019974394120209e-12, -6.2190482554379714e-12, 
    -6.3238715276539034e-12, -6.4146265154843611e-12, 
    -6.4902646904039425e-12, -6.5504444715882716e-12, 
    -6.5953812566574182e-12, -6.62568535920219e-12, -6.6421799200187626e-12, 
    -6.6457945274421957e-12, -6.637435433618189e-12, -6.6179800880247343e-12, 
    -6.5882494314988963e-12, -6.5490764537279441e-12, 
    -6.5013445312945496e-12, -6.4460799955983562e-12, 
    -6.3844930221776659e-12, -6.3180103855367566e-12, 
    -6.2482495763558317e-12, -6.1769971116625689e-12, -6.106091410504812e-12, 
    -6.037361141598868e-12, -5.9724867545616626e-12, -5.9129147622604488e-12, 
    -5.8597470306252319e-12, -5.8137138301764887e-12, 
    -5.7751100653911748e-12, -5.7438160675492621e-12, 
    -5.7192962004274988e-12, -5.7006671681412601e-12, 
    -5.6867438875012972e-12, -5.6761155772640282e-12, -5.66721661834871e-12, 
    -5.6584252306807665e-12, -5.6481186130760671e-12, 
    -5.6347803919232932e-12, -5.6170586609897075e-12, -5.593834339697868e-12, 
    -5.5642614658576743e-12, -5.5277988166580896e-12, 
    -5.4841987378382515e-12, -5.4334998125527155e-12, 
    -5.3759766272762621e-12, -5.31207795204008e-12, -5.2423748891041867e-12, 
    -5.1675034980310742e-12, -5.0881388528848113e-12, -5.004981647907925e-12, 
    -4.9187633978524641e-12, -4.8303031314749088e-12, -4.740537444925375e-12, 
    -4.6505678355026367e-12, -4.5616703167046625e-12, -4.475294518499445e-12, 
    -4.3929928279560239e-12, -4.3163170372198376e-12, 
    -4.2466694954685744e-12, -4.1851419838212051e-12, 
    -4.1323460580232278e-12, -4.0882740810965758e-12, 
    -4.0522096771967154e-12, -4.0227089723581711e-12, 
    -3.9976883396196103e-12, -3.9745630644606343e-12, 
    -3.9504955742070263e-12, -3.9226848831304519e-12, 
    -3.8886638876650318e-12, -3.8466331715846512e-12, 
    -3.7957017711533899e-12, -3.7360677733239243e-12, 
    -3.6691012171625761e-12, -3.5973142807626622e-12, 
    -3.5242016338337623e-12, -3.4540139895233714e-12, 
    -3.3914030321384144e-12, -3.3410524897475087e-12, 
    -3.3073509117947463e-12, -3.2939667127305072e-12, 
    -3.3035864413597738e-12, -3.337711521218835e-12, -3.3965536177452094e-12, 
    -3.4790521229345064e-12, -3.5829837599179936e-12, 
    -3.7051828924519477e-12, -3.8418043130802063e-12, 
    -3.9886438783511604e-12, -4.1414716651108654e-12, 
    -4.2963138202684159e-12, -4.4497088255561099e-12, 
    -4.5989097980573984e-12, -4.7419724096179602e-12, 
    -4.8777828487872949e-12, -5.0060134495887482e-12, -5.126985641516468e-12, 
    -5.241501426647076e-12, -5.3506480259596318e-12, -5.4555667166604463e-12, 
    -5.5572734114597297e-12, -5.6564586855160384e-12, 
    -5.7533696816033048e-12, -5.8477198941749941e-12, 
    -5.9386633124326498e-12, -6.0248100718279911e-12, 
    -6.1043121454866319e-12, -6.1749678024057343e-12, -6.234371981281596e-12, 
    -6.2800697484436691e-12, -6.3097422394592134e-12, -6.321364572143435e-12, 
    -6.3133608954194803e-12, -6.2847401320880551e-12, 
    -6.2351951577664056e-12, -6.1651748531936761e-12, 
    -6.0759228054687611e-12, -5.969463707000497e-12, -5.8485768167025605e-12, 
    -5.7167231901617894e-12, -5.5779179880960973e-12, 
    -5.4366199827034174e-12, -5.297547762887491e-12, -5.1654945386379435e-12, 
    -5.0451368361238185e-12, -4.9408179029527463e-12, 
    -4.8563461617957496e-12, -4.7948080611617308e-12, 
    -4.7584105836117774e-12, -4.7483570011712519e-12, 
    -4.7647997245953187e-12, -4.8068255310246289e-12, 
    -4.8725351162421273e-12, -4.9591526856833028e-12, 
    -5.0632228791597321e-12, -5.1808157260224058e-12, 
    -5.3077613369683882e-12, -5.4398776344631795e-12, 
    -5.5731674147961345e-12, -5.703964326990583e-12, -5.8290366999501427e-12, 
    -5.94562220491151e-12, -6.0514039368196941e-12, -6.1444431235481569e-12, 
    -6.2230891411954655e-12, -6.2858843538538175e-12, 
    -6.3314794838968236e-12, -6.3585782315175414e-12, 
    -6.3659407647487384e-12, -6.3524196466800552e-12, 
    -6.3170470741917544e-12, -6.2591641890711009e-12, 
    -6.1785483134973714e-12, -6.0755515523076675e-12, -5.951210395811299e-12, 
    -5.8073143442255171e-12, -5.6464100279333666e-12, 
    -5.4717570462308954e-12, -5.287192741054949e-12, -5.0969651426140686e-12, 
    -4.9055102243489841e-12, -4.7172047619651066e-12, 
    -4.5361138489960285e-12, -4.3657544724742721e-12, -4.208906074905801e-12, 
    -4.0674371949863459e-12, -3.942256708130714e-12, -3.8332978055520437e-12, 
    -3.7395582997962172e-12, -3.6592332778795209e-12, 
    -3.5899253101163425e-12, -3.5288739743283079e-12, -3.473203184415345e-12, 
    -3.4201944866980463e-12, -3.3675653918519815e-12, 
    -3.3136527280259399e-12, -3.2575816294686046e-12, 
    -3.1993538820513499e-12, -3.1398137911381228e-12, 
    -3.0805577730812022e-12, -3.0237583219329579e-12, 
    -2.9719054436860809e-12, -2.9275205088144192e-12, 
    -2.8928447290882117e-12, -2.8695839298214195e-12, 
    -2.8586780344862153e-12, -2.8601729838510507e-12, 
    -2.8731763952497494e-12, -2.8959429842938588e-12, 
    -2.9260337656283074e-12, -2.9605745659441195e-12, 
    -2.9965410824418947e-12, -3.0310898596621021e-12, 
    -3.0618320024581462e-12, -3.0870940401808013e-12, 
    -3.1060788081711346e-12, -3.1189345281289271e-12, 
    -3.1267097634369904e-12, -3.1312849558950105e-12, 
    -3.1351392849311465e-12, -3.1411525705154687e-12, 
    -3.1523177037151213e-12, -3.1715117173368141e-12, 
    -3.2012549315326108e-12, -3.243544249161357e-12, -3.2997182602611389e-12, 
    -3.3704054782667412e-12, -3.4555045014702434e-12, 
    -3.5542120742793654e-12, -3.6650709109696387e-12, 
    -3.7860532134133349e-12, -3.9146265450715806e-12, 
    -4.0478191907402175e-12, -4.1822750895899912e-12, 
    -4.3143063209140326e-12, -4.4399536893108405e-12, 
    -4.5550465214080216e-12, -4.6552855219736021e-12, 
    -4.7363794440633443e-12, -4.794201878884177e-12, -4.8249662563822445e-12, 
    -4.8254598461351834e-12, -4.7932585876882576e-12, 
    -4.7269422903774784e-12, -4.626285042212032e-12, -4.492376717329513e-12, 
    -4.3276826789103674e-12, -4.1360116739479479e-12, 
    -3.9223987992833131e-12, -3.6929173737278201e-12, 
    -3.4543955930568642e-12, -3.2140976731995865e-12, 
    -2.9793825868828203e-12, -2.7573273752338773e-12, 
    -2.5544114855593913e-12, -2.3762003458410454e-12, 
    -2.2271197022557071e-12, -2.1102468145439447e-12, 
    -2.0272600241995719e-12, -1.9783859212256707e-12, 
    -1.9624506325821874e-12, -1.9769780576837466e-12, 
    -2.0183965578264703e-12, -2.0822326677993884e-12, 
    -2.1633756889093529e-12, -2.2563497227237108e-12, 
    -2.3556309584823905e-12, -2.455897317737757e-12, -2.5523350423566326e-12, 
    -2.6408543170839458e-12, -2.7183168433262065e-12, 
    -2.7826408799277032e-12, -2.8329259249389177e-12, 
    -2.8694054429016717e-12, -2.8934381562976455e-12, 
    -2.9073275532756426e-12, -2.9141667153142833e-12, 
    -2.9175536889916994e-12, -2.9213770916652794e-12, 
    -2.9294817202151385e-12, -2.9454542903400949e-12, 
    -2.9723463868576154e-12, -3.0125168747813658e-12, 
    -3.0674775683978874e-12, -3.1378393645138063e-12, 
    -3.2233017157359568e-12, -3.322710343696947e-12, -3.4341391599815796e-12, 
    -3.5550339160152436e-12, -3.6823623196060463e-12, 
    -3.8127576512095504e-12, -3.9426753021867671e-12, 
    -4.0685304580127686e-12, -4.186824942016042e-12, -4.2942381154821959e-12, 
    -4.3877465706066614e-12, -4.4646573067516034e-12, 
    -4.5227360125665516e-12, -4.5602182341474074e-12, 
    -4.5759185020197865e-12, -4.5692462564161383e-12, 
    -4.5403030920018486e-12, -4.4898552431348388e-12, 
    -4.4193951348136707e-12, -4.3310807341762439e-12, 
    -4.2277102431174269e-12, -4.1125895045818872e-12, 
    -3.9894351238386748e-12, -3.8621624014856224e-12, 
    -3.7347455616381064e-12, -3.6109409149261677e-12, 
    -3.4941421277662522e-12, -3.3871550794739213e-12, 
    -3.2920640212474377e-12, -3.2101076812832936e-12, 
    -3.1416610881753295e-12, -3.0862155077714911e-12, 
    -3.0424785616602099e-12, -3.0085002802955466e-12, 
    -2.9818438952291574e-12, -2.9598014405152951e-12, 
    -2.9396233915867964e-12, -2.9187171547098039e-12, 
    -2.8948549932712581e-12, -2.8663280196867613e-12, 
    -2.8320487918566645e-12, -2.7916114769085631e-12, 
    -2.7452788817127637e-12, -2.693907356191946e-12, -2.6388326487773651e-12, 
    -2.5817015523279713e-12, -2.524287605553545e-12, -2.4682906309285365e-12, 
    -2.4151524695440319e-12, -2.365886427782174e-12, -2.320959010483421e-12, 
    -2.2802256655407295e-12, -2.2429397332672663e-12, 
    -2.2077886683073639e-12, -2.1730094326588676e-12, 
    -2.1365823576326155e-12, -2.0964160121622047e-12, 
    -2.0505516320808213e-12, -1.9973955534269804e-12, 
    -1.9358829969020973e-12, -1.8656449611131939e-12, 
    -1.7870842695026113e-12, -1.7014225491750672e-12, 
    -1.6106498591966348e-12, -1.5174441663865217e-12, -1.425011458146724e-12, 
    -1.3369099756120345e-12, -1.2568234833758619e-12, 
    -1.1883534169399045e-12, -1.1347784566703984e-12, 
    -1.0988734102232168e-12, -1.0827422253451021e-12, 
    -1.0877068979951111e-12, -1.1142210860310269e-12, 
    -1.1619035837962451e-12, -1.2295305821918167e-12, 
    -1.3151579007689636e-12, -1.4162708264141085e-12, 
    -1.5299483602232448e-12, -1.6530480146394008e-12, 
    -1.7824456641517984e-12, -1.9151857178766554e-12, 
    -2.0486805979257627e-12, -2.1808150046157909e-12, 
    -2.3100391235880435e-12, -2.435391187091139e-12, -2.5564812718367837e-12, 
    -2.6733982939222797e-12, -2.7866187421588433e-12, 
    -2.8968570016250429e-12, -3.004919692083293e-12, -3.1115899004958326e-12, 
    -3.2174971546929643e-12, -3.3230354638933891e-12, 
    -3.4283269323688602e-12, -3.533179220132318e-12, -3.6370923407912082e-12, 
    -3.7392973006582424e-12, -3.8387661638669455e-12, 
    -3.9342355458449048e-12, -4.0242483002990647e-12, 
    -4.1071349346053769e-12, -4.1810204560435647e-12, 
    -4.2438505446983485e-12, -4.2933858456694778e-12, 
    -4.3272443116500062e-12, -4.3429541233217028e-12, 
    -4.3380417800213565e-12, -4.3101462258864965e-12, 
    -4.2571569794447349e-12, -4.177358110195247e-12, -4.0695824578673107e-12, 
    -3.9333339576391277e-12, -3.7689053762736959e-12, 
    -3.5774370850700577e-12, -3.3609359038916688e-12, 
    -3.1222495330007785e-12, -2.8650068537179417e-12, 
    -2.5934953660854018e-12, -2.3125394559691864e-12, 
    -2.0273465581348757e-12, -1.7433530862995929e-12, 
    -1.4660709287002226e-12, -1.200958619428882e-12, -9.5329846236381237e-13, 
    -7.2807409699546473e-13, -5.2989365400905419e-13, 
    -3.6289707821868056e-13, -2.3070288936052142e-13, -1.363138938010777e-13, 
    -8.2066682227070205e-14, -6.9566831166777157e-14, 
    -9.9628179272201675e-14, -1.7222419500167976e-13, 
    -2.8646339379040014e-13, -4.405648575823255e-13, -6.3187367801462361e-13, 
    -8.5691070055029627e-13, -1.111444490695212e-12, -1.3905970744159227e-12, 
    -1.6889813521163987e-12, -2.0008433810551161e-12, 
    -2.3202432147662536e-12, -2.6411980862582216e-12, 
    -2.9578506402688323e-12, -3.2646043831771846e-12, 
    -3.5562402161024115e-12, -3.8280226425762232e-12, -4.075748265101267e-12, 
    -4.2958091739705543e-12, -4.4852280835226434e-12, -4.641664927343802e-12, 
    -4.7634397730336681e-12, -4.8495373974810784e-12, 
    -4.8996136251489269e-12, -4.9140114645812616e-12, 
    -4.8937649531831008e-12, -4.8405915621067812e-12, 
    -4.7568962685650049e-12, -4.6457220122134668e-12, 
    -4.5107156188690071e-12, -4.3560335481803339e-12, 
    -4.1862337538235674e-12, -4.0061281740371304e-12, -3.820594248984967e-12, 
    -3.6344128588206373e-12, -3.4520373513803697e-12, 
    -3.2774213227264338e-12, -3.1138368399870887e-12, 
    -2.9637459061656543e-12, -2.8287301258993637e-12, 
    -2.7094684545011898e-12, -2.6057875920290301e-12, 
    -2.5167925385871064e-12, -2.4410470028649589e-12, 
    -2.3767608765657638e-12, -2.3220385733949292e-12, 
    -2.2751110518801022e-12, -2.2345312228515277e-12, 
    -2.1993194036564824e-12, -2.1690624171720819e-12, 
    -2.1439078061764953e-12, -2.1245011114880135e-12, 
    -2.1118419140827918e-12, -2.1070837930931995e-12, 
    -2.1112959993262018e-12, -2.1252448416391761e-12, 
    -2.1491234477097829e-12, -2.1823972688753202e-12, 
    -2.2236951001799085e-12, -2.2707957168708146e-12, 
    -2.3206856601219206e-12, -2.3697623285369875e-12, 
    -2.4140699907417281e-12, -2.4496523403523566e-12, 
    -2.4728960897328305e-12, -2.48087450750456e-12, -2.4716647978600445e-12, 
    -2.4445638072545747e-12, -2.4001968602659104e-12, 
    -2.3404959884320351e-12, -2.2685437406250408e-12, 
    -2.1882957848542158e-12, -2.104188410928657e-12, -2.0207182278477091e-12, 
    -1.9419911975462723e-12, -1.871323110991132e-12, -1.8109412424124777e-12, 
    -1.7617963977841657e-12, -1.7235586309363364e-12, 
    -1.6947521279507821e-12, -1.6730412764398757e-12, 
    -1.6556199801796355e-12, -1.639671437496663e-12, -1.6228215605284508e-12, 
    -1.6035424285835074e-12, -1.5814406256477563e-12, 
    -1.5573858661168837e-12, -1.5334788173725671e-12, 
    -1.5128471422916898e-12, -1.4992839142700745e-12, 
    -1.4967854344049183e-12, -1.5090356623709614e-12, 
    -1.5388883771073791e-12, -1.5879533307691611e-12, 
    -1.6562691082424627e-12, -1.7421753674968835e-12, 
    -1.8423390417474099e-12, -1.9519912215164471e-12, 
    -2.0652786324383278e-12, -2.1757596193805039e-12, -2.27693881133122e-12, 
    -2.3628132764779956e-12, -2.4283425973468186e-12, 
    -2.4698388298229247e-12, -2.4851909844438645e-12, 
    -2.4739876996084309e-12, -2.4374200704899197e-12, 
    -2.3780979398933774e-12, -2.2997910575222808e-12, 
    -2.2070569237736267e-12, -2.1048655089236308e-12, 
    -1.9982524647670384e-12, -1.8919850341576397e-12, 
    -1.7903216918308367e-12, -1.6968211618522914e-12, 
    -1.6142455684731362e-12, -1.5445209957270327e-12, 
    -1.4887592235608164e-12, -1.4473356321875467e-12, 
    -1.4199984829347191e-12, -1.4059741426448854e-12, 
    -1.4041293694438876e-12, -1.4130757322612619e-12, -1.431312782518698e-12, 
    -1.4573245323345098e-12, -1.4896747047804322e-12, 
    -1.5270817301203637e-12, -1.5684821561012501e-12, 
    -1.6130532063681823e-12, -1.660221057809022e-12, -1.7096822280803276e-12, 
    -1.7614023312600922e-12, -1.8155699150493972e-12, 
    -1.8725789070035479e-12, -1.9329988902151619e-12, 
    -1.9975322745885653e-12, -2.0669442051004979e-12, 
    -2.1420035808958373e-12, -2.2233948004644763e-12, 
    -2.3116262570116213e-12, -2.4069243132705099e-12, 
    -2.5091263898247469e-12, -2.6175776993152315e-12, 
    -2.7310534045531003e-12, -2.8476950892032364e-12, 
    -2.9650004131199151e-12, -3.0798611173378171e-12, 
    -3.1886644427222243e-12, -3.2874178626400647e-12, 
    -3.3719560052678842e-12, -3.438182776185575e-12, -3.482299635594808e-12, 
    -3.5010797740231253e-12, -3.492084772632106e-12, -3.4538617931687263e-12, 
    -3.3860740591820589e-12, -3.2895739756569692e-12, 
    -3.1663980772979166e-12, -3.0196945251461575e-12, 
    -2.8535911165698736e-12, -2.673019370322449e-12, -2.4834593266765424e-12, 
    -2.2907434872227143e-12, -2.100791247550559e-12, -1.919355120038084e-12, 
    -1.7518074753440633e-12, -1.6029373649990909e-12, 
    -1.4767859542695587e-12, -1.3765052775783703e-12, 
    -1.3042478119255148e-12, -1.2611162754913445e-12, 
    -1.2471265447091712e-12, -1.2612237373930151e-12, 
    -1.3013454799736671e-12, -1.3645139731348986e-12, 
    -1.4469717991510632e-12, -1.5443709884004147e-12, 
    -1.6519754149384644e-12, -1.7648796737535156e-12, -1.878252558245169e-12, 
    -1.9875536623573942e-12, -2.0887291895705789e-12, 
    -2.1783716957004116e-12, -2.2538558008583706e-12, 
    -2.3133485314090709e-12, -2.3558475477424542e-12, 
    -2.3810963366710587e-12, -2.3895118621925807e-12, 
    -2.3820426637602619e-12, -2.3600351310411259e-12, 
    -2.3250924528472667e-12, -2.2789651799061613e-12, 
    -2.2234502408424413e-12, -2.1603399305659897e-12, 
    -2.0913868599199682e-12, -2.0183046750616204e-12, 
    -1.9427981848757852e-12, -1.8665825306423276e-12, 
    -1.7914166800969154e-12, -1.719108123218557e-12, -1.651522018933917e-12, 
    -1.5905436214428195e-12, -1.5380318992329438e-12, 
    -1.4957566973584639e-12, -1.4653132390899595e-12, 
    -1.4480369162038795e-12, -1.4449262141594372e-12, 
    -1.4565804652367635e-12, -1.4831282458930638e-12, 
    -1.5242092800006552e-12, -1.578978016519992e-12, -1.6461212188993666e-12, 
    -1.7239142929846511e-12, -1.8102978896561225e-12, 
    -1.9029916785018416e-12, -1.9995900962254428e-12, 
    -2.0977153646850806e-12, -2.1951040960962549e-12, -2.289733367400685e-12, 
    -2.3798703728914139e-12, -2.4641300245223754e-12, 
    -2.5414603297057252e-12, -2.6110955911954503e-12, 
    -2.6724828064966789e-12, -2.7251771287952426e-12, 
    -2.7687532881398547e-12, -2.802706803807119e-12, -2.8263961557763048e-12, 
    -2.8390647721466346e-12, -2.8398861217881551e-12, 
    -2.8280664073026288e-12, -2.8030188924070572e-12, 
    -2.7645361802034266e-12, -2.7129832587121977e-12, 
    -2.6494619541564043e-12, -2.5759134991169743e-12, 
    -2.4951518602235018e-12, -2.4108282550546987e-12, 
    -2.3272363013457711e-12, -2.2490904752391824e-12, 
    -2.1812128088066311e-12, -2.1281689462989052e-12, 
    -2.0938853019214919e-12, -2.081314952198914e-12, -2.0921290417060467e-12, 
    -2.1265155151075927e-12, -2.1830811134340576e-12, -2.258865825088056e-12, 
    -2.349478935924397e-12, -2.4493483198203991e-12, -2.5520439984296037e-12, 
    -2.6506670053701098e-12, -2.7382752466542281e-12, 
    -2.8082989846264237e-12, -2.8549043220095607e-12, 
    -2.8733413984938547e-12, -2.860167948370234e-12, -2.8134474074723466e-12, 
    -2.7328001417871227e-12, -2.6194163750000122e-12, 
    -2.4759806084030076e-12, -2.3065399763831538e-12, 
    -2.1163050911043473e-12, -1.9114395097495371e-12, 
    -1.6987890623581619e-12, -1.4856338999456999e-12, 
    -1.2793547401989202e-12, -1.0872065864499645e-12, 
    -9.1596229617325688e-13, -7.7165860723307131e-13, 
    -6.5936103320841919e-13, -5.8293964949635206e-13, 
    -5.4488806582769763e-13, -5.4622794444771757e-13, 
    -5.8645046225633205e-13, -6.6355760873218048e-13, 
    -7.7414244506144788e-13, -9.1356968430633758e-13, 
    -1.0761688425197241e-12, -1.2555387182481815e-12, 
    -1.4448054884418154e-12, -1.6369593192958586e-12, 
    -1.8251576146678204e-12, -2.0030265142211001e-12, 
    -2.1649076257230497e-12, -2.3060927205802119e-12, 
    -2.4229552984006395e-12, -2.5130582685206967e-12, 
    -2.5751716741175675e-12, -2.6092295439760264e-12, 
    -2.6162218039499055e-12, -2.5980489552719751e-12, 
    -2.5573104315777467e-12, -2.4971051753888243e-12, 
    -2.4207987931863263e-12, -2.3318199748321163e-12, 
    -2.2334709542703768e-12, -2.1287803574016553e-12, 
    -2.0203920532568795e-12, -1.9105138416226798e-12, -1.8008847187154e-12, 
    -1.6928178035337673e-12, -1.5872392257065366e-12, -1.484750950637849e-12, 
    -1.3857403006449881e-12, -1.290460464532735e-12, -1.1991070227672558e-12, 
    -1.1118995972913748e-12, -1.0291402206059624e-12, 
    -9.5127214203333151e-13, -8.7892029341921088e-13, 
    -8.1290440666943421e-13, -7.5428755061406933e-13, -7.043621292137932e-13, 
    -6.6467386186337521e-13, -6.3698607479190597e-13, 
    -6.2325512973179261e-13, -6.2556143728203148e-13, 
    -6.4600637391683891e-13, -6.8657616641515903e-13, 
    -7.4898390784074762e-13, -8.3446962836260063e-13, 
    -9.4360095409148157e-13, -1.0760661225435507e-12, 
    -1.2305251675624722e-12, -1.4044835396817506e-12, 
    -1.5942556680377804e-12, -1.7950087860285462e-12, 
    -2.0009271008759891e-12, -2.2054455523826553e-12, 
    -2.4015978738754926e-12, -2.5824116153626219e-12, 
    -2.7413589677736534e-12, -2.8728029991326213e-12, 
    -2.9724013259750001e-12, -3.0374563826466294e-12, 
    -3.0671525364638732e-12, -3.0626634134525422e-12, 
    -3.0271361095805898e-12, -2.9655166591776365e-12, 
    -2.8842417917381274e-12, -2.7908345932634697e-12, 
    -2.6933902600681357e-12, -2.6000388127073525e-12, 
    -2.5183756204564955e-12, -2.4549441804030893e-12, 
    -2.4147750389331408e-12, -2.4010323910662701e-12,
  // Sqw-F(1, 0-1999)
    0.11657913759996912, 0.11607557541154639, 0.11458146934983199, 
    0.11214557078821014, 0.10884591742533103, 0.10478530219515197, 
    0.10008547763039144, 0.09488056969922927, 0.089310216504517578, 
    0.083512936078982442, 0.077620168518573632, 0.071751341056230752, 
    0.066010184275696757, 0.060482398897984686, 0.055234650158844843, 
    0.050314762914332248, 0.045752913638652977, 0.04156356942523156, 
    0.03774790875296323, 0.034296470400424758, 0.031191809307218543, 
    0.02841098400476675, 0.025927752027079285, 0.023714400910449303, 
    0.021743187956204016, 0.019987398616644531, 0.018422059703778061, 
    0.017024359673745579, 0.015773835202830246, 0.014652383031755251, 
    0.013644150774530713, 0.012735352156953372, 0.011914042748669328, 
    0.011169883021980411, 0.010493907377246271, 0.0098783110536559658, 
    0.0093162616868766243, 0.0088017385399296964, 0.0083293998542192122, 
    0.0078944770443102191, 0.0074926933248741518, 0.0071202036110016229, 
    0.0067735520512131921, 0.0064496432808726131, 0.006145723412662815, 
    0.005859366920192878, 0.0055884659268092204, 0.0053312189707526722, 
    0.005086117039862858, 0.0048519254895979117, 0.0046276612971187479, 
    0.0044125658785492154, 0.0042060743333263151, 0.0040077824267509398, 
    0.0038174128547556973, 0.003634782357748465, 0.0034597710929179667, 
    0.0032922953849550984, 0.0031322846115115011, 0.0029796625996563824, 
    0.0028343335625838867, 0.0026961723272750262, 0.0025650184122270156, 
    0.002440673411637844, 0.0023229011167681481, 0.0022114298357633387, 
    0.0021059564355011104, 0.0020061516999562534, 0.00191166666136009, 
    0.0018221396028469188, 0.0017372034519936616, 0.0016564932880717021, 
    0.0015796536806923279, 0.0015063455741957863, 0.0014362524398853042, 
    0.001369085443321713, 0.0013045874185976583, 0.0012425355039804521, 
    0.0011827423684296317, 0.001125056039155052, 0.0010693584188919047, 
    0.0010155626509444036, 0.00096360954487177946, 0.00091346331258703904, 
    0.00086510688229208339, 0.00081853705659791769, 0.0007737597632876005, 
    0.00073078561538581855, 0.00068962595501151098, 0.0006502895067482359, 
    0.00061277971489119294, 0.00057709278874482105, 0.00054321643465940071, 
    0.00051112921570284429, 0.00048080045198656485, 0.00045219055797253763, 
    0.0004252517077320002, 0.0003999287241325087, 0.00037616010128513404, 
    0.00035387908850260323, 0.0003330147852839851, 0.00031349321725120745, 
    0.00029523837974477644, 0.0002781732469896477, 0.00026222074946550378, 
    0.00024730472061816459, 0.00023335080763421797, 0.00022028733178803048, 
    0.00020804607438343144, 0.00019656295706173502, 0.00018577858227268997, 
    0.00017563860224316537, 0.0001660938930401086, 0.00015710052348312967, 
    0.00014861952498359092, 0.00014061648555569462, 0.00013306100673890934, 
    0.00012592607371084271, 0.00011918739476842297, 0.00011282276580621106, 
    0.00010681150858315278, 0.00010113401953223141, 9.5771450427931161e-05, 
    9.0705525590349502e-05, 8.5918484714014965e-05, 8.1393127809179471e-05, 
    7.7112930494005688e-05, 7.3062194607525813e-05, 6.9226200678681495e-05, 
    6.5591334375222663e-05, 6.2145167369338341e-05, 5.8876482578786593e-05, 
    5.5775242979452951e-05, 5.2832510910773579e-05, 5.0040330183012586e-05, 
    4.7391586001563837e-05, 4.4879857852868204e-05, 4.2499278520596148e-05, 
    4.0244409009789866e-05, 3.8110135122902734e-05, 3.6091587461959324e-05, 
    3.4184083283651483e-05, 3.2383086253897916e-05, 3.0684178873428913e-05, 
    2.9083042126426926e-05, 2.7575437562366554e-05, 2.6157188300132709e-05, 
    2.4824157067602473e-05, 2.3572221092183892e-05, 2.2397245217498484e-05, 
    2.1295055859001989e-05, 2.0261419209673385e-05, 1.9292027391875912e-05, 
    1.8382496009790764e-05, 1.7528375816355462e-05, 1.6725180053960894e-05, 
    1.5968427578349145e-05, 1.5253700290889294e-05, 1.4576711855929564e-05, 
    1.393338334477944e-05, 1.3319920474504878e-05, 1.2732886614219789e-05, 
    1.2169265770383099e-05, 1.1626510340110078e-05, 1.1102569479257633e-05, 
    1.0595895370499339e-05, 1.0105426356561383e-05, 9.6305476751381771e-06, 
    9.1710322354001207e-06, 8.7269653722373774e-06, 8.2986586783174054e-06, 
    7.8865587581540852e-06, 7.4911570145362749e-06, 7.1129063513988517e-06, 
    6.7521499791490899e-06, 6.409066403758947e-06, 6.0836332649127822e-06, 
    5.7756110911157834e-06, 5.4845464039120576e-06, 5.2097920827035807e-06, 
    4.9505416337171786e-06, 4.7058731074266989e-06, 4.4747979504785672e-06, 
    4.2563100883937445e-06, 4.0494309860230453e-06, 3.8532472526916317e-06, 
    3.6669384351682548e-06, 3.4897938433084778e-06, 3.3212184396636517e-06, 
    3.1607288720823538e-06, 3.0079415352663347e-06, 2.8625550532295902e-06, 
    2.7243297559630925e-06, 2.5930666013188021e-06, 2.4685876187509897e-06, 
    2.3507194046894953e-06, 2.23928056847162e-06, 2.134073405705387e-06, 
    2.0348795392042173e-06, 1.9414588761650061e-06, 1.8535510136852581e-06, 
    1.7708781861803453e-06, 1.6931489616204918e-06, 1.6200621142980313e-06, 
    1.5513103698509311e-06, 1.4865839748521619e-06, 1.425574234665679e-06, 
    1.3679772559206766e-06, 1.3134981092736448e-06, 1.2618555070789716e-06, 
    1.2127868990789795e-06, 1.1660536749241263e-06, 1.1214459743568165e-06, 
    1.0787864914643405e-06, 1.0379326489176095e-06, 9.9877662490032507e-07, 
    9.612429278967275e-07, 9.2528350395716029e-07, 8.9087068109486278e-07, 
    8.5798855699781558e-07, 8.2662366854570356e-07, 7.9675590970497597e-07, 
    7.6835066490337831e-07, 7.4135300013785745e-07, 7.1568451934910754e-07, 
    6.9124318579390185e-07, 6.6790606863350111e-07, 6.4553465135917471e-07, 
    6.2398207093812356e-07, 6.0310147676392414e-07, 5.8275462169967418e-07, 
    5.6281982718785313e-07, 5.4319858512193706e-07, 5.2382025020720718e-07, 
    5.0464450544319038e-07, 4.8566152138790841e-07, 4.6688994696403634e-07, 
    4.4837304721574069e-07, 4.3017342630300886e-07, 4.1236684125690515e-07, 
    3.95035624861757e-07, 3.7826220563369484e-07, 3.6212314922661425e-07, 
    3.4668406236630167e-07, 3.3199560595663366e-07, 3.1809076874217979e-07, 
    3.0498345928843454e-07, 2.9266838910055347e-07, 2.8112214242922834e-07, 
    2.7030526468582475e-07, 2.6016515081769915e-07, 2.5063948273412192e-07, 
    2.4165995059061007e-07, 2.3315599936339225e-07, 2.2505836605127361e-07, 
    2.173022132101061e-07, 2.098297134350697e-07, 2.0259199333062496e-07, 
    1.9555039572658137e-07, 1.8867706322081239e-07, 1.8195487927652701e-07, 
    1.7537682716985714e-07, 1.6894484191432878e-07, 1.6266824073934158e-07, 
    1.5656182559066177e-07, 1.506437605830066e-07, 1.4493333763281701e-07, 
    1.3944875492659023e-07, 1.3420504140583108e-07, 1.2921226343861423e-07, 
    1.2447414211710666e-07, 1.199871900540374e-07, 1.1574044277152596e-07, 
    1.1171581497339407e-07, 1.0788905851640033e-07, 1.0423124436121854e-07, 
    1.0071063985002608e-07, 9.7294813971266511e-08, 9.3952780380627387e-08, 
    9.0656985538389177e-08, 8.7384966911464593e-08, 8.4120542694126833e-08, 
    8.085444445420461e-08, 7.7584362438535775e-08, 7.431443154790644e-08, 
    7.1054239309198236e-08, 6.781747743767688e-08, 6.4620384665985672e-08, 
    6.1480136041259553e-08, 5.8413325714771766e-08, 5.5434667164730726e-08, 
    5.2556002021838791e-08, 4.9785669709863482e-08, 4.7128251089855857e-08, 
    4.4584662828581813e-08, 4.215255044828628e-08, 3.9826907127823006e-08, 
    3.7600835206256881e-08, 3.5466365828019998e-08, 3.3415259858063386e-08, 
    3.143972647850187e-08, 2.9533014019562965e-08, 2.7689846482208831e-08, 
    2.5906698086292717e-08, 2.4181913139766412e-08, 2.2515690156269438e-08, 
    2.0909954672143591e-08, 1.9368146575536523e-08, 1.7894944408447398e-08, 
    1.6495944051266345e-08, 1.5177302707384886e-08, 1.3945354966995412e-08, 
    1.2806205376094561e-08, 1.1765304196330462e-08, 1.0827017504331739e-08, 
    9.9942105579241654e-09, 9.2678704662288517e-09, 8.6468005361442794e-09, 
    8.1274202508171383e-09, 7.703702306518142e-09, 7.3672688190490691e-09, 
    7.1076559944410371e-09, 6.912738978037501e-09, 6.7692916630002886e-09, 
    6.6636398408412448e-09, 6.5823552278770418e-09, 6.5129320172662207e-09, 
    6.4443895290467886e-09, 6.3677521768764893e-09, 6.2763718152816246e-09, 
    6.1660736665445601e-09, 6.0351251604182556e-09, 5.8840429196772739e-09, 
    5.7152669908661957e-09, 5.5327398473398604e-09, 5.3414324101343209e-09, 
    5.1468583366241032e-09, 4.9546138646649102e-09, 4.7699725782140804e-09, 
    4.597555791663763e-09, 4.441089237734198e-09, 4.3032481627267025e-09, 
    4.1855849478876308e-09, 4.0885285643311205e-09, 4.0114415762109734e-09, 
    3.9527203102218051e-09, 3.9099245920526024e-09, 3.8799266199324501e-09, 
    3.859071363023242e-09, 3.8433443387872382e-09, 3.8285443926168913e-09, 
    3.8104603280570037e-09, 3.7850490488374965e-09, 3.7486114071181137e-09, 
    3.6979588291812358e-09, 3.630561462554154e-09, 3.5446665106981052e-09, 
    3.4393754739530209e-09, 3.3146702334578351e-09, 3.1713821142138334e-09, 
    3.0111027485690811e-09, 2.8360421191686161e-09, 2.6488448570217146e-09, 
    2.4523811487228316e-09, 2.2495314520029312e-09, 2.0429852216473045e-09, 
    1.8350718051259472e-09, 1.627637934200643e-09, 1.4219803385797528e-09, 
    1.2188360950059393e-09, 1.0184268189354118e-09, 8.2054804567737417e-10, 
    6.2469130846768192e-10, 4.301848850383497e-10, 2.363388789789644e-10, 
    4.2582006825453541e-11, -1.514205677767006e-10, -3.4567602359329408e-10, 
    -5.3980436483270804e-10, -7.3301317218906772e-10, 
    -9.2410715778765426e-10, -1.1115313419052287e-09, 
    -1.2934452287257803e-09, -1.4678238271996327e-09, 
    -1.6325800127569353e-09, -1.7857009343970925e-09, 
    -1.9253898458884715e-09, -2.0502031950513316e-09, -2.159172232179182e-09, 
    -2.2518982467117448e-09, -2.3286118375423763e-09, 
    -2.3901885146428595e-09, -2.438116468905794e-09, -2.4744161095977272e-09, 
    -2.5015156549396477e-09, -2.5220911057655596e-09, -2.538883038577953e-09, 
    -2.5545049152166612e-09, -2.5712591922212574e-09, 
    -2.5909769655060307e-09, -2.6148951500997901e-09, 
    -2.6435815728211159e-09, -2.6769144792437693e-09, 
    -2.7141175571299881e-09, -2.7538470564339426e-09, 
    -2.7943226833851923e-09, -2.8334905688374288e-09, 
    -2.8692038999723039e-09, -2.8994057895362578e-09, 
    -2.9222991945279954e-09, -2.9364904248317963e-09, 
    -2.9410954087166071e-09, -2.9358016105716977e-09, 
    -2.9208824850830752e-09, -2.8971655553867946e-09, 
    -2.8659589162182093e-09, -2.8289442132050133e-09, 
    -2.7880463622267202e-09, -2.7452915317906311e-09, -2.702664835953695e-09, 
    -2.6619785770413427e-09, -2.6247598847281824e-09, 
    -2.5921644754850402e-09, -2.5649205913945854e-09, -2.543304582495722e-09, 
    -2.5271470906099013e-09, -2.5158669413355471e-09, 
    -2.5085280376570926e-09, -2.503913862631253e-09, -2.5006133999942999e-09, 
    -2.4971126038307539e-09, -2.4918856229133563e-09, 
    -2.4834808828009998e-09, -2.4705978038170682e-09, 
    -2.4521510156876354e-09, -2.4273196277800847e-09, 
    -2.3955803406103526e-09, -2.3567236126720315e-09, 
    -2.3108532160544705e-09, -2.2583698279296647e-09, 
    -2.1999402424279409e-09, -2.1364540478235373e-09, 
    -2.0689704945569211e-09, -1.9986584357296117e-09, 
    -1.9267329457489535e-09, -1.8543922930343037e-09, 
    -1.7827591412440675e-09, -1.7128295983183845e-09, 
    -1.6454332708131709e-09, -1.5812067047535865e-09, 
    -1.5205816033111747e-09, -1.4637878874342568e-09, 
    -1.4108706751626567e-09, -1.3617187893020969e-09, 
    -1.3161018666538426e-09, -1.2737121898413645e-09, 
    -1.2342075244849122e-09, -1.1972511010643173e-09, 
    -1.1625457677512012e-09, -1.1298598015830973e-09, 
    -1.0990431422069744e-09, -1.0700334847288504e-09, 
    -1.0428528021892566e-09, -1.0175953402871872e-09, 
    -9.9440885836233456e-10, -9.7347101600016912e-10, 
    -9.5496304278008815e-10, -9.3904268975689543e-10, -9.258184723543555e-10, 
    -9.1532688916251632e-10, -9.0751424842274877e-10, 
    -9.0222429515864519e-10, -8.9919275876682639e-10, 
    -8.9804934095982902e-10, -8.9832752689008451e-10, 
    -8.9948184682059985e-10, -9.0091199207511235e-10, 
    -9.0199241346269756e-10, -9.0210589265719477e-10, 
    -9.0067886484139737e-10, -8.9721644991150298e-10, 
    -8.9133469025553984e-10, -8.8278792054861922e-10, 
    -8.7148914716909398e-10, -8.575219262812048e-10, -8.411424118393661e-10, 
    -8.2277109384106667e-10, -8.0297408823687237e-10, 
    -7.8243469975590904e-10, -7.619165123738223e-10, -7.4222015054480979e-10, 
    -7.2413610081673119e-10, -7.0839685320259154e-10, -6.956315587318788e-10, 
    -6.8632661871226795e-10, -6.8079516020577732e-10, 
    -6.7915795525477654e-10, -6.8133726242330847e-10, 
    -6.8706423049601878e-10, -6.9589924536632075e-10, 
    -7.0726357626803779e-10, -7.2047972326901424e-10, 
    -7.3481720974014393e-10, -7.4954010138904967e-10, 
    -7.6395265806227606e-10, -7.7743964805048972e-10, 
    -7.8949855320464231e-10, -7.9976160760968819e-10, -8.08006554326732e-10, 
    -8.1415592762903057e-10, -8.182656170495716e-10, -8.2050422964128603e-10, 
    -8.211254657881839e-10, -8.2043611546707629e-10, -8.1876255026229862e-10, 
    -8.1641854373457981e-10, -8.1367701577345851e-10, -8.107478581279298e-10, 
    -8.0776336410205513e-10, -8.0477211910284698e-10, 
    -8.0174136932899384e-10, -7.9856720374689295e-10, 
    -7.9509121491252309e-10, -7.9112179862066651e-10, 
    -7.8645794172296098e-10, -7.8091328900753435e-10, 
    -7.7433827197899775e-10, -7.6663851975133914e-10, 
    -7.5778812631391721e-10, -7.4783684159432473e-10, 
    -7.3691087922123384e-10, -7.2520758943403851e-10, 
    -7.1298467171676991e-10, -7.0054502394273216e-10, 
    -6.8821859574582944e-10, -6.7634272385428485e-10, -6.652424562584289e-10, 
    -6.5521222381074759e-10, -6.4650006261643602e-10, 
    -6.3929526799936544e-10, -6.3372011324903716e-10, 
    -6.2982588570019242e-10, -6.2759323955912417e-10, 
    -6.2693661252974372e-10, -6.2771219168859268e-10, 
    -6.2972877057588165e-10, -6.3276080504240258e-10, 
    -6.3656273236270481e-10, -6.40883756755904e-10, -6.4548224269023731e-10, 
    -6.5013887650940593e-10, -6.5466780775654188e-10, -6.589251965007476e-10, 
    -6.628145425133287e-10, -6.6628856638061273e-10, -6.6934745163879915e-10, 
    -6.7203364713060509e-10, -6.7442354743864767e-10, -6.766167715594326e-10, 
    -6.7872377373159967e-10, -6.808528520400479e-10, -6.8309751775104043e-10, 
    -6.8552526987304642e-10, -6.8816861235729996e-10, 
    -6.9101910818682715e-10, -6.940247516004484e-10, -6.9709097458729221e-10, 
    -7.000850141707888e-10, -7.0284339354799595e-10, -7.0518175617023402e-10, 
    -7.0690646610274308e-10, -7.0782691824756799e-10, 
    -7.0776791658795387e-10, -7.0658111023207259e-10, 
    -7.0415488062408928e-10, -7.0042202109427687e-10, 
    -6.9536487871483325e-10, -6.8901755435960683e-10, 
    -6.8146529603985542e-10, -6.7284096476833233e-10, 
    -6.6331903253872417e-10, -6.5310730616487567e-10, 
    -6.4243704420696796e-10, -6.3155186637489721e-10, 
    -6.2069626402059835e-10, -6.1010414276677235e-10, 
    -5.9998818418492951e-10, -5.9053043486990134e-10, 
    -5.8187476065577874e-10, -5.7412133828099104e-10, 
    -5.6732364987816683e-10, -5.6148787510749381e-10, 
    -5.5657486603288682e-10, -5.5250432743346935e-10, 
    -5.4916114979407096e-10, -5.4640329950620607e-10, 
    -5.4407095616854521e-10, -5.419962148385851e-10, -5.4001291938201167e-10, 
    -5.3796586744146632e-10, -5.3571898903843504e-10, 
    -5.3316182677707896e-10, -5.3021406187519908e-10, 
    -5.2682767410382065e-10, -5.2298675723933373e-10, 
    -5.1870496257104945e-10, -5.1402096253589607e-10, 
    -5.0899227837444156e-10, -5.0368815977203845e-10, -4.98182101429588e-10, 
    -4.9254481988391192e-10, -4.8683818014791903e-10, 
    -4.8111076709690968e-10, -4.753953044301649e-10, -4.6970818696993839e-10, 
    -4.6405096380604701e-10, -4.5841357891346523e-10, 
    -4.5277881860907639e-10, -4.4712752426345602e-10, 
    -4.4144383466540353e-10, -4.3571999069245282e-10, 
    -4.2996007573193046e-10, -4.2418241522522219e-10, 
    -4.1842031065796202e-10, -4.1272119172187666e-10, 
    -4.0714418822867441e-10, -4.0175651227249146e-10, 
    -3.9662894556518176e-10, -3.9183097195603602e-10, -3.8742589726638e-10, 
    -3.834664714546527e-10, -3.7999126290460106e-10, -3.7702208124576711e-10, 
    -3.745625023582008e-10, -3.725975231218274e-10, -3.7109422891203119e-10, 
    -3.7000337156217338e-10, -3.6926154219425514e-10, 
    -3.6879390849606593e-10, -3.6851716122891241e-10, 
    -3.6834265026529058e-10, -3.6817952797975264e-10, 
    -3.6793786646916006e-10, -3.6753164501750175e-10, 
    -3.6688163992443549e-10, -3.6591809000915046e-10, 
    -3.6458311460897008e-10, -3.6283282424772033e-10, 
    -3.6063900076639819e-10, -3.5799028757496811e-10, 
    -3.5489275897672065e-10, -3.5136982109340205e-10, 
    -3.4746143053781166e-10, -3.4322255126624381e-10, 
    -3.3872093428397723e-10, -3.3403426896181216e-10, 
    -3.2924684278726568e-10, -3.2444582349015748e-10, 
    -3.1971736859805266e-10, -3.1514272192723707e-10, 
    -3.1079457240952657e-10, -3.0673378681090437e-10, 
    -3.0300682451522686e-10, -2.9964390863611235e-10, 
    -2.9665820172712012e-10, -2.94045986184601e-10, -2.9178793945197103e-10, 
    -2.8985142389011979e-10, -2.8819369803450203e-10, 
    -2.8676581111702892e-10, -2.8551688965416226e-10, -2.843984960945611e-10, 
    -2.8336869167979613e-10, -2.8239539805520973e-10, 
    -2.8145881134809269e-10, -2.8055251356033579e-10, 
    -2.7968328531268054e-10, -2.7886949512283292e-10, 
    -2.7813831138692024e-10, -2.7752193828194188e-10, 
    -2.7705330889898611e-10, -2.7676162499188757e-10, 
    -2.7666829491924964e-10, -2.7678357017870625e-10, 
    -2.7710432856270426e-10, -2.7761314963964539e-10, -2.782788123729181e-10, 
    -2.7905806202914534e-10, -2.7989851752500003e-10, 
    -2.8074231515969211e-10, -2.8153017642474779e-10, 
    -2.8220542968670065e-10, -2.8271770578374334e-10, 
    -2.8302589484799488e-10, -2.8310027450869056e-10, 
    -2.8292360923066733e-10, -2.8249132313971881e-10, -2.818107664266102e-10, 
    -2.808998061768192e-10, -2.7978488230151473e-10, -2.7849880830832739e-10, 
    -2.7707843269259012e-10, -2.7556240010564851e-10, 
    -2.7398904428356593e-10, -2.7239458569411846e-10, 
    -2.7081158116229839e-10, -2.6926774463891765e-10, -2.677850408492091e-10, 
    -2.6637914619043143e-10, -2.6505918134700064e-10, 
    -2.6382781229499387e-10, -2.6268160517291004e-10, 
    -2.6161168806376459e-10, -2.606046366839843e-10, -2.5964358292904372e-10, 
    -2.5870941497741534e-10, -2.5778204810420786e-10, 
    -2.5684163538201507e-10, -2.558697083363615e-10, -2.5485009856143421e-10, 
    -2.5376969334281662e-10, -2.5261890592712785e-10, 
    -2.5139196430645291e-10, -2.5008692199358225e-10, 
    -2.4870554201578476e-10, -2.4725294767825494e-10, 
    -2.4573722204704929e-10, -2.4416883056186233e-10, 
    -2.4256001537332848e-10, -2.409240991342144e-10, -2.392747485172039e-10, 
    -2.3762521398006182e-10, -2.3598760003847169e-10, 
    -2.3437213572782178e-10, -2.3278660664999542e-10, 
    -2.3123585711358702e-10, -2.2972152413942761e-10, 
    -2.2824194817526822e-10, -2.2679235536260775e-10, 
    -2.2536525367768691e-10, -2.2395105857463316e-10, 
    -2.2253888994456807e-10, -2.2111751848114458e-10, 
    -2.1967632292460134e-10, -2.1820628523176415e-10, 
    -2.1670083341127779e-10, -2.1515657103015996e-10, 
    -2.1357376464995424e-10, -2.1195658991269845e-10, 
    -2.1031309625434661e-10, -2.0865498754114361e-10, 
    -2.0699711485190216e-10, -2.0535682795934876e-10, 
    -2.0375319020969924e-10, -2.0220614097406733e-10, 
    -2.0073558880241768e-10, -1.9936054848735846e-10, 
    -1.9809825047488667e-10, -1.9696330931751594e-10, 
    -1.9596688593128794e-10, -1.951159312964886e-10, -1.9441245038529019e-10, 
    -1.9385289178615569e-10, -1.934276738949511e-10, -1.9312094987647523e-10, 
    -1.9291062469034217e-10, -1.9276879991679765e-10, 
    -1.9266255221242203e-10, -1.9255514575616836e-10, 
    -1.9240759009123531e-10, -1.9218054071160149e-10, 
    -1.9183628568107229e-10, -1.9134081846035628e-10, 
    -1.9066573092599003e-10, -1.8978979599278007e-10, 
    -1.8870013796586913e-10, -1.8739289986159129e-10, 
    -1.8587329630361899e-10, -1.8415520027973703e-10, 
    -1.8226018344762753e-10, -1.8021620671589806e-10, 
    -1.7805603473503846e-10, -1.7581553239007524e-10, 
    -1.7353191798930882e-10, -1.7124213133128988e-10, 
    -1.6898134311192896e-10, -1.6678169186965449e-10, 
    -1.6467124151785133e-10, -1.6267321780576548e-10, 
    -1.6080544817960215e-10, -1.5908011691897998e-10, 
    -1.5750371368938774e-10, -1.5607724412537766e-10, 
    -1.5479668491998342e-10, -1.5365368249430775e-10, 
    -1.5263643301278354e-10, -1.5173074588728091e-10, 
    -1.5092119203313173e-10, -1.5019229407508824e-10, 
    -1.4952960983905107e-10, -1.4892067067348497e-10, 
    -1.4835563789368498e-10, -1.478276569123977e-10, -1.4733281001989889e-10, 
    -1.4686975886715826e-10, -1.4643904594587224e-10, -1.460421960252373e-10, 
    -1.45680682350598e-10, -1.4535496191733147e-10, -1.4506362585342099e-10, 
    -1.4480281462049986e-10, -1.4456599229458221e-10, 
    -1.4434408606636864e-10, -1.4412596765846601e-10, 
    -1.4389929453151445e-10, -1.4365150129946911e-10, 
    -1.4337092412356107e-10, -1.4304784945948408e-10, 
    -1.4267544387512638e-10, -1.4225038282654984e-10, 
    -1.4177319539748095e-10, -1.4124821955889398e-10, 
    -1.4068327756212705e-10, -1.4008902438537955e-10, 
    -1.3947813889416057e-10, -1.3886436436433541e-10, 
    -1.3826155539128512e-10, -1.3768275387841327e-10, 
    -1.3713939292669516e-10, -1.3664064594998755e-10, 
    -1.3619293809400556e-10, -1.3579959342192979e-10, -1.354606841529611e-10, 
    -1.3517294170803421e-10, -1.3492984156862148e-10, 
    -1.3472176275087604e-10, -1.345362832725446e-10, -1.3435858692407837e-10, 
    -1.3417202106579432e-10, -1.3395878449346857e-10, 
    -1.3370076364417424e-10, -1.3338048294470635e-10, 
    -1.3298214063455975e-10, -1.3249264459490302e-10, 
    -1.3190264121258097e-10, -1.3120735933114212e-10, 
    -1.3040728301271636e-10, -1.2950849573071069e-10, 
    -1.2852274961905371e-10, -1.2746711044776357e-10, 
    -1.2636329181302604e-10, -1.2523663804564996e-10, 
    -1.2411487790800372e-10, -1.2302667472534363e-10, 
    -1.2200012924800755e-10, -1.2106127219481355e-10, 
    -1.2023270632285935e-10, -1.1953240381546859e-10, 
    -1.1897279916994901e-10, -1.1856015357260121e-10, 
    -1.1829423924300003e-10, -1.1816835437119535e-10, 
    -1.1816964804703697e-10, -1.1827973602993105e-10, 
    -1.1847557069269408e-10, -1.18730527771303e-10, -1.1901569060333895e-10, 
    -1.1930121721124863e-10, -1.1955779205206408e-10, 
    -1.1975802876454901e-10, -1.1987779854993701e-10, 
    -1.1989734431475428e-10, -1.198021765858363e-10, -1.1958362426717889e-10, 
    -1.1923905339172757e-10, -1.1877173107350923e-10, 
    -1.1819033046859886e-10, -1.1750817149263874e-10, 
    -1.1674224381180843e-10, -1.1591210225783525e-10, 
    -1.1503873917420146e-10, -1.1414348745473619e-10, 
    -1.1324707370036385e-10, -1.123688171458234e-10, -1.1152600379986811e-10, 
    -1.1073344047438713e-10, -1.1000318198262294e-10, 
    -1.0934436923078746e-10, -1.0876315469408891e-10, 
    -1.0826269502030212e-10, -1.0784319726644968e-10, 
    -1.0750200578448789e-10, -1.0723371159104247e-10, 
    -1.0703032355414242e-10, -1.0688153128347478e-10, 
    -1.0677500960271198e-10, -1.0669685044520477e-10, 
    -1.0663204524598439e-10, -1.0656508031467245e-10, 
    -1.0648057186310298e-10, -1.0636392047285747e-10, 
    -1.0620197261734059e-10, -1.0598365218400129e-10, 
    -1.0570046861453532e-10, -1.0534695067305373e-10, 
    -1.0492088074893698e-10, -1.0442338303867176e-10, 
    -1.0385878408137889e-10, -1.0323429776898724e-10, 
    -1.0255949981258897e-10, -1.0184565880794072e-10, 
    -1.0110494179257001e-10, -1.0034957479353484e-10, 
    -9.9590985659372778e-11, -9.8839073150686554e-11, 
    -9.8101565030164583e-11, -9.7383614565317819e-11, -9.668760682046006e-11, 
    -9.6013225121883002e-11, -9.5357743574781341e-11, -9.471653591218157e-11, 
    -9.4083723686868883e-11, -9.3452918185242667e-11, 
    -9.2817965965405547e-11, -9.2173653167686621e-11, 
    -9.1516284239974387e-11, -9.084409163291993e-11, -9.0157474229011755e-11, 
    -8.9459042708208967e-11, -8.8753475576280383e-11, 
    -8.8047242979941905e-11, -8.7348213411421138e-11, 
    -8.6665181076242581e-11, -8.6007348870849625e-11, 
    -8.5383842962410853e-11, -8.4803208608947255e-11, 
    -8.4272955771964979e-11, -8.3799138446832605e-11, 
    -8.3385996599362636e-11, -8.3035649058191581e-11, 
    -8.2747861781243381e-11, -8.251986969918921e-11, -8.2346385295562547e-11, 
    -8.2219660733544955e-11, -8.2129747055946148e-11, 
    -8.2064880205451384e-11, -8.2012061616339477e-11, 
    -8.1957723767490837e-11, -8.188852384161889e-11, -8.1792138427968517e-11, 
    -8.1658047652980391e-11, -8.1478153109969513e-11, 
    -8.1247306362138754e-11, -8.0963513859055115e-11, 
    -8.0627959455327993e-11, -8.0244710503676237e-11, 
    -7.9820264557555986e-11, -7.9362861774909727e-11, 
    -7.8881762653716857e-11, -7.8386457850360582e-11, 
    -7.7886010557899369e-11, -7.7388467529907298e-11, 
    -7.6900513235364297e-11, -7.6427255811382251e-11, 
    -7.5972258145430031e-11, -7.5537646545223696e-11, 
    -7.5124375833477725e-11, -7.4732471231850281e-11, 
    -7.4361285422226887e-11, -7.4009638135563912e-11, 
    -7.3675926138981256e-11, -7.335806680733805e-11, -7.3053448884114416e-11, 
    -7.2758789707774398e-11, -7.2470028589298163e-11, 
    -7.2182281645477849e-11, -7.1889902976949435e-11, 
    -7.1586647942571615e-11, -7.1265981216050054e-11, 
    -7.0921451955875547e-11, -7.0547191589556676e-11, 
    -7.0138358031295782e-11, -6.9691619595566052e-11, 
    -6.9205501166628148e-11, -6.8680627641319729e-11, 
    -6.8119814866512032e-11, -6.7528020442481417e-11, 
    -6.6912107880224874e-11, -6.628053587093969e-11, -6.5642913951785459e-11, 
    -6.5009514462368624e-11, -6.4390741319606218e-11, 
    -6.3796653867384255e-11, -6.3236473617325349e-11, 
    -6.2718175397234843e-11, -6.2248132522036514e-11, 
    -6.1830869819806697e-11, -6.1468876205444257e-11, 
    -6.1162546101403562e-11, -6.0910203793538977e-11, 
    -6.0708260579531015e-11, -6.055146997360209e-11, -6.0433304876238148e-11, 
    -6.0346409894121152e-11, -6.0283145691268554e-11, 
    -6.0236158496583853e-11, -6.0198969280205405e-11, 
    -6.0166486218831288e-11, -6.013545328525625e-11, -6.0104728615284721e-11, 
    -6.0075384702894101e-11, -6.0050618661941123e-11, 
    -6.0035426517654955e-11, -6.0036103063027944e-11, 
    -6.0059564724805384e-11, -6.0112576343924548e-11, 
    -6.0200943831777428e-11, -6.0328735030085528e-11, 
    -6.0497639970532536e-11, -6.0706492724311508e-11, 
    -6.0951037985802076e-11, -6.122393681780242e-11, -6.1515045013927654e-11, 
    -6.1811902743180334e-11, -6.2100423912350065e-11, 
    -6.2365681332907751e-11, -6.2592785180102318e-11, 
    -6.2767710428942109e-11, -6.2878071300517765e-11, 
    -6.2913761330100394e-11, -6.2867461665477297e-11, 
    -6.2734946813204684e-11, -6.2515248234994908e-11, 
    -6.2210623455906102e-11, -6.1826407881685025e-11, 
    -6.1370697789435055e-11, -6.0853998323187061e-11, 
    -6.0288719966011462e-11, -5.9688714794347976e-11, 
    -5.9068710094996046e-11, -5.8443804948307842e-11, 
    -5.7828940273383229e-11, -5.7238436891288179e-11, 
    -5.6685535685268946e-11, -5.6182034759021187e-11, 
    -5.5737933615825357e-11, -5.5361181549184977e-11, 
    -5.5057433638633574e-11, -5.4829922525160724e-11, 
    -5.4679357863250679e-11, -5.4603931259353852e-11, 
    -5.4599364504526819e-11, -5.46591266506973e-11, -5.4774659347169037e-11, 
    -5.4935755916625867e-11, -5.5130980069125349e-11, 
    -5.5348189296942404e-11, -5.5575030721711805e-11, -5.579949184197322e-11, 
    -5.6010355568489253e-11, -5.6197620729770369e-11, 
    -5.6352774149444947e-11, -5.6468993846843807e-11, 
    -5.6541168746920972e-11, -5.6565855955951285e-11, 
    -5.6541099711988811e-11, -5.6466246286571758e-11, 
    -5.6341661425311635e-11, -5.616854143782822e-11, -5.5948664695708263e-11, 
    -5.568428692097947e-11, -5.5378005113859362e-11, -5.5032741928859678e-11, 
    -5.4651709252821102e-11, -5.4238446613603392e-11, 
    -5.3796799075275967e-11, -5.333094660283199e-11, -5.2845368806742187e-11, 
    -5.2344798720124779e-11, -5.1834156329356842e-11, 
    -5.1318496864190536e-11, -5.0802904025076081e-11, 
    -5.0292457608558442e-11, -4.9792135013669284e-11, 
    -4.9306775583391534e-11, -4.8841003204155943e-11, 
    -4.8399141473607511e-11, -4.7985095789633165e-11, 
    -4.7602228536417279e-11, -4.7253163366403028e-11, 
    -4.6939611955280203e-11, -4.6662175886393108e-11, 
    -4.6420192230914868e-11, -4.6211660923166305e-11, 
    -4.6033227023086705e-11, -4.588033067485002e-11, -4.5747442662055433e-11, 
    -4.562844451364285e-11, -4.5517099950228757e-11, -4.5407575991264396e-11, 
    -4.5294969713527339e-11, -4.5175784798136112e-11, 
    -4.5048268219701113e-11, -4.4912616102865448e-11, 
    -4.4770957322928792e-11, -4.4627144795134037e-11, 
    -4.4486346508227397e-11, -4.4354484760634945e-11, -4.423755747609827e-11, 
    -4.4140931604474282e-11, -4.4068680171600799e-11, 
    -4.4023005345399007e-11, -4.4003835907489091e-11, 
    -4.4008629559465367e-11, -4.4032386589392607e-11, -4.406788307457235e-11, 
    -4.4106108459263781e-11, -4.4136850187660514e-11, 
    -4.4149360501965219e-11, -4.4133078327725534e-11, 
    -4.4078329565002082e-11, -4.3976963685305829e-11, 
    -4.3822871244016187e-11, -4.3612366539522048e-11, 
    -4.3344450998848261e-11, -4.3020901653071191e-11, -4.264623202393414e-11, 
    -4.2227531931936254e-11, -4.177419590463553e-11, -4.129757641903652e-11, 
    -4.0810562502453958e-11, -4.0327083855493752e-11, 
    -3.9861599616351316e-11, -3.9428527742052059e-11, 
    -3.9041640375136106e-11, -3.8713468607095071e-11, 
    -3.8454690500159552e-11, -3.8273536533696123e-11, 
    -3.8175286809047227e-11, -3.8161829049395759e-11, 
    -3.8231348404660028e-11, -3.8378207835290233e-11, 
    -3.8593006831668354e-11, -3.8862867666558387e-11, 
    -3.9171953741950806e-11, -3.9502211836440133e-11, 
    -3.9834251247105485e-11, -4.0148383844498952e-11, 
    -4.0425718277378533e-11, -4.0649218219983234e-11, 
    -4.0804664719110727e-11, -4.0881448810028222e-11, 
    -4.0873111242228051e-11, -4.0777620171084199e-11, 
    -4.0597340995254165e-11, -4.0338737628745019e-11, 
    -4.0011790319657704e-11, -3.9629250452025024e-11, 
    -3.9205727832199229e-11, -3.875675740296044e-11, -3.8297828100987482e-11, 
    -3.784353621262164e-11, -3.7406836245701082e-11, -3.6998492065684096e-11, 
    -3.6626675158385869e-11, -3.6296791763722918e-11, 
    -3.6011483918222085e-11, -3.5770797527093184e-11, 
    -3.5572468675041143e-11, -3.5412352271043038e-11, 
    -3.5284870598498842e-11, -3.5183526398822491e-11, 
    -3.5101383354621237e-11, -3.5031542371187696e-11, 
    -3.4967503486327687e-11, -3.4903497175044743e-11, 
    -3.4834665549549262e-11, -3.4757180045405093e-11, 
    -3.4668237993046047e-11, -3.456597483118308e-11, -3.4449331417970327e-11, 
    -3.4317874545806401e-11, -3.4171611840889454e-11, 
    -3.4010844599076715e-11, -3.3836075284168631e-11, 
    -3.3648000290540014e-11, -3.3447554979337606e-11, 
    -3.3236070142998854e-11, -3.3015465249497084e-11, 
    -3.2788485733585826e-11, -3.2558891548568994e-11, -3.23316245349753e-11, 
    -3.2112839432816314e-11, -3.1909814048675319e-11, 
    -3.1730694350619919e-11, -3.1584076725919983e-11, 
    -3.1478431337873259e-11, -3.1421440822083659e-11, 
    -3.1419276200405081e-11, -3.1475892834252597e-11, 
    -3.1592427119887477e-11, -3.1766760421789755e-11, 
    -3.1993308693080012e-11, -3.2263087178902331e-11, 
    -3.2564057080983164e-11, -3.288177179068653e-11, -3.3200226785306759e-11, 
    -3.3502910587155172e-11, -3.377392192086279e-11, -3.399907970957556e-11, 
    -3.4166925486001689e-11, -3.4269503577998288e-11, 
    -3.4302874640464931e-11, -3.4267267723617206e-11, 
    -3.4166920705414788e-11, -3.4009559063772282e-11, 
    -3.3805602774538016e-11, -3.3567166555934802e-11, 
    -3.3306947468232812e-11, -3.3037136343715527e-11, 
    -3.2768405537763865e-11, -3.2509127902789134e-11, 
    -3.2264844168095952e-11, -3.203805750796962e-11, -3.1828321493838143e-11, 
    -3.1632619520529358e-11, -3.1445977851161389e-11, 
    -3.1262208623030226e-11, -3.1074721494424503e-11, 
    -3.0877296094772672e-11, -3.0664752166765858e-11, 
    -3.0433430822808925e-11, -3.0181495693034513e-11, 
    -2.9909010597815624e-11, -2.9617812634891791e-11, 
    -2.9311218997424062e-11, -2.8993682093171764e-11, 
    -2.8670301343740357e-11, -2.8346445471891324e-11, 
    -2.8027318241650071e-11, -2.7717705602820346e-11, -2.742172808864986e-11, 
    -2.7142782313230369e-11, -2.6883474965811434e-11, 
    -2.6645719728322103e-11, -2.6430758448627232e-11, 
    -2.6239342597825487e-11, -2.6071758739906506e-11, 
    -2.5927980224917813e-11, -2.5807684723751933e-11, 
    -2.5710365020613701e-11, -2.5635322555580426e-11, 
    -2.5581779459141317e-11, -2.5548865117257501e-11, 
    -2.5535744721817941e-11, -2.5541613430290944e-11, 
    -2.5565798517859582e-11, -2.5607732615807256e-11, 
    -2.5666983417579938e-11, -2.5743134632132949e-11, 
    -2.5835726238501389e-11, -2.5944044362130568e-11, 
    -2.6066959162257409e-11, -2.6202699564852609e-11, -2.634870183348933e-11, 
    -2.6501463177637618e-11, -2.6656534903208532e-11, -2.680856862407166e-11, 
    -2.6951541044621747e-11, -2.7079025425498664e-11, -2.718461369769376e-11, 
    -2.7262351110189455e-11, -2.7307217393462727e-11, 
    -2.7315526683834385e-11, -2.7285301669856103e-11, 
    -2.7216457961801625e-11, -2.7110882988456455e-11, 
    -2.6972311321187687e-11, -2.6806075268811719e-11, 
    -2.6618691020916123e-11, -2.6417369901951427e-11, 
    -2.6209466013259212e-11, -2.6001935329553024e-11, 
    -2.5800829765766108e-11, -2.5610913699990807e-11, 
    -2.5435376829325309e-11, -2.5275708749779581e-11, 
    -2.5131706633046551e-11, -2.5001644779325022e-11, 
    -2.4882549647812588e-11, -2.4770553961435792e-11, 
    -2.4661328902165992e-11, -2.4550514531291275e-11, -2.443412005884487e-11, 
    -2.4308889932234899e-11, -2.4172551309724379e-11, 
    -2.4023973176186557e-11, -2.3863198871617321e-11, 
    -2.3691368149640087e-11, -2.3510516261940702e-11, 
    -2.3323344021581211e-11, -2.3132901773217501e-11, 
    -2.2942282338652741e-11, -2.2754352912685811e-11, 
    -2.2571552562750468e-11, -2.2395766118536055e-11, 
    -2.2228297134815431e-11, -2.2069925993458608e-11, 
    -2.1921040957973968e-11, -2.1781794836471847e-11, 
    -2.1652257538004285e-11, -2.1532534976432253e-11, 
    -2.1422818205405387e-11, -2.1323355333479271e-11, 
    -2.1234335275077525e-11, -2.1155703398441959e-11, 
    -2.1086964729912606e-11, -2.1026972711881155e-11, 
    -2.0973804636651057e-11, -2.0924688851198631e-11, 
    -2.0876096814825214e-11, -2.0823927693321468e-11, 
    -2.0763843637889383e-11, -2.0691682083495834e-11, 
    -2.0603921332454787e-11, -2.0498129286894111e-11, 
    -2.0373375329151606e-11, -2.0230497847782939e-11, 
    -2.0072243668074939e-11, -1.990319653887411e-11, -1.9729573120822477e-11, 
    -1.955881156001462e-11, -1.9399067415840515e-11, -1.9258615358314523e-11, 
    -1.9145231767499631e-11, -1.9065651180560182e-11, 
    -1.9025055067234936e-11, -1.9026723463603394e-11, 
    -1.9071862261711471e-11, -1.9159566397376855e-11, 
    -1.9286970265135996e-11, -1.9449528645637397e-11, 
    -1.9641419467931376e-11, -1.9855987616420292e-11, 
    -2.0086260775277486e-11, -2.0325415191632786e-11, 
    -2.0567199873503207e-11, -2.080627668983089e-11, -2.1038478445726489e-11, 
    -2.1260922357147691e-11, -2.147205105068668e-11, -2.1671522164284669e-11, 
    -2.1860058690683314e-11, -2.2039195632679951e-11, 
    -2.2211001462352774e-11, -2.2377744351555858e-11, -2.254162602085182e-11, 
    -2.2704470295965865e-11, -2.2867507728276568e-11, 
    -2.3031183741605594e-11, -2.3195069893298892e-11, 
    -2.3357810802459557e-11, -2.3517184046787972e-11, 
    -2.3670190802652175e-11, -2.3813233614722156e-11, -2.394230542675662e-11, 
    -2.4053243702869078e-11, -2.4141959835547147e-11, 
    -2.4204691213144315e-11, -2.4238207656916813e-11, 
    -2.4240010502992107e-11, -2.4208468701369941e-11, 
    -2.4142936871442157e-11, -2.4043803418265686e-11, -2.391252800470785e-11, 
    -2.3751612687146116e-11, -2.3564569523269213e-11, 
    -2.3355830862649853e-11, -2.3130663529305009e-11, 
    -2.2895025586153485e-11, -2.2655431474087826e-11, 
    -2.2418749651429664e-11, -2.2192008308965332e-11, 
    -2.1982148857019651e-11, -2.1795772541659957e-11, 
    -2.1638869970133215e-11, -2.1516567022533068e-11, 
    -2.1432868918937643e-11, -2.1390469667643592e-11, 
    -2.1390586389242806e-11, -2.1432878031248487e-11, 
    -2.1515432017058691e-11, -2.1634824300352534e-11, 
    -2.1786247195284655e-11, -2.1963704997630726e-11, -2.216024036349612e-11, 
    -2.236821180806982e-11, -2.2579572527970931e-11, -2.2786140542107718e-11, 
    -2.297985669225039e-11, -2.3153039268632001e-11, -2.3298578686445049e-11, 
    -2.3410124605165097e-11, -2.3482233103211702e-11, 
    -2.3510503024549836e-11, -2.3491674757114962e-11, 
    -2.3423717780276136e-11, -2.3305905012767607e-11, 
    -2.3138842451013945e-11, -2.2924482515989995e-11, 
    -2.2666098504848465e-11, -2.2368189593119649e-11, 
    -2.2036349683451233e-11, -2.1677046774559632e-11, 
    -2.1297355034201206e-11, -2.0904619740030751e-11, 
    -2.0506098056870162e-11, -2.0108572879564689e-11, 
    -1.9718004042257283e-11, -1.9339192587718133e-11, 
    -1.8975594113225605e-11, -1.8629152656720237e-11, 
    -1.8300354280157018e-11, -1.7988348386966519e-11, 
    -1.7691198472388675e-11, -1.7406230785156069e-11, 
    -1.7130470431378667e-11, -1.6861065434985783e-11, 
    -1.6595694814157021e-11, -1.6332902348747704e-11, 
    -1.6072356252740773e-11, -1.5814933332520886e-11, 
    -1.5562710400910073e-11, -1.531879070556419e-11, -1.5087032962529031e-11, 
    -1.4871665384647358e-11, -1.4676909700412906e-11, 
    -1.4506545028974462e-11, -1.4363542053821402e-11, 
    -1.4249756778877051e-11, -1.4165747366603423e-11, 
    -1.4110699101573415e-11, -1.408247439107502e-11, -1.4077791479071621e-11, 
    -1.409250365452891e-11, -1.4121952006577409e-11, -1.4161367828299177e-11, 
    -1.4206271894927441e-11, -1.425286061303649e-11, -1.4298313834758817e-11, 
    -1.4341027833095152e-11, -1.4380731064408271e-11, -1.441847569316435e-11, 
    -1.4456512171972533e-11, -1.4498069139072489e-11, 
    -1.4547015647140101e-11, -1.4607506952905574e-11, -1.468356621437717e-11, 
    -1.4778719864266599e-11, -1.4895659311069599e-11, 
    -1.5035999599266974e-11, -1.5200124916936288e-11, 
    -1.5387156295680887e-11, -1.5595012403875399e-11, 
    -1.5820557229200234e-11, -1.6059785314222278e-11, 
    -1.6308079230767987e-11, -1.6560411399703417e-11, 
    -1.6811547350237919e-11, -1.7056176743312256e-11, 
    -1.7289010169523199e-11, -1.7504812104603965e-11, 
    -1.7698408590808689e-11, -1.7864675327703382e-11, 
    -1.7998568675534631e-11, -1.809518734534382e-11, -1.8149884328660294e-11, 
    -1.8158464195190446e-11, -1.8117438735419088e-11, 
    -1.8024307860130588e-11, -1.7877878623730093e-11, 
    -1.7678529424994475e-11, -1.7428437837776432e-11, 
    -1.7131681638516907e-11, -1.6794255642372933e-11, 
    -1.6423913391238371e-11, -1.6029906148892661e-11, 
    -1.5622574340668554e-11, -1.5212884543445642e-11, 
    -1.4811863167433481e-11, -1.443007187350075e-11, -1.4077059609684069e-11, 
    -1.3760927851591593e-11, -1.3487934950263895e-11, 
    -1.3262299874819025e-11, -1.3086060719235999e-11, 
    -1.2959099692761222e-11, -1.2879267460268238e-11, 
    -1.2842649339859496e-11, -1.2843882703210543e-11, -1.287655060518273e-11, 
    -1.2933612923962229e-11, -1.3007872121892963e-11, 
    -1.3092384198687888e-11, -1.318090480907909e-11, -1.3268218776229972e-11, 
    -1.3350448050251653e-11, -1.3425226466634581e-11, 
    -1.3491809604981275e-11, -1.3551023609361456e-11, -1.360515306408592e-11, 
    -1.3657663894387097e-11, -1.3712881496696856e-11, 
    -1.3775554632041362e-11, -1.3850448776639925e-11, 
    -1.3941866762753604e-11, -1.405328263941874e-11, -1.4186998333778982e-11, 
    -1.4343922680463921e-11, -1.4523460087988266e-11, 
    -1.4723526089986774e-11, -1.4940643637693304e-11, 
    -1.5170169982411503e-11, -1.5406532264967864e-11, 
    -1.5643550105311793e-11, -1.5874726209140647e-11, 
    -1.6093529011753246e-11, -1.6293642373284685e-11, 
    -1.6469187951354683e-11, -1.6614885810927076e-11, 
    -1.6726185706030187e-11, -1.6799386143527349e-11, 
    -1.6831694850737395e-11, -1.6821326781084124e-11, 
    -1.6767532924943232e-11, -1.6670651414885258e-11, 
    -1.6532130444472886e-11, -1.6354524391140858e-11, 
    -1.6141434830108392e-11, -1.5897440311714377e-11, 
    -1.5627954195633912e-11, -1.5339048171108677e-11, 
    -1.5037234142885803e-11, -1.4729198891109473e-11, 
    -1.4421536012782601e-11, -1.4120479818468627e-11, 
    -1.3831618684055205e-11, -1.3559673537162871e-11, 
    -1.3308327479772955e-11, -1.3080084452758977e-11, 
    -1.2876241592262771e-11, -1.2696906990295461e-11, 
    -1.2541105529782124e-11, -1.2406932614661338e-11, 
    -1.2291789195233138e-11, -1.2192618310796115e-11, 
    -1.2106167609363126e-11, -1.2029255863432637e-11, 
    -1.1958986014396579e-11, -1.1892938046555762e-11, -1.182929501604511e-11, 
    -1.1766905775317201e-11, -1.1705291431881879e-11, 
    -1.1644574768607416e-11, -1.1585361073970135e-11, 
    -1.1528563772578547e-11, -1.147520750343289e-11, -1.1426201334492557e-11, 
    -1.138212532237904e-11, -1.1343026002737188e-11, -1.1308267556789099e-11, 
    -1.1276430915314007e-11, -1.1245296708122158e-11, 
    -1.1211921148504836e-11, -1.1172774856093107e-11, 
    -1.1123959343996039e-11, -1.1061536371244722e-11, 
    -1.0981830044992234e-11, -1.0881767945101803e-11, 
    -1.0759200601546619e-11, -1.061315088292694e-11, -1.0444007235737884e-11, 
    -1.0253599111420411e-11, -1.0045194498969031e-11, 
    -9.8233791362855381e-12, -9.5938687978443139e-12, -9.363254525197686e-12, 
    -9.1386943360914001e-12, -8.927605675174351e-12, -8.7373432518511428e-12, 
    -8.574899365785028e-12, -8.4466232162442242e-12, -8.3580007064710922e-12, 
    -8.3134506080479874e-12, -8.3161661530928464e-12, 
    -8.3680363714267759e-12, -8.469560127725799e-12, -8.6198475585107233e-12, 
    -8.8167010934196607e-12, -9.0567045468984602e-12, 
    -9.3353834558370704e-12, -9.6474246134863688e-12, -9.986899561509523e-12, 
    -1.0347509807329158e-11, -1.0722833401789828e-11, 
    -1.1106532651121199e-11, -1.1492541697028901e-11, 
    -1.1875197077650578e-11, -1.2249310743395112e-11, 
    -1.2610227022725817e-11, -1.2953809293296287e-11, 
    -1.3276446522242575e-11, -1.357502778147029e-11, -1.3846940018208619e-11, 
    -1.4090058034543353e-11, -1.4302772268684925e-11, 
    -1.4483977693206067e-11, -1.4633087292958118e-11, 
    -1.4750008622589917e-11, -1.4835097003199251e-11, 
    -1.4889043740089738e-11, -1.491278064733846e-11, -1.4907287435688308e-11, 
    -1.4873449982915903e-11, -1.4811893165714452e-11, 
    -1.4722874942468326e-11, -1.4606191379000751e-11, 
    -1.4461200447863802e-11, -1.4286861929709172e-11, 
    -1.4081897667580488e-11, -1.3844963953872703e-11, -1.357490680099658e-11, 
    -1.3270989301764338e-11, -1.2933142677823983e-11, -1.256216824608797e-11, 
    -1.2159928319246351e-11, -1.1729412942827922e-11, 
    -1.1274810712197478e-11, -1.0801471974689799e-11, 
    -1.0315838582939983e-11, -9.8252904138547795e-12, 
    -9.3379859578727326e-12, -8.8626353695034955e-12, 
    -8.4082757877118085e-12, -7.984008997834443e-12, -7.5987623149042012e-12, 
    -7.2609889744466484e-12, -6.9784376292284828e-12, 
    -6.7578807639314533e-12, -6.6049158996916371e-12, 
    -6.5237365203359129e-12, -6.5169986395870278e-12, 
    -6.5857116223077561e-12, -6.7291957629157637e-12, 
    -6.9451133381019536e-12, -7.2295725099308979e-12, 
    -7.5772765407629834e-12, -7.9817438853919755e-12, -8.435566892880284e-12, 
    -8.9306761433078579e-12, -9.4585993835923246e-12, 
    -1.0010700789560302e-11, -1.0578356974436581e-11, 
    -1.1153101317331158e-11, -1.172666399058418e-11, -1.2291007837131054e-11, 
    -1.2838287452502938e-11, -1.3360820077295472e-11, 
    -1.3851060393644132e-11, -1.4301604591060648e-11, 
    -1.4705264386856649e-11, -1.5055216657343872e-11, 
    -1.5345200808782528e-11, -1.5569820750061114e-11, 
    -1.5724840588952161e-11, -1.5807527320625551e-11, 
    -1.5816953675014385e-11, -1.5754243995309173e-11, 
    -1.5622713825851862e-11, -1.5427902512079942e-11, 
    -1.5177434240585515e-11, -1.4880771708738201e-11, 
    -1.4548778423553039e-11, -1.4193218412231563e-11, 
    -1.3826124935486294e-11, -1.3459162977210102e-11, -1.310299994126433e-11, 
    -1.2766713723727842e-11, -1.2457360141927584e-11, 
    -1.2179653893811148e-11, -1.193585421866003e-11, -1.1725840266881818e-11, 
    -1.1547378865720247e-11, -1.1396540433589086e-11, 
    -1.1268273740416412e-11, -1.115701790449771e-11, -1.1057329717251525e-11, 
    -1.096445936019043e-11, -1.0874830116176932e-11, -1.0786325252877134e-11, 
    -1.0698422850144267e-11, -1.06121084206315e-11, -1.0529609814296666e-11, 
    -1.045397585443636e-11, -1.0388549406003658e-11, -1.0336370913117927e-11, 
    -1.0299626650049696e-11, -1.0279160201836566e-11, 
    -1.0274105783652327e-11, -1.028170294974896e-11, -1.0297357608083625e-11, 
    -1.0314857766184755e-11, -1.0326819984132507e-11, 
    -1.0325268756519058e-11, -1.0302356236017548e-11, -1.025108751128701e-11, 
    -1.0166041983787711e-11, -1.0043957174340221e-11, 
    -9.8841857112686718e-12, -9.6888954057273321e-12, 
    -9.4630601953735396e-12, -9.2141671841431461e-12, 
    -8.9517218094238385e-12, -8.686544646689654e-12, -8.429950402393863e-12, 
    -8.1928706299759631e-12, -7.9850268496965359e-12, 
    -7.8141940888296716e-12, -7.6856694445092357e-12, 
    -7.6019644137672465e-12, -7.5627766408512139e-12, 
    -7.5652019132649014e-12, -7.6042076064562277e-12, 
    -7.6732666235091949e-12, -7.7651140383772413e-12, 
    -7.8725005156092295e-12, -7.9889135737816698e-12, 
    -8.1091315330004831e-12, -8.229567287339063e-12, -8.3483830303313747e-12, 
    -8.4653672389885413e-12, -8.5815748194065834e-12, 
    -8.6988227699696169e-12, -8.8190766281315936e-12, 
    -8.9438466089098703e-12, -9.0736409800159148e-12, 
    -9.2075847574321028e-12, -9.3432226236035513e-12, 
    -9.4765591241609392e-12, -9.6023078206395284e-12, 
    -9.7143253917888774e-12, -9.806181822458725e-12, -9.8717929316801741e-12, 
    -9.9060266309051285e-12, -9.905242373468398e-12, -9.8676610819500816e-12, 
    -9.7935824263199203e-12, -9.6854123732846388e-12, 
    -9.5474685331886004e-12, -9.3856502899915951e-12, 
    -9.2070270224832885e-12, -9.0193127457155411e-12, 
    -8.8303464405873921e-12, -8.6476095079598171e-12, 
    -8.4778109432407703e-12, -8.326561463347838e-12, -8.1981640191006341e-12, 
    -8.0955088832395391e-12, -8.0200797673451302e-12, 
    -7.9720433649569324e-12, -7.950420757140885e-12, -7.9533127889459074e-12, 
    -7.9781476461986573e-12, -8.0219642354801577e-12, 
    -8.0816643806546453e-12, -8.154266205614349e-12, -8.237104886663315e-12, 
    -8.3280028483538226e-12, -8.425368912136834e-12, -8.52827237303091e-12, 
    -8.6364368941860594e-12, -8.7501983301661931e-12, 
    -8.8704365925396491e-12, -8.9984859363873678e-12, 
    -9.1359896458288855e-12, -9.2847762534793497e-12, 
    -9.4467253702098951e-12, -9.6236113238428838e-12, 
    -9.8169473361342333e-12, -1.0027811280440422e-11, 
    -1.0256686656262761e-11, -1.0503273280957621e-11, 
    -1.0766326181348358e-11, -1.1043505923101e-11, -1.1331255857549943e-11, 
    -1.1624744149499785e-11, -1.1917874482514035e-11, 
    -1.2203369281205649e-11, -1.2472959615181867e-11, 
    -1.2717651914188101e-11, -1.29280947191228e-11, -1.3094978361337468e-11, 
    -1.3209534068612564e-11, -1.326398368046872e-11, -1.325203394403135e-11, 
    -1.3169273735817472e-11, -1.3013538158720073e-11, 
    -1.2785133009039737e-11, -1.24869944699903e-11, -1.212466820760344e-11, 
    -1.1706206117308426e-11, -1.1241906638190349e-11, 
    -1.0743971769924878e-11, -1.0226020460340682e-11, 
    -9.7025929173152347e-12, -9.1885604235644034e-12, 
    -8.6985057137438739e-12, -8.2461354590575397e-12, 
    -7.8437063154445277e-12, -7.5015179154333506e-12, 
    -7.2274855036989721e-12, -7.0268071321932805e-12, 
    -6.9017787452483678e-12, -6.8517133074386345e-12, 
    -6.8730250003056943e-12, -6.9594497277050608e-12, 
    -7.1023875218766268e-12, -7.2913672789450682e-12, 
    -7.5146157194086093e-12, -7.759664407843725e-12, -8.0139948852285776e-12, 
    -8.2656695160560624e-12, -8.5038904797536687e-12, 
    -8.7194863848027785e-12, -8.905272654186107e-12, -9.0562875578814364e-12, 
    -9.1698484164819603e-12, -9.2454964745282495e-12, 
    -9.2847928823462016e-12, -9.2910169172282156e-12, 
    -9.2687729489755481e-12, -9.2235557356656182e-12, 
    -9.1613100543573765e-12, -9.087993901770945e-12, -9.0091966505403797e-12, 
    -8.9298304269445368e-12, -8.8538793312271884e-12, 
    -8.7842667918919678e-12, -8.7227957947379406e-12, 
    -8.6701821488650074e-12, -8.6261653613396542e-12, 
    -8.5896867529027412e-12, -8.5591172198114006e-12, 
    -8.5325238322821159e-12, -8.5079360463607889e-12, 
    -8.4836247700728232e-12, -8.4583343960487752e-12, 
    -8.4314759774172043e-12, -8.4032513346647655e-12, 
    -8.3747108338992845e-12, -8.3476998415937067e-12, 
    -8.3247431790914087e-12, -8.3088388361440463e-12, 
    -8.3032107501809653e-12, -8.3109947974986178e-12, 
    -8.3349457895174525e-12, -8.3771464179600218e-12, 
    -8.4387608853115463e-12, -8.5198733095979604e-12, 
    -8.6193886010851698e-12, -8.7350289336824181e-12, 
    -8.8634145624210886e-12, -9.0002198645963327e-12, 
    -9.1403991606911119e-12, -9.2784196571891525e-12, 
    -9.4085598429043045e-12, -9.525173455932162e-12, -9.622989872873365e-12, 
    -9.6973501566977054e-12, -9.7444246803048636e-12, 
    -9.7614437813773729e-12, -9.7468348280697573e-12, 
    -9.7003437892690352e-12, -9.6231219246872819e-12, 
    -9.5177409689377342e-12, -9.3881682842093178e-12, 
    -9.2396938267357032e-12, -9.0787595132786517e-12, 
    -8.9127787141759802e-12, -8.7498605350286004e-12, 
    -8.5984739304207844e-12, -8.4670739873080833e-12, 
    -8.3637127863926625e-12, -8.2955889890730891e-12, 
    -8.2686348158822034e-12, -8.2871051100652006e-12, 
    -8.3532373565483351e-12, -8.4669739795567503e-12, -8.625808980964554e-12, 
    -8.8247534606681878e-12, -9.0564466867887587e-12, 
    -9.3114141331780255e-12, -9.5784666112355144e-12, 
    -9.8452226183146255e-12, -1.0098713225981801e-11, 
    -1.0326061551402722e-11, -1.0515138951301203e-11, 
    -1.0655212767010301e-11, -1.073750426139619e-11, -1.0755658956607865e-11, 
    -1.0706051444506979e-11, -1.0587986619663537e-11, 
    -1.0403728895260444e-11, -1.0158411262314694e-11, 
    -9.8597982083432282e-12, -9.5179652035259007e-12, 
    -9.1448579288671169e-12, -8.7538137873290083e-12, 
    -8.3589692538585135e-12, -7.9747208132839138e-12, 
    -7.6150606215006718e-12, -7.2929909168624073e-12, 
    -7.0199658272546521e-12, -6.8053610845333359e-12, 
    -6.6560360760387552e-12, -6.5760300908950516e-12, 
    -6.5663533208427281e-12, -6.6249704927844596e-12, 
    -6.7468975732958893e-12, -6.9244857366799333e-12, 
    -7.1478018628191986e-12, -7.4051749197604078e-12, 
    -7.6837522091139203e-12, -7.9701598091918809e-12, 
    -8.2511359522582035e-12, -8.5141521034141856e-12, 
    -8.7479416510200847e-12, -8.942977272545331e-12, -9.0918020222076241e-12, 
    -9.1892715157780071e-12, -9.2326507967051186e-12, 
    -9.2216095712435944e-12, -9.1580920242565894e-12, 
    -9.0461171677785733e-12, -8.8914648258021044e-12, 
    -8.7013444772498355e-12, -8.4839966578309022e-12, -8.248297216171536e-12, 
    -8.003358324508707e-12, -7.758148952937275e-12, -7.5211454630907042e-12, 
    -7.300040929988993e-12, -7.101482620243678e-12, -6.9309031767902807e-12, 
    -6.7923678263679807e-12, -6.688496906578232e-12, -6.620466770012618e-12, 
    -6.588028820260299e-12, -6.5896014320951144e-12, -6.6224034779818101e-12, 
    -6.6826384404180062e-12, -6.7657318621526124e-12, 
    -6.8665915247802436e-12, -6.9799161975809376e-12, 
    -7.1005089624180391e-12, -7.2236025790495975e-12, 
    -7.3451642763700795e-12, -7.4621527074681513e-12, 
    -7.5727059276213984e-12, -7.6762484778254612e-12, 
    -7.7734693144210413e-12, -7.8662087503135935e-12, 
    -7.9572070274399179e-12, -8.0497821303293018e-12, 
    -8.1474022891191567e-12, -8.2532550888520908e-12, -8.369791844034503e-12, 
    -8.4983570805690602e-12, -8.6388762284057226e-12, 
    -8.7896943964958004e-12, -8.947558155314976e-12, -9.107766729871781e-12, 
    -9.2644514856464549e-12, -9.4110251103873481e-12, 
    -9.5406935948329661e-12, -9.6470454253239736e-12, 
    -9.7246300361284093e-12, -9.7694879254406512e-12, 
    -9.7795717125968773e-12, -9.7550355453989685e-12, 
    -9.6983424342256131e-12, -9.6141881936280682e-12, 
    -9.5092218229604606e-12, -9.3916146305296863e-12, 
    -9.2704715918632795e-12, -9.1551698026683642e-12, 
    -9.0546375842158984e-12, -8.9766739306873362e-12, 
    -8.9273339889197905e-12, -8.9104523428262026e-12,
  // Sqw-F(2, 0-1999)
    0.08231993264695131, 0.082096344679358169, 0.081431394683803865, 
    0.08034222115697881, 0.078856401429921757, 0.077010552647195085, 
    0.07484852692387535, 0.072419335378246963, 0.069774949674564588, 
    0.06696812955546208, 0.064050411465848722, 0.061070369076795465, 
    0.058072224670461109, 0.055094854862362215, 0.052171198955709375, 
    0.049328046822985777, 0.046586158235754974, 0.043960648601443796, 
    0.041461567590112672, 0.039094596605556017, 0.036861797136928082, 
    0.03476235287475591, 0.032793262045948693, 0.030949950760693821, 
    0.029226791626363189, 0.027617523281877096, 0.026115575164620597, 
    0.024714307554353492, 0.023407179962136048, 0.022187861745333898, 
    0.021050298074148176, 0.019988742708301852, 0.018997767035721081, 
    0.01807225289815452, 0.017207375124698571, 0.016398578489721625, 
    0.015641552954166416, 0.014932210409472945, 0.014266665570585424, 
    0.013641223033146486, 0.013052371750894808, 0.012496787301878122, 
    0.011971341358205566, 0.011473116858045116, 0.010999426619710807, 
    0.010547832642128241, 0.010116163173842516, 0.0097025248247115201, 
    0.0093053075090272427, 0.008923180769790753, 0.0085550809348524468, 
    0.0082001894784893819, 0.0078579037950805512, 0.0075278022448699404, 
    0.0072096057469451819, 0.0069031383487327298, 0.006608289105771238, 
    0.0063249772996330691, 0.0060531225641908826, 0.0057926209488084563, 
    0.0055433273888958537, 0.0053050445385627101, 0.0050775174915158481, 
    0.0048604336022527173, 0.0046534264296479418, 0.0044560827531015569, 
    0.0042679516392922223, 0.0040885546395989913, 0.0039173963461282225, 
    0.0037539747013486595, 0.003597790620697637, 0.0034483566337889645, 
    0.0033052043694872094, 0.0031678908006234617, 0.0030360032275425848, 
    0.0029091630207671816, 0.0027870281677176202, 0.0026692946824451477, 
    0.0025556969456984927, 0.0024460070492831644, 0.0023400332264064527, 
    0.0022376174603532979, 0.0021386323782260565, 0.0020429775543975978, 
    0.0019505753684356001, 0.0018613665821260901, 0.0017753058165050381, 
    0.0016923571187015343, 0.0016124898063026739, 0.001535674761258493, 
    0.001461881315124382, 0.0013910748239245438, 0.001323214977585608, 
    0.0012582548311218962, 0.0011961404890921551, 0.0011368113280066112, 
    0.0010802006091236963, 0.0010262363203445593, 0.00097484209202958422, 
    0.00092593805606603242, 0.00087944155631826621, 0.00083526766561752008, 
    0.00079332951253459968, 0.00075353846320616656, 0.00071580423343389321, 
    0.00068003502016446933, 0.00064613773790780037, 0.00061401842608035592, 
    0.00058358286158594129, 0.00055473737292114982, 0.00052738981430646207, 
    0.00050145062712911314, 0.00047683389634904297, 0.00045345830435991331, 
    0.00043124789446593947, 0.00041013257850071864, 0.00039004835403377521, 
    0.00037093723077528999, 0.00035274689770477529, 0.00033543018743260726, 
    0.00031894440922600723, 0.00030325062585838413, 0.00028831294282785863, 
    0.00027409786403261575, 0.00026057374917130784, 0.00024771038867546464, 
    0.00023547869509979398, 0.00022385049779053245, 0.00021279842121050402, 
    0.00020229582614947358, 0.00019231679582654176, 0.00018283615371372355, 
    0.00017382950485337497, 0.00016527329600037307, 0.00015714489126719352, 
    0.00014942265905004557, 0.00014208606350098177, 0.00013511575076131306, 
    0.00012849361777154595, 0.00012220285072277079, 0.00011622792168154453, 
    0.00011055453563721464, 0.00010516952569073092, 0.00010006070044664424, 
    9.5216653812551683e-05, 9.062655233172873e-05, 8.6279918093370064e-05, 
    8.2166425784581962e-05, 7.8275730595993594e-05, 7.4597339889506328e-05, 
    7.1120536475968924e-05, 6.7834355861621585e-05, 6.4727614698309322e-05, 
    6.1788983550057668e-05, 5.9007094347376529e-05, 5.6370671643628203e-05, 
    5.3868676855256996e-05, 5.1490455717544691e-05, 4.9225880778283407e-05, 
    4.7065482455190731e-05, 4.5000563656206646e-05, 4.3023294018226532e-05, 
    4.1126780434916134e-05, 3.9305110850897625e-05, 3.7553368528732194e-05, 
    3.5867614419497858e-05, 3.4244836118414487e-05, 3.2682863303736308e-05, 
    3.1180251534839435e-05, 2.9736138677588999e-05, 2.8350080749820172e-05, 
    2.702187628152063e-05, 2.5751389985585886e-05, 2.4538387318564378e-05, 
    2.3382391168514657e-05, 2.2282570393575685e-05, 2.1237667366652016e-05, 
    2.0245968335525588e-05, 1.9305316663348045e-05, 1.8413165310023558e-05, 
    1.7566661666951326e-05, 1.6762755416055508e-05, 1.5998318674099778e-05, 
    1.5270267396269655e-05, 1.4575673793781459e-05, 1.391186119988969e-05, 
    1.3276475137948871e-05, 1.2667527007572116e-05, 1.2083409507566528e-05, 
    1.1522885392913698e-05, 1.0985053207684095e-05, 1.0469295113135991e-05, 
    9.9752127773988635e-06, 9.5025575211053165e-06, 9.0511605850295084e-06, 
    8.6208686114686613e-06, 8.2114883412797318e-06, 7.8227432690431646e-06, 
    7.4542437044027776e-06, 7.1054704822183349e-06, 6.7757715376719995e-06, 
    6.4643697774628826e-06, 6.1703801559250832e-06, 5.8928335977723809e-06, 
    5.6307053580264032e-06, 5.3829455224822069e-06, 5.1485095671494136e-06, 
    4.9263871612606256e-06, 4.7156276759098886e-06, 4.5153611329493342e-06, 
    4.3248135970042425e-06, 4.1433162947913929e-06, 3.9703080600092614e-06, 
    3.8053310664116127e-06, 3.648020225747388e-06, 3.4980870750746975e-06, 
    3.3552994192743434e-06, 3.2194583801509841e-06, 3.0903747735404218e-06, 
    2.9678468439221821e-06, 2.8516412975803481e-06, 2.741479287127646e-06, 
    2.6370285336651118e-06, 2.5379021790737806e-06, 2.4436643070880853e-06, 
    2.3538414364649196e-06, 2.2679387441347111e-06, 2.1854593812522227e-06, 
    2.105925035775049e-06, 2.0288958838315278e-06, 1.953988242487842e-06, 
    1.8808885552894828e-06, 1.8093627577399986e-06, 1.7392605298020755e-06, 
    1.6705143925269329e-06, 1.6031340043844518e-06, 1.5371963280553522e-06, 
    1.4728325577266464e-06, 1.4102128176885909e-06, 1.3495296780558614e-06, 
    1.2909814986642253e-06, 1.2347565292404121e-06, 1.1810185790237082e-06, 
    1.1298949369245435e-06, 1.0814670788886e-06, 1.0357645461197705e-06, 
    9.9276221265645644e-07, 9.523809838066961e-07, 9.1449177836485766e-07, 
    8.7892245535101394e-07, 8.4546716184334802e-07, 8.1389742010415193e-07, 
    7.8397415746525698e-07, 7.5545982832150181e-07, 7.2812979357212611e-07, 
    7.0178221148134421e-07, 6.762458455461346e-07, 6.5138539384205745e-07, 
    6.2710416511136013e-07, 6.0334414594749217e-07, 5.800836952290627e-07, 
    5.5733325063661341e-07, 5.3512952644492547e-07, 5.1352872258793419e-07, 
    4.9259925747704409e-07, 4.7241449436868425e-07, 4.5304586582868153e-07, 
    4.3455672656319584e-07, 4.169971901191947e-07, 4.0040013561308035e-07, 
    3.8477850645224922e-07, 3.7012396317477187e-07, 3.5640689239978627e-07, 
    3.4357771236932957e-07, 3.3156935082449903e-07, 3.2030070680227186e-07, 
    3.0968084831871686e-07, 2.9961365052290242e-07, 2.9000255008259928e-07, 
    2.807550878629821e-07, 2.7178693532209817e-07, 2.6302515088455034e-07, 
    2.5441048521406553e-07, 2.4589864248096553e-07, 2.3746049642472009e-07, 
    2.2908134733012987e-07, 2.2075937673509761e-07, 2.1250350628658708e-07, 
    2.0433088988290953e-07, 1.9626426616950821e-07, 1.8832937363564136e-07, 
    1.8055259079194453e-07, 1.7295891538523862e-07, 1.6557034873669228e-07, 
    1.5840470831707669e-07, 1.5147486003238725e-07, 1.4478834060450571e-07, 
    1.3834733085212446e-07, 1.3214893793765193e-07, 1.2618574643173954e-07, 
    1.2044659877524441e-07, 1.1491756439830633e-07, 1.0958305006203715e-07, 
    1.044269946298652e-07, 9.9434079214738176e-08, 9.4590874094027588e-08, 
    8.9886837962084632e-08, 8.531508791588421e-08, 8.0872869960239748e-08, 
    7.65616815024643e-08, 7.2387025694496828e-08, 6.8357811877315657e-08, 
    6.4485450132182247e-08, 6.0782719406084161e-08, 5.7262511360875013e-08, 
    5.3936565269832217e-08, 5.0814309135439652e-08, 4.7901910618563993e-08, 
    4.5201617924320869e-08, 4.2711440058326383e-08, 4.0425179806029234e-08, 
    3.8332797671225589e-08, 3.6421052816828357e-08, 3.4674343392509069e-08, 
    3.3075654359248941e-08, 3.1607518420066389e-08, 3.0252903472804439e-08, 
    2.8995957333249939e-08, 2.7822563499654985e-08, 2.6720687857032798e-08, 
    2.56805209335666e-08, 2.46944412840713e-08, 2.3756839702926677e-08, 
    2.2863851179877688e-08, 2.2013040676738336e-08, 2.1203082556348128e-08, 
    2.0433462500304563e-08, 1.970421865135605e-08, 1.9015726463465285e-08, 
    1.8368522692080386e-08, 1.7763157657921902e-08, 1.720006354008607e-08, 
    1.6679427800176366e-08, 1.6201065892332671e-08, 1.5764293201110919e-08, 
    1.5367802748820144e-08, 1.5009560003709308e-08, 1.4686729514940787e-08, 
    1.4395647898260643e-08, 1.4131855458918727e-08, 1.3890193042335541e-08, 
    1.3664964044610173e-08, 1.3450153067001068e-08, 1.3239685644677293e-08, 
    1.3027707086234682e-08, 1.2808855359730915e-08, 1.257850256305682e-08, 
    1.2332942954160435e-08, 1.2069511274166348e-08, 1.1786623639437271e-08, 
    1.1483741843196491e-08, 1.1161270511386831e-08, 1.0820402729672947e-08, 
    1.0462933806350474e-08, 1.009106301183371e-08, 9.7072013372579868e-09, 
    9.3137985590008461e-09, 8.9131979671813366e-09, 8.5075216652126932e-09, 
    8.0985858357303004e-09, 7.6878429845339927e-09, 7.2763483192027716e-09, 
    6.8647483737225852e-09, 6.4532923334550077e-09, 6.0418676639226487e-09, 
    5.6300626851873301e-09, 5.2172570257722212e-09, 4.8027385213612125e-09, 
    4.3858405773690275e-09, 3.9660898482599655e-09, 3.5433498231623543e-09, 
    3.1179438803373181e-09, 2.6907410954732319e-09, 2.2631910818413741e-09, 
    1.8372989459411944e-09, 1.4155387802178364e-09, 1.0007114737150765e-09, 
    5.9576039770047496e-10, 2.0356394898535778e-10, -1.7327230361136374e-10, 
    -5.3260117375391513e-10, -8.7287658639386362e-10, 
    -1.1932387303866414e-09, -1.493533654383276e-09, -1.7742675882271575e-09, 
    -2.0365035893592198e-09, -2.2817148082142619e-09, 
    -2.5116123327803406e-09, -2.727967648078472e-09, -2.9324484052838693e-09, 
    -3.1264833298124512e-09, -3.3111669963938628e-09, 
    -3.4872100267286933e-09, -3.6549342711644905e-09, 
    -3.8143082019471766e-09, -3.965013657763672e-09, -4.1065332981239305e-09, 
    -4.2382471288686834e-09, -4.359527298571592e-09, -4.4698216845585256e-09, 
    -4.5687193749592098e-09, -4.6559933939661691e-09, 
    -4.7316190877082615e-09, -4.7957689077203326e-09, 
    -4.8487869384237455e-09, -4.8911481283963443e-09, 
    -4.9234087844052806e-09, -4.9461552779774965e-09, 
    -4.9599579849652025e-09, -4.9653360609013783e-09, 
    -4.9627373571799155e-09, -4.9525349159506796e-09, 
    -4.9350393418138213e-09, -4.9105235107374326e-09, 
    -4.8792544890806992e-09, -4.8415261794332782e-09, 
    -4.7976865836607166e-09, -4.7481543224728463e-09, 
    -4.6934213798816868e-09, -4.6340412852054515e-09, 
    -4.5706048848578631e-09, -4.5037077383723764e-09, 
    -4.4339150346596498e-09, -4.3617299710357261e-09, 
    -4.2875712921179952e-09, -4.2117636735970664e-09, 
    -4.1345427602484279e-09, -4.0560738449448648e-09, 
    -3.9764811124076627e-09, -3.8958824159307702e-09, 
    -3.8144238988278534e-09, -3.7323085642005155e-09, 
    -3.6498143621975428e-09, -3.5672985557906827e-09, -3.485187938211159e-09, 
    -3.4039561836215024e-09, -3.3240919265260556e-09, 
    -3.2460622268013803e-09, -3.1702767990855636e-09, -3.097057865256112e-09, 
    -3.0266196841187228e-09, -2.9590598856906782e-09, 
    -2.8943632867629688e-09, -2.8324167190127801e-09, 
    -2.7730323611691409e-09, -2.7159759074885475e-09, 
    -2.6609959584002418e-09, -2.6078511239926522e-09, 
    -2.5563324299778835e-09, -2.506279340707776e-09, -2.4575891178389991e-09, 
    -2.410219767962619e-09, -2.3641876826012228e-09, -2.3195609922340782e-09, 
    -2.2764498424143372e-09, -2.234994224483348e-09, -2.1953500157159836e-09, 
    -2.1576733312298656e-09, -2.1221036722433924e-09, 
    -2.0887462071756742e-09, -2.0576542817704931e-09, -2.028813356769259e-09, 
    -2.0021282870045859e-09, -1.9774156804070111e-09, 
    -1.9544032089182027e-09, -1.9327370087407683e-09, 
    -1.9119977537234383e-09, -1.8917247416041884e-09, 
    -1.8714466518657699e-09, -1.8507163642889134e-09, 
    -1.8291470015705375e-09, -1.8064456767833952e-09, 
    -1.7824418954661206e-09, -1.757107703806136e-09, -1.7305676952887949e-09, 
    -1.7030976792139291e-09, -1.6751120055081411e-09, 
    -1.6471402984879118e-09, -1.6197953645434226e-09, 
    -1.5937344992233999e-09, -1.5696170925782643e-09, 
    -1.5480613634354426e-09, -1.5296033955850381e-09, 
    -1.5146612169917198e-09, -1.5035065098663277e-09, 
    -1.4962458717955253e-09, -1.4928130761992949e-09, 
    -1.4929728239251387e-09, -1.496335840561616e-09, -1.5023841731683674e-09, 
    -1.5105048713998209e-09, -1.5200294404487791e-09, -1.530276105623746e-09, 
    -1.5405915222739155e-09, -1.5503888656604374e-09, 
    -1.5591792962292616e-09, -1.5665946675179201e-09, 
    -1.5723999802479397e-09, -1.5764951546002128e-09, 
    -1.5789065064381113e-09, -1.5797693255527899e-09, 
    -1.5793034631456953e-09, -1.577784518694096e-09, -1.5755131177610763e-09, 
    -1.572785026592474e-09, -1.5698642340740569e-09, -1.5669610458309806e-09, 
    -1.5642163250738977e-09, -1.5616927934219013e-09, 
    -1.5593734288076747e-09, -1.5571668475374868e-09, 
    -1.5549187299717549e-09, -1.552428397725289e-09, -1.5494690156683682e-09, 
    -1.5458099680759832e-09, -1.5412396110165715e-09, -1.535586724418015e-09, 
    -1.5287388970995237e-09, -1.5206564886039936e-09, 
    -1.5113807976750168e-09, -1.5010358532820934e-09, 
    -1.4898234569947838e-09, -1.4780119482350848e-09, 
    -1.4659194777322705e-09, -1.4538933159659859e-09, -1.442286862133699e-09, 
    -1.4314364206575161e-09, -1.4216395790370547e-09, 
    -1.4131370217805879e-09, -1.4060989908159897e-09, 
    -1.4006173388710122e-09, -1.3967033074725542e-09, 
    -1.3942908782940992e-09, -1.3932448380011012e-09, 
    -1.3933726181137383e-09, -1.394438556979065e-09, -1.3961795127214583e-09, 
    -1.3983205234019809e-09, -1.4005897286630783e-09, 
    -1.4027317772597006e-09, -1.4045193445280779e-09, 
    -1.4057623648772631e-09, -1.4063149536548909e-09, 
    -1.4060797800214612e-09, -1.4050099366510764e-09, -1.403108126576253e-09, 
    -1.4004232287230467e-09, -1.3970441557877853e-09, 
    -1.3930913218742212e-09, -1.3887059182555086e-09, 
    -1.3840377042668307e-09, -1.3792319968795468e-09, 
    -1.3744168710818962e-09, -1.3696915194206671e-09, 
    -1.3651169093741874e-09, -1.3607094296822629e-09, -1.356438301995072e-09, 
    -1.3522269442436831e-09, -1.3479583406243576e-09, 
    -1.3434838972637037e-09, -1.3386351986069604e-09, 
    -1.3332376032679924e-09, -1.3271246988021342e-09, 
    -1.3201524340824977e-09, -1.3122118844684506e-09, 
    -1.3032396985032529e-09, -1.2932254905961367e-09, 
    -1.2822156263657219e-09, -1.2703131812477962e-09, 
    -1.2576739716723474e-09, -1.2444990437035615e-09, 
    -1.2310239309779565e-09, -1.2175055538384114e-09, 
    -1.2042074452463427e-09, -1.1913844539708655e-09, -1.179267780262803e-09, 
    -1.1680515053523205e-09, -1.157881412974946e-09, -1.1488469813914938e-09, 
    -1.1409769954329499e-09, -1.1342391414648319e-09, 
    -1.1285435300299507e-09, -1.123749885656253e-09, -1.1196777655738463e-09, 
    -1.1161190930388725e-09, -1.1128519103921696e-09, 
    -1.1096544075841607e-09, -1.1063180850409012e-09, 
    -1.1026592012645502e-09, -1.0985276529509218e-09, 
    -1.0938128696851454e-09, -1.0884464081235938e-09, 
    -1.0824013834291066e-09, -1.0756889677012926e-09, 
    -1.0683525537204439e-09, -1.0604601783056858e-09, 
    -1.0520960027260102e-09, -1.0433515339477088e-09, 
    -1.0343173019718197e-09, -1.0250755582738678e-09, 
    -1.0156944742969405e-09, -1.0062241520943148e-09, 
    -9.9669465516584325e-10, -9.8711607528648552e-10, 
    -9.7748059104296035e-10, -9.6776625238490181e-10, 
    -9.5794220490294246e-10, -9.4797484253404344e-10, 
    -9.3783438798219978e-10, -9.2750129160155382e-10, 
    -9.1697185244341249e-10, -9.0626248771433066e-10, -8.954122495121051e-10, 
    -8.8448323490886379e-10, -8.7355885621347313e-10, 
    -8.6274000316405617e-10, -8.5213950266318487e-10, 
    -8.4187524738349788e-10, -8.3206269967683062e-10, 
    -8.2280732008005571e-10, -8.1419762733097657e-10, 
    -8.0629936933544132e-10, -7.9915132793701983e-10, 
    -7.9276290873111104e-10, -7.8711368556755939e-10, 
    -7.8215479214829421e-10, -7.7781198980603824e-10, 
    -7.7399002815453003e-10, -7.7057803877698875e-10, 
    -7.6745542523704085e-10, -7.6449797771936606e-10, 
    -7.6158376814638649e-10, -7.5859857446393569e-10, 
    -7.5544052256286131e-10, -7.5202383996347398e-10, 
    -7.4828148745071904e-10, -7.4416672235352674e-10, 
    -7.3965347454328907e-10, -7.3473570507114961e-10, 
    -7.2942576261533403e-10, -7.2375197988885364e-10, 
    -7.1775566786357917e-10, -7.1148783810888085e-10, 
    -7.0500578957102547e-10, -6.9836991642795266e-10, 
    -6.9164083032932364e-10, -6.8487706977139074e-10, 
    -6.7813330125606935e-10, -6.7145916113032262e-10, 
    -6.6489852340135683e-10, -6.5848921923831245e-10, 
    -6.5226291856434694e-10, -6.4624522430547739e-10, 
    -6.4045574193992313e-10, -6.3490826073186835e-10, 
    -6.2961096830319059e-10, -6.2456685198599476e-10, 
    -6.1977433330688484e-10, -6.1522828035799792e-10, 
    -6.1092133550605033e-10, -6.0684560500358644e-10, 
    -6.0299447043567795e-10, -5.9936444427738881e-10, 
    -5.9595666719629492e-10, -5.9277792585601401e-10, 
    -5.8984082062575721e-10, -5.8716307188772117e-10, 
    -5.8476580656931906e-10, -5.8267104064234079e-10, 
    -5.8089847511583378e-10, -5.7946206393097399e-10, 
    -5.7836662384870738e-10, -5.7760506156736948e-10, 
    -5.7715643108605477e-10, -5.7698523447624171e-10, 
    -5.7704202512889276e-10, -5.772653844535731e-10, -5.7758501765177973e-10, 
    -5.7792580042689964e-10, -5.7821223428488937e-10, 
    -5.7837301685998905e-10, -5.783451626169871e-10, -5.7807743144208906e-10, 
    -5.7753264386277407e-10, -5.7668887056632004e-10, 
    -5.7553935758907954e-10, -5.7409140334586396e-10, -5.723642969206354e-10, 
    -5.7038666643493923e-10, -5.6819348802165313e-10, -5.658230858350743e-10, 
    -5.6331433476255022e-10, -5.6070431307865054e-10, 
    -5.5802644602380431e-10, -5.5530929423172352e-10, -5.525758672516439e-10, 
    -5.4984350708020501e-10, -5.4712417211544156e-10, 
    -5.4442507073421462e-10, -5.4174948633187152e-10, 
    -5.3909775782463822e-10, -5.364682256947259e-10, -5.3385817103083752e-10, 
    -5.3126457175606595e-10, -5.2868475961865008e-10, 
    -5.2611682071073926e-10, -5.2355984345421381e-10, 
    -5.2101393586682831e-10, -5.1848012529614895e-10, 
    -5.1596007611020467e-10, -5.1345577464734344e-10, -5.109691176328726e-10, 
    -5.0850155340361106e-10, -5.0605371125513492e-10, 
    -5.0362512195181746e-10, -5.01213967143486e-10, -4.9881696069039207e-10, 
    -4.9642924501065466e-10, -4.9404440752778667e-10, 
    -4.9165454474752394e-10, -4.8925041190017243e-10, 
    -4.8682165378366494e-10, -4.8435713712978745e-10, 
    -4.8184535364180152e-10, -4.7927497434431675e-10, 
    -4.7663543436060681e-10, -4.7391762504191378e-10, 
    -4.7111457900212288e-10, -4.6822213502334661e-10, 
    -4.6523948522825286e-10, -4.6216957414396561e-10, 
    -4.5901925403470108e-10, -4.5579919101088608e-10, 
    -4.5252347297991532e-10, -4.4920899511383025e-10, 
    -4.4587460203488985e-10, -4.4254013327502463e-10, 
    -4.3922541695887871e-10, -4.3594935004710016e-10, 
    -4.3272910090576431e-10, -4.295796036516157e-10, -4.2651324475044952e-10, 
    -4.2353983507996774e-10, -4.206667743957255e-10, -4.1789935362660912e-10, 
    -4.1524107391334822e-10, -4.1269393687435798e-10, 
    -4.1025855186131152e-10, -4.0793408172709174e-10, 
    -4.0571794855995361e-10, -4.0360541266715387e-10, 
    -4.0158900052276258e-10, -3.9965797733345476e-10, 
    -3.9779792262693972e-10, -3.9599055889851017e-10, 
    -3.9421389593187992e-10, -3.9244282304748231e-10, 
    -3.9065004420719359e-10, -3.8880741544135327e-10, 
    -3.8688751051052271e-10, -3.8486536436012386e-10, 
    -3.8272012629718959e-10, -3.8043656896345714e-10, 
    -3.7800620596543927e-10, -3.7542798896675826e-10, 
    -3.7270842531128984e-10, -3.6986122801534111e-10, -3.669063806232084e-10, 
    -3.638688807851973e-10, -3.6077714685475841e-10, -3.57661329145439e-10, 
    -3.545516323997937e-10, -3.5147680683698864e-10, -3.4846290374340033e-10, 
    -3.4553238184815134e-10, -3.4270356931103092e-10, 
    -3.3999050985588687e-10, -3.3740308415785397e-10, 
    -3.3494742703497605e-10, -3.3262645240137271e-10, 
    -3.3044048784778592e-10, -3.2838788053973391e-10, 
    -3.2646554021473629e-10, -3.2466936730843671e-10, 
    -3.2299455083568542e-10, -3.2143571604788369e-10, -3.199869867053016e-10, 
    -3.186419180794619e-10, -3.1739341356010778e-10, -3.162335920349532e-10, 
    -3.1515368697568927e-10, -3.1414395377827549e-10, 
    -3.1319365224766066e-10, -3.1229105219272841e-10, 
    -3.1142351377893194e-10, -3.1057761841145927e-10, 
    -3.0973935300778242e-10, -3.0889433470393524e-10, 
    -3.0802812863661296e-10, -3.0712660278114242e-10, 
    -3.0617633351043785e-10, -3.0516510682648614e-10, 
    -3.0408244328723753e-10, -3.029201435716713e-10, -3.0167285990766759e-10, 
    -3.0033857474631511e-10, -2.9891901332310197e-10, 
    -2.9741987865748992e-10, -2.9585090664795835e-10, 
    -2.9422568195882983e-10, -2.9256121579069285e-10, 
    -2.9087727234861828e-10, -2.8919551601828241e-10, 
    -2.8753847537967477e-10, -2.8592843610277736e-10, 
    -2.8438630827904793e-10, -2.8293054755230525e-10, 
    -2.8157620894395976e-10, -2.8033415780385654e-10, 
    -2.7921050785985805e-10, -2.782062809549389e-10, -2.7731729410600747e-10, 
    -2.7653431209036812e-10, -2.7584337766517396e-10, 
    -2.7522638064316296e-10, -2.7466178766830226e-10, 
    -2.7412556175755375e-10, -2.735921893521868e-10, -2.7303583732485235e-10, 
    -2.7243155166202685e-10, -2.717564694487947e-10, -2.7099096774873851e-10, 
    -2.7011969596846278e-10, -2.691324011625775e-10, -2.6802452286758315e-10, 
    -2.6679747618675279e-10, -2.6545863124178724e-10, 
    -2.6402095783512339e-10, -2.6250241444468339e-10, 
    -2.6092506167578946e-10, -2.5931401145184625e-10, 
    -2.5769624797317826e-10, -2.5609942176395886e-10, 
    -2.5455063716930721e-10, -2.5307530920236924e-10, 
    -2.5169611415574538e-10, -2.504320674104899e-10, -2.4929772808234375e-10, 
    -2.4830255945668471e-10, -2.4745046373322011e-10, 
    -2.4673948750065421e-10, -2.461617522109741e-10, -2.4570363699207213e-10, 
    -2.4534622322326094e-10, -2.4506601761933694e-10, 
    -2.4483597450290629e-10, -2.446267687592222e-10, -2.4440824515223791e-10, 
    -2.4415100220856235e-10, -2.4382794522422268e-10, 
    -2.4341574284082657e-10, -2.4289601904518998e-10, 
    -2.4225623218939328e-10, -2.4149011549789951e-10, 
    -2.4059772711539409e-10, -2.3958506293057638e-10, 
    -2.3846332395391353e-10, -2.3724794507144021e-10, 
    -2.3595747449961798e-10, -2.3461242861117838e-10, 
    -2.3323423072375585e-10, -2.3184425759250978e-10, 
    -2.3046311063584125e-10, -2.291100140062845e-10, -2.2780239447390405e-10, 
    -2.2655551383365778e-10, -2.2538220639823411e-10, 
    -2.2429256872519606e-10, -2.2329366869819721e-10, 
    -2.2238921402202282e-10, -2.2157928668485531e-10, 
    -2.2086009593790038e-10, -2.2022389063601199e-10, 
    -2.1965902177865783e-10, -2.1915025168012955e-10, 
    -2.1867926184458816e-10, -2.1822541812098159e-10, 
    -2.1776668646481003e-10, -2.1728071344550039e-10, 
    -2.1674593456023601e-10, -2.161426687874722e-10, -2.1545412220341874e-10, 
    -2.1466722995814855e-10, -2.1377326938994335e-10, 
    -2.1276824405197184e-10, -2.1165297452684908e-10, -2.104329451051952e-10, 
    -2.091178571781824e-10, -2.0772098306015804e-10, -2.0625829963045031e-10, 
    -2.0474749100812082e-10, -2.0320687097882684e-10, 
    -2.0165429828111196e-10, -2.0010615887164569e-10, 
    -1.9857651205775453e-10, -1.9707643416806568e-10, 
    -1.9561365703082628e-10, -1.9419250228883292e-10, 
    -1.9281414369165113e-10, -1.9147714298379665e-10, 
    -1.9017824315702867e-10, -1.8891329278227764e-10, 
    -1.8767823898322428e-10, -1.8647004975438577e-10, 
    -1.8528749678094009e-10, -1.8413167932134231e-10, 
    -1.8300623639207952e-10, -1.8191724728371775e-10, 
    -1.8087282191273806e-10, -1.7988239781674895e-10, 
    -1.7895589684604512e-10, -1.7810276453666442e-10, 
    -1.7733102694796427e-10, -1.7664644484465056e-10, -1.760518966291131e-10, 
    -1.755469189361501e-10, -1.7512755312529586e-10, -1.7478638802291655e-10, 
    -1.7451283817449907e-10, -1.7429355274970916e-10, 
    -1.7411294976745737e-10, -1.7395377488609614e-10, 
    -1.7379774939020208e-10, -1.7362614804671792e-10, 
    -1.7342042314336074e-10, -1.7316278353096011e-10, 
    -1.7283681055473351e-10, -1.7242802110177851e-10, 
    -1.7192447173416184e-10, -1.7131726649958066e-10, 
    -1.7060105540456417e-10, -1.6977434311080953e-10, 
    -1.6883974393171065e-10, -1.67803944433337e-10, -1.6667752976662081e-10, 
    -1.6547453164651892e-10, -1.6421183324045831e-10, 
    -1.6290837843661764e-10, -1.6158430778449503e-10, 
    -1.6026004398224402e-10, -1.5895543250268318e-10, 
    -1.5768894807699419e-10, -1.5647706542382922e-10, -1.553337539648957e-10, 
    -1.5427015496224424e-10, -1.5329436819666277e-10, -1.524113793910123e-10, 
    -1.5162304228940886e-10, -1.5092813476111324e-10, 
    -1.5032244101134231e-10, -1.4979888657760965e-10, 
    -1.4934770071571924e-10, -1.4895668174305271e-10, 
    -1.4861154304154611e-10, -1.4829634742683482e-10, -1.47994088531437e-10, 
    -1.4768737877172695e-10, -1.4735918962770067e-10, 
    -1.4699364356344094e-10, -1.465767647637169e-10, -1.4609715908034298e-10, 
    -1.4554652425768722e-10, -1.4492001177498186e-10, 
    -1.4421634489603381e-10, -1.4343775160258148e-10, 
    -1.4258968511459087e-10, -1.4168040776333419e-10, 
    -1.4072044066011717e-10, -1.3972197163583917e-10, 
    -1.3869822842793706e-10, -1.3766287613114897e-10, -1.366294512641069e-10, 
    -1.3561087536264064e-10, -1.3461900718960311e-10, 
    -1.3366427765236588e-10, -1.3275535908528858e-10, 
    -1.3189892862177123e-10, -1.310994583297782e-10, -1.3035910720025971e-10, 
    -1.2967768216475125e-10, -1.2905271768531743e-10, -1.284796746691595e-10, 
    -1.2795227739317197e-10, -1.2746296573466053e-10, 
    -1.2700350200752809e-10, -1.2656561446935926e-10, 
    -1.2614175211368397e-10, -1.2572576208087387e-10, 
    -1.2531353978074865e-10, -1.2490350340201969e-10, 
    -1.2449687993323646e-10, -1.2409772853619049e-10, 
    -1.2371271294021507e-10, -1.2335057718118418e-10, -1.230214104061697e-10, 
    -1.2273570123981057e-10, -1.2250332794975247e-10, 
    -1.2233250571216086e-10, -1.2222886317211594e-10, -1.221946719657485e-10, 
    -1.2222834888804937e-10, -1.22324247424403e-10, -1.2247277495804604e-10, 
    -1.226607953229007e-10, -1.2287230867638778e-10, -1.2308928634545531e-10, 
    -1.2329267318113827e-10, -1.2346336959741709e-10, -1.235832233880644e-10, 
    -1.2363588591428208e-10, -1.2360757209222177e-10, 
    -1.2348760748097709e-10, -1.2326884002685375e-10, 
    -1.2294784972563648e-10, -1.2252501295986284e-10, 
    -1.2200440150810533e-10, -1.2139357659074613e-10, 
    -1.2070323703092188e-10, -1.1994679832781779e-10, 
    -1.1913987059105542e-10, -1.1829969363254128e-10, 
    -1.1744450880787463e-10, -1.1659293036456758e-10, 
    -1.1576328946528097e-10, -1.1497303026260192e-10, 
    -1.1423812102169889e-10, -1.1357254942022528e-10, 
    -1.1298786405227024e-10, -1.1249283242827014e-10, 
    -1.1209317393365898e-10, -1.1179139485910782e-10, 
    -1.1158672319504121e-10, -1.1147518126659491e-10, 
    -1.1144973211714612e-10, -1.1150056350909704e-10, 
    -1.1161545959936829e-10, -1.1178030237932984e-10, 
    -1.1197961160947032e-10, -1.1219718007002148e-10, -1.124167038986249e-10, 
    -1.1262242362004861e-10, -1.127996799205515e-10, -1.1293542541858137e-10, 
    -1.1301857293655885e-10, -1.1304024914774057e-10, 
    -1.1299386473401222e-10, -1.1287510315501702e-10, 
    -1.1268174733195332e-10, -1.1241346957390643e-10, 
    -1.1207152892181485e-10, -1.1165849291985079e-10, 
    -1.1117794987267147e-10, -1.1063426632333409e-10, 
    -1.1003239521881057e-10, -1.0937774332049281e-10, -1.086760678290761e-10, 
    -1.0793345772389678e-10, -1.0715629012014396e-10, 
    -1.0635122858816898e-10, -1.05525210246387e-10, -1.0468541483624151e-10, 
    -1.038392050995576e-10, -1.0299406060609168e-10, -1.021574473370873e-10, 
    -1.0133669695983897e-10, -1.0053883388880055e-10, 
    -9.9770398967745112e-11, -9.9037252595096653e-11, 
    -9.8344406050834763e-11, -9.7695826440483011e-11, 
    -9.7094296549755812e-11, -9.6541306483511833e-11, 
    -9.6036982929828972e-11, -9.5580118478232673e-11, -9.516823550050569e-11, 
    -9.4797772162180835e-11, -9.4464307446967471e-11, 
    -9.4162878826441651e-11, -9.3888342214815882e-11, 
    -9.3635743160252379e-11, -9.340067892749062e-11, -9.3179618965679968e-11, 
    -9.2970113754239035e-11, -9.2770911998163287e-11, 
    -9.2581918669618643e-11, -9.2404031006057786e-11, 
    -9.2238825184813949e-11, -9.2088159480090269e-11, 
    -9.1953688035966795e-11, -9.1836381488344519e-11, 
    -9.1736071353783841e-11, -9.1651095022831381e-11, 
    -9.1578053193342355e-11, -9.1511738136821629e-11, 
    -9.1445209519932101e-11, -9.1370028675360471e-11, 
    -9.1276648530577101e-11, -9.11548949826589e-11, -9.099451226032459e-11, 
    -9.0785748731461901e-11, -9.0519944036249996e-11, 
    -9.0190084144393925e-11, -8.979128989760113e-11, -8.9321233229024678e-11, 
    -8.8780475854484732e-11, -8.8172687578843594e-11, 
    -8.7504730366669531e-11, -8.6786617251786098e-11, 
    -8.6031311162428326e-11, -8.5254344072887992e-11, 
    -8.4473282929706756e-11, -8.3707015847730626e-11, -8.297490730741288e-11, 
    -8.2295847276009765e-11, -8.1687245220814634e-11, 
    -8.1164038004368702e-11, -8.0737787828633445e-11, 
    -8.0415898558475336e-11, -8.0201092134588582e-11, 
    -8.0091110693229232e-11, -8.0078714713904862e-11, 
    -8.0151982281085378e-11, -8.029490558432188e-11, -8.0488195856163674e-11, 
    -8.0710326927706405e-11, -8.0938665237044158e-11, 
    -8.1150652121124872e-11, -8.1324957380589737e-11, 
    -8.1442533423683784e-11, -8.1487490363376288e-11, 
    -8.1447767793019149e-11, -8.131556260003398e-11, -8.1087506163828829e-11, 
    -8.0764592896874859e-11, -8.0351893331882026e-11, -7.985807068971725e-11, 
    -7.9294759914346947e-11, -7.8675845504939718e-11, 
    -7.8016679934861041e-11, -7.7333296926759118e-11, 
    -7.6641640536425913e-11, -7.5956846569843551e-11, 
    -7.5292618171165814e-11, -7.4660695270911303e-11, -7.407043879935024e-11, 
    -7.3528558265088637e-11, -7.3039001881366629e-11, 
    -7.2602992844223178e-11, -7.2219225765246352e-11, 
    -7.1884223974826448e-11, -7.1592816048934692e-11, -7.133870688442098e-11, 
    -7.1115086807493187e-11, -7.0915246096707192e-11, 
    -7.0733082621497545e-11, -7.0563523863604914e-11, 
    -7.0402735608908541e-11, -7.0248187149898359e-11, 
    -7.0098485952552132e-11, -6.9953089292196273e-11, -6.981188807243779e-11, 
    -6.9674775329951878e-11, -6.9541231528797482e-11, 
    -6.9410038040225255e-11, -6.9279158960972098e-11, 
    -6.9145818828789845e-11, -6.9006774682872882e-11, 
    -6.8858765660778162e-11, -6.8699049360663885e-11, 
    -6.8525991936070811e-11, -6.8339542979674745e-11, 
    -6.8141601466862131e-11, -6.7936125301888023e-11, 
    -6.7728999483393524e-11, -6.7527628047595106e-11, 
    -6.7340308588355805e-11, -6.7175424113263233e-11, 
    -6.7040585216361281e-11, -6.6941785023369087e-11, 
    -6.6882703063652707e-11, -6.686420375483124e-11, -6.6884135709967887e-11, 
    -6.693740429787785e-11, -6.7016354304402834e-11, -6.711137884609355e-11, 
    -6.7211721609108853e-11, -6.7306344038905698e-11, 
    -6.7384820111346958e-11, -6.7438111919956728e-11, 
    -6.7459220164485738e-11, -6.7443597253091848e-11, 
    -6.7389370960953176e-11, -6.7297279679937012e-11, 
    -6.7170440246077309e-11, -6.7013915117467933e-11, 
    -6.6834156537749882e-11, -6.6638354396733408e-11, -6.643379053349647e-11, 
    -6.6227190428457566e-11, -6.6024168980782893e-11, 
    -6.5828772351814722e-11, -6.5643174508426631e-11, 
    -6.5467517969539665e-11, -6.5299929442404537e-11, -6.513668314827856e-11, 
    -6.4972507842769881e-11, -6.480101045002495e-11, -6.4615172238902631e-11, 
    -6.4407888101776402e-11, -6.4172480862638595e-11, 
    -6.3903195541085654e-11, -6.3595572912529905e-11, 
    -6.3246735094889336e-11, -6.2855533684496897e-11, 
    -6.2422557148943264e-11, -6.194999892565087e-11, -6.1441470248830189e-11, 
    -6.0901660628268212e-11, -6.0336026583116257e-11, 
    -5.9750403970397986e-11, -5.9150711487760659e-11, 
    -5.8542629077679534e-11, -5.7931425572986339e-11, 
    -5.7321792316454929e-11, -5.6717831342240938e-11, 
    -5.6123037585987636e-11, -5.5540446746016399e-11, 
    -5.4972721048957692e-11, -5.4422357886901426e-11, 
    -5.3891827963713037e-11, -5.3383761933532136e-11, -5.290104536237268e-11, 
    -5.2446938382189309e-11, -5.2025059655485632e-11, -5.163940285581131e-11, 
    -5.1294190118720813e-11, -5.0993761780007242e-11, 
    -5.0742333038007301e-11, -5.0543761937285797e-11, 
    -5.0401241067500692e-11, -5.0317038870736793e-11, 
    -5.0292172513211663e-11, -5.0326191560726545e-11, 
    -5.0416942255146352e-11, -5.0560469260230908e-11, 
    -5.0750965165492294e-11, -5.0980862599769367e-11, 
    -5.1241007099135782e-11, -5.1520987381910932e-11, 
    -5.1809524084522423e-11, -5.2094968252474486e-11, 
    -5.2365833561924458e-11, -5.2611366324776156e-11, 
    -5.2822037815965508e-11, -5.29900520913684e-11, -5.3109664691764042e-11, 
    -5.3177437359043449e-11, -5.3192291334743092e-11, 
    -5.3155455254721927e-11, -5.3070224383307467e-11, 
    -5.2941637734102012e-11, -5.2776023234002141e-11, 
    -5.2580525153367176e-11, -5.2362573878748221e-11, 
    -5.2129441361082728e-11, -5.1887789072764944e-11, 
    -5.1643363239343972e-11, -5.1400740449919251e-11, 
    -5.1163233548209821e-11, -5.0932853698767968e-11, 
    -5.0710403788982444e-11, -5.0495612331567336e-11, 
    -5.0287336881554369e-11, -5.0083756537691212e-11, 
    -4.9882607838597106e-11, -4.9681363458753297e-11, 
    -4.9477407729189879e-11, -4.9268165412909067e-11, 
    -4.9051227912030575e-11, -4.8824423758909706e-11, 
    -4.8585948049431077e-11, -4.8334432679711831e-11, 
    -4.8069077826930687e-11, -4.7789749407842753e-11, 
    -4.7497131901128293e-11, -4.7192815875686578e-11, 
    -4.6879385780580899e-11, -4.6560407845600045e-11, 
    -4.6240384113603055e-11, -4.5924553345310695e-11, 
    -4.5618624314038073e-11, -4.532837931114017e-11, -4.5059243228844318e-11, 
    -4.4815782128284283e-11, -4.4601245703089957e-11, 
    -4.4417139560711587e-11, -4.4262975382866397e-11, -4.413613287792769e-11, 
    -4.403195151422089e-11, -4.3944001478314192e-11, -4.3864560102420495e-11, 
    -4.3785226080514544e-11, -4.3697643867732087e-11, 
    -4.3594244394115349e-11, -4.346894452857047e-11, -4.3317719194447176e-11, 
    -4.3139033169322272e-11, -4.2934008484662105e-11, -4.270640444158748e-11, 
    -4.2462320812093364e-11, -4.2209761497790882e-11, -4.195797921011088e-11, 
    -4.1716790837128391e-11, -4.1495816935302354e-11, 
    -4.1303802751562572e-11, -4.1148026036319632e-11, 
    -4.1033847357338972e-11, -4.0964435662724358e-11, 
    -4.0940699842867323e-11, -4.09613715651839e-11, -4.1023272891703433e-11, 
    -4.1121680286034865e-11, -4.1250796886441564e-11, 
    -4.1404228838450359e-11, -4.1575493471407772e-11, 
    -4.1758455377251208e-11, -4.1947710511950325e-11, 
    -4.2138865474761631e-11, -4.2328744425919565e-11, 
    -4.2515461581658662e-11, -4.269842625745068e-11, -4.287822440896079e-11, 
    -4.3056470665679571e-11, -4.3235541947631088e-11, 
    -4.3418303954643186e-11, -4.3607757062039996e-11, 
    -4.3806722682363353e-11, -4.4017468714563267e-11, 
    -4.4241406529251318e-11, -4.4478787942502833e-11, 
    -4.4728521688431097e-11, -4.4988030413744826e-11, 
    -4.5253266268409294e-11, -4.5518804673695863e-11, 
    -4.5778093400580461e-11, -4.6023782694502838e-11, 
    -4.6248188191682902e-11, -4.6443769051646651e-11, 
    -4.6603665346843773e-11, -4.6722186891618315e-11, 
    -4.6795248811254096e-11, -4.6820692298639206e-11, 
    -4.6798485762924312e-11, -4.6730750554883737e-11, 
    -4.6621646251154526e-11, -4.6477094825486947e-11, -4.630440001591211e-11, 
    -4.6111748980973881e-11, -4.5907680233156738e-11, 
    -4.5700544833377713e-11, -4.5498002199835477e-11, 
    -4.5306586457464687e-11, -4.5131392385193273e-11, 
    -4.4975880281590752e-11, -4.484181637923246e-11, -4.4729348335332961e-11, 
    -4.463720100635866e-11, -4.4562958300415359e-11, -4.4503414362076142e-11, 
    -4.4454932656413436e-11, -4.4413815547035868e-11, -4.437660206246949e-11, 
    -4.4340318394650747e-11, -4.4302624898925458e-11, 
    -4.4261871881349244e-11, -4.4217047226865545e-11, 
    -4.4167682482583846e-11, -4.4113650691262337e-11, 
    -4.4054969530613304e-11, -4.3991561499946816e-11, 
    -4.3923062249723551e-11, -4.3848649512085181e-11, 
    -4.3766933970128087e-11, -4.3675909943713173e-11, 
    -4.3573002529688452e-11, -4.3455152928824253e-11, -4.331900400838931e-11, 
    -4.3161113778662139e-11, -4.2978214530936403e-11, 
    -4.2767473218631255e-11, -4.2526774635849911e-11, -4.225493350901973e-11, 
    -4.1951870348401309e-11, -4.1618701082316698e-11, 
    -4.1257743796456673e-11, -4.087240620764732e-11, -4.0467007819355479e-11, 
    -4.0046498020604456e-11, -3.9616137668476184e-11, 
    -3.9181143265900466e-11, -3.87463676240107e-11, -3.8315997471597897e-11, 
    -3.7893378450354422e-11, -3.748090248842533e-11, -3.7080018292069332e-11, 
    -3.6691325279540325e-11, -3.6314790424859377e-11, 
    -3.5949964019347355e-11, -3.5596237355157994e-11, 
    -3.5253045281118838e-11, -3.4920057084132684e-11, 
    -3.4597218489080882e-11, -3.4284772948922921e-11, 
    -3.3983156135773808e-11, -3.3692850000011806e-11, 
    -3.3414181975858309e-11, -3.3147184341618193e-11, 
    -3.2891436716833469e-11, -3.264602903549158e-11, -3.2409567699033078e-11, 
    -3.2180333743448697e-11, -3.1956472142861534e-11, 
    -3.1736277185947482e-11, -3.1518475004605441e-11, 
    -3.1302533287731557e-11, -3.1088888406387732e-11, -3.087912360049992e-11, 
    -3.0676018501817668e-11, -3.0483524708401638e-11, -3.030659238322766e-11, 
    -3.0150929948283099e-11, -3.0022662986394239e-11, -2.992795473169639e-11, 
    -2.9872577413637531e-11, -2.986153645228921e-11, -2.9898666807905062e-11, 
    -2.9986354568652964e-11, -3.0125289681293105e-11, 
    -3.0314349736095238e-11, -3.0550584843362736e-11, 
    -3.0829314205998407e-11, -3.1144314658057679e-11, 
    -3.1488135960263273e-11, -3.1852439023336094e-11, 
    -3.2228391475629786e-11, -3.2607037591134459e-11, 
    -3.2979679810743087e-11, -3.3338129036364279e-11, 
    -3.3674922221745605e-11, -3.3983392991740946e-11, -3.425770235758332e-11, 
    -3.4492746758728933e-11, -3.4684060684042721e-11, 
    -3.4827686688005335e-11, -3.492011334799798e-11, -3.4958254884354569e-11, 
    -3.4939537572250309e-11, -3.4862067186957094e-11, 
    -3.4724909615013103e-11, -3.4528384834655327e-11, 
    -3.4274410307043725e-11, -3.3966761546347829e-11, 
    -3.3611268829923462e-11, -3.321583473358485e-11, -3.2790311796093248e-11, 
    -3.2346164093068604e-11, -3.1895988803779801e-11, 
    -3.1452861428187358e-11, -3.102964856007044e-11, -3.063825557741031e-11, 
    -3.0288963692818411e-11, -2.9989851133043319e-11, 
    -2.9746404810724506e-11, -2.9561290733455647e-11, 
    -2.9434374513503579e-11, -2.9362890420394303e-11, 
    -2.9341794483576068e-11, -2.9364202882020979e-11, 
    -2.9421961635099117e-11, -2.9506159637270312e-11, 
    -2.9607674901802983e-11, -2.9717629685302035e-11, 
    -2.9827812327359725e-11, -2.9930970183490585e-11, 
    -3.0021075545038615e-11, -3.0093466968774211e-11, 
    -3.0144984764097919e-11, -3.0173994275638025e-11, 
    -3.0180418374239536e-11, -3.0165659338565366e-11, 
    -3.0132530406131984e-11, -3.0085066450824993e-11, 
    -3.0028329843386965e-11, -2.9968101487601435e-11, 
    -2.9910570939416274e-11, -2.9861932593754753e-11, 
    -2.9828004541686636e-11, -2.9813824562555152e-11, 
    -2.9823289990189282e-11, -2.9858849204792034e-11, 
    -2.9921300499033668e-11, -3.0009657492615643e-11, -3.012115600029161e-11, 
    -3.0251340789285268e-11, -3.039427843173521e-11, -3.0542832417969974e-11, 
    -3.0689003695753083e-11, -3.082429975121841e-11, -3.0940141982495272e-11, 
    -3.1028226287217554e-11, -3.1080887449410916e-11, 
    -3.1091395905125748e-11, -3.1054226127919283e-11, 
    -3.0965261487179591e-11, -3.0821931636947593e-11, -3.062330901075034e-11, 
    -3.0370154622573222e-11, -3.0064906635988502e-11, 
    -2.9711628990756047e-11, -2.9315919198026068e-11, 
    -2.8884775942730482e-11, -2.8426425043045361e-11, 
    -2.7950102638455134e-11, -2.7465802341279663e-11, 
    -2.6983978749287411e-11, -2.6515221399620095e-11, -2.606987052727313e-11, 
    -2.5657646884526605e-11, -2.528724807118216e-11, -2.4965964772589676e-11, 
    -2.4699342896557825e-11, -2.4490899235266622e-11, 
    -2.4341913560519878e-11, -2.4251340682270949e-11, 
    -2.4215839092255373e-11, -2.4229924300413272e-11, -2.428623864005219e-11, 
    -2.4375958304713802e-11, -2.44892402276809e-11, -2.4615762257424753e-11, 
    -2.4745255763867972e-11, -2.4868011865229421e-11, -2.497534237628123e-11, 
    -2.5059921926202205e-11, -2.5116022324377304e-11, 
    -2.5139612174032257e-11, -2.5128326837460359e-11, -2.508132548999973e-11, 
    -2.4999049368460752e-11, -2.4882939752811084e-11, 
    -2.4735114663958611e-11, -2.4558083508056305e-11, 
    -2.4354502002547548e-11, -2.4127020428823639e-11, 
    -2.3878187230944002e-11, -2.3610453268610476e-11, 
    -2.3326268147936677e-11, -2.3028192186368765e-11, 
    -2.2719034343690305e-11, -2.2401993301558963e-11, 
    -2.2080732687405008e-11, -2.1759425213139808e-11, 
    -2.1442710043468509e-11, -2.1135597969304186e-11, -2.084332603489876e-11, 
    -2.0571183433297995e-11, -2.0324320203075655e-11, 
    -2.0107588397486288e-11, -1.9925401448258765e-11, 
    -1.9781648623892123e-11, -1.9679627782761687e-11, 
    -1.9622026444702271e-11, -1.9610926706588538e-11, 
    -1.9647808725015315e-11, -1.9733535442474808e-11, 
    -1.9868358305064449e-11, -2.005184882240449e-11, -2.0282852409106569e-11, 
    -2.0559446813130644e-11, -2.0878871088515432e-11, 
    -2.1237505801642119e-11, -2.1630877484428616e-11, 
    -2.2053696249764558e-11, -2.2499948547379111e-11, 
    -2.2963023683972973e-11, -2.3435862782267824e-11, 
    -2.3911148533237373e-11, -2.4381480871212056e-11, -2.48395581437588e-11, 
    -2.5278351986916928e-11, -2.5691245800665637e-11, 
    -2.6072172044622443e-11, -2.64157277860832e-11, -2.6717257980872821e-11, 
    -2.6972945409613634e-11, -2.7179882059154571e-11, 
    -2.7336100727995153e-11, -2.7440611768193499e-11, 
    -2.7493410874988092e-11, -2.749544491034389e-11, -2.7448538084143031e-11, 
    -2.7355303334738273e-11, -2.7218981371010471e-11, 
    -2.7043266501635339e-11, -2.683213040398453e-11, -2.6589608465641068e-11, 
    -2.6319616873962062e-11, -2.6025789826731071e-11, 
    -2.5711355951500961e-11, -2.5379060512646714e-11, 
    -2.5031153984712068e-11, -2.4669421081130542e-11, 
    -2.4295271358216616e-11, -2.3909847858212452e-11, 
    -2.3514206685925677e-11, -2.310947609169784e-11, -2.2697038308266358e-11, 
    -2.2278693000550532e-11, -2.185682143693521e-11, -2.1434498808141835e-11, 
    -2.1015583684716819e-11, -2.0604746119357043e-11, 
    -2.0207475303932844e-11, -1.9829988204662265e-11, 
    -1.9479126667179861e-11, -1.9162166340497029e-11, 
    -1.8886583434320077e-11, -1.8659779910079124e-11, 
    -1.8488774979857221e-11, -1.8379881494303189e-11, 
    -1.8338388209834239e-11, -1.8368254629881131e-11, 
    -1.8471889368977768e-11, -1.864994865208938e-11, -1.8901264531336917e-11, 
    -1.9222854460325318e-11, -1.9610014377758085e-11, 
    -2.0056521255057889e-11, -2.0554911199246352e-11, 
    -2.1096792319735421e-11, -2.1673201144907597e-11, 
    -2.2274924495817791e-11, -2.2892800905331967e-11, 
    -2.3517951466251428e-11, -2.4141924102672397e-11, 
    -2.4756757209869569e-11, -2.535498459304259e-11, -2.5929554213236569e-11, 
    -2.6473744056895466e-11, -2.6981053815687265e-11, 
    -2.7445150908245277e-11, -2.7859861189677289e-11, 
    -2.8219236978797968e-11, -2.8517711046152884e-11, 
    -2.8750317658899767e-11, -2.8912978652969539e-11, 
    -2.9002812993391963e-11, -2.901843080882241e-11, -2.8960193530386542e-11, 
    -2.883037874735444e-11, -2.8633230268990388e-11, -2.8374889160446013e-11, 
    -2.8063164136703764e-11, -2.7707197367886213e-11, 
    -2.7317003957371701e-11, -2.6902949180466018e-11, 
    -2.6475210515554188e-11, -2.6043240638713379e-11, 
    -2.5615322138739901e-11, -2.5198227352262048e-11, 
    -2.4797012628397565e-11, -2.4414979445159038e-11, -2.405378247707171e-11, 
    -2.3713670147169419e-11, -2.3393841280538615e-11, 
    -2.3092856449467064e-11, -2.2809045388905551e-11, 
    -2.2540896455645058e-11, -2.2287376327342936e-11, 
    -2.2048115329944544e-11, -2.1823485885805672e-11, 
    -2.1614539287699979e-11, -2.1422815560784684e-11, 
    -2.1250066432497368e-11, -2.1097897923172439e-11, 
    -2.0967394190391125e-11, -2.0858766227701695e-11, 
    -2.0771067565628192e-11, -2.0701989112569615e-11, 
    -2.0647806601710598e-11, -2.0603489596335008e-11, 
    -2.0562950387747091e-11, -2.0519436641375831e-11, 
    -2.0466042151311301e-11, -2.039629853942433e-11, -2.0304771691372043e-11, 
    -2.018762265607208e-11, -2.0043056074949965e-11, -1.9871630708703096e-11, 
    -1.967636161753018e-11, -1.9462606084957063e-11, -1.9237748607702989e-11, 
    -1.90106775796144e-11, -1.8791128421030446e-11, -1.8588931976159254e-11, 
    -1.8413239794023149e-11, -1.8271817569926202e-11, 
    -1.8170435643956555e-11, -1.8112453917078324e-11, 
    -1.8098595708076208e-11, -1.8126961774212183e-11, 
    -1.8193241225470834e-11, -1.8291128801666366e-11, 
    -1.8412865838123547e-11, -1.8549873645373404e-11, 
    -1.8693404493534042e-11, -1.8835155035720077e-11, 
    -1.8967787023238469e-11, -1.9085301613192721e-11, 
    -1.9183256222903463e-11, -1.9258826689798134e-11, 
    -1.9310693239809213e-11, -1.9338825530201445e-11, 
    -1.9344154125898154e-11, -1.9328220786893436e-11, 
    -1.9292834658422995e-11, -1.9239776756220035e-11, 
    -1.9170593584865064e-11, -1.9086505024190184e-11, -1.898841036196918e-11, 
    -1.8877006634920594e-11, -1.8752976972067215e-11, 
    -1.8617226029531576e-11, -1.8471112471883437e-11, -1.831665020731553e-11, 
    -1.8156627617869699e-11, -1.7994647999674813e-11, 
    -1.7835065410619873e-11, -1.7682798415693817e-11, 
    -1.7543061988695561e-11, -1.742107274834065e-11, -1.732167508341348e-11, 
    -1.7249002900940053e-11, -1.720616509664526e-11, -1.7195012974577602e-11, 
    -1.7215982739485942e-11, -1.7268060491033786e-11, 
    -1.7348843698155838e-11, -1.7454726685811287e-11, 
    -1.7581159910514461e-11, -1.7723019678831769e-11, 
    -1.7874994857774068e-11, -1.8032018564555447e-11, 
    -1.8189676134963323e-11, -1.8344565889072877e-11, 
    -1.8494577941429569e-11, -1.8639086425233173e-11, -1.877899055186197e-11, 
    -1.8916657044217767e-11, -1.9055713940549487e-11, 
    -1.9200758065997937e-11, -1.9356955205886746e-11, 
    -1.9529625172631327e-11, -1.9723797775753772e-11, 
    -1.9943779642350974e-11, -2.0192776529988335e-11, 
    -2.0472620897486162e-11, -2.078353378913619e-11, -2.1124011220848408e-11, 
    -2.1490781564042243e-11, -2.1878856610962068e-11, 
    -2.2281633202905093e-11, -2.2691077477905395e-11, 
    -2.3097948625059564e-11, -2.3492070866463957e-11, 
    -2.3862644870389513e-11, -2.4198608238559964e-11, 
    -2.4488998870446105e-11, -2.4723366820023307e-11, 
    -2.4892168249214864e-11, -2.4987163124114043e-11, 
    -2.5001758304484387e-11, -2.4931346451811068e-11, 
    -2.4773516860431699e-11, -2.4528230244303866e-11, 
    -2.4197871536344778e-11, -2.3787218275367117e-11, 
    -2.3303298890057409e-11, -2.27551907241459e-11, -2.2153719794889795e-11, 
    -2.1511123657233083e-11, -2.0840668386096296e-11, 
    -2.0156266151550194e-11, -1.9472049096962769e-11, -1.880201647103398e-11, 
    -1.8159651106769728e-11, -1.7557574451608455e-11, 
    -1.7007239393727076e-11, -1.6518655044651889e-11, 
    -1.6100131457217743e-11, -1.5758069664810092e-11, 
    -1.5496780590055939e-11, -1.5318357435171058e-11, 
    -1.5222584239243884e-11, -1.5206919140210245e-11, 
    -1.5266544739118365e-11, -1.5394489290385759e-11, 
    -1.5581847665261455e-11, -1.5818089533426015e-11, 
    -1.6091454442625084e-11, -1.6389420475159051e-11, 
    -1.6699249822045828e-11, -1.7008539960685597e-11, 
    -1.7305798870850499e-11, -1.7580988559408242e-11, 
    -1.7825987273728642e-11, -1.8034932269366945e-11, 
    -1.8204451240044456e-11, -1.8333712347305607e-11, 
    -1.8424310887787215e-11, -1.8479989676997142e-11, 
    -1.8506205400259773e-11, -1.8509588980150794e-11, 
    -1.8497323381155688e-11, -1.8476500017434673e-11, 
    -1.8453515105794935e-11, -1.8433531791354151e-11, 
    -1.8420087282525717e-11, -1.8414858451144788e-11, 
    -1.8417597783898489e-11, -1.8426272169679344e-11, 
    -1.8437361086060257e-11, -1.8446304990682897e-11, 
    -1.8448058031167531e-11, -1.8437681588603082e-11, 
    -1.8410951335369342e-11, -1.8364889005915084e-11, 
    -1.8298198431018951e-11, -1.8211547862125742e-11, 
    -1.8107686129814072e-11, -1.7991353331171723e-11, 
    -1.7869034689800986e-11, -1.7748538348531908e-11, 
    -1.7638455287431608e-11, -1.7547540886580903e-11, 
    -1.7484056329390735e-11, -1.7455144931223847e-11, 
    -1.7466269284765544e-11, -1.752076314782617e-11, -1.7619526138361862e-11, 
    -1.7760868755622318e-11, -1.7940535093899117e-11, 
    -1.8151880801778768e-11, -1.8386217304021379e-11, 
    -1.8633236716648699e-11, -1.8881581386310644e-11, 
    -1.9119443524417628e-11, -1.9335226719505958e-11, 
    -1.9518162570728337e-11, -1.9658908756446065e-11, 
    -1.9750091596063358e-11, -1.9786727612518311e-11, 
    -1.9766528278211658e-11, -1.9690084394257146e-11, 
    -1.9560884367826996e-11, -1.9385205245258055e-11, 
    -1.9171855665431591e-11, -1.8931787655026743e-11, 
    -1.8677607247989086e-11, -1.8423004941545349e-11, -1.818209062500506e-11, 
    -1.7968725100261177e-11, -1.7795832404540288e-11, 
    -1.7674737529745644e-11, -1.761452738312095e-11, -1.7621531126847447e-11, 
    -1.7698872909997482e-11, -1.7846190275487274e-11, 
    -1.8059478999331289e-11, -1.8331158970289197e-11, 
    -1.8650287325970588e-11, -1.9002992435942352e-11, 
    -1.9373048248354218e-11, -1.9742624437263793e-11, 
    -2.0093107881686211e-11, -2.0406014308628324e-11, 
    -2.0663872427919926e-11, -2.0851097809034142e-11, 
    -2.0954731452364643e-11, -2.0965093483449642e-11, 
    -2.0876234033851333e-11, -2.0686260117672098e-11, 
    -2.0397434947909003e-11, -2.0016148794633636e-11, 
    -1.9552678359858907e-11, -1.9020830402880528e-11, 
    -1.8437402875855354e-11, -1.7821552404334285e-11, 
    -1.7193988383044713e-11, -1.6576144233718521e-11, 
    -1.5989190490954081e-11, -1.5453079116076015e-11, 
    -1.4985571728014915e-11, -1.4601341803629593e-11, 
    -1.4311173865556317e-11, -1.4121389742541664e-11, 
    -1.4033465084356208e-11, -1.4043950109530615e-11, 
    -1.4144655993897816e-11, -1.4323156495007996e-11, 
    -1.4563506342189653e-11, -1.4847227350657434e-11, -1.515436612960831e-11, 
    -1.5464674483774666e-11, -1.5758741131715164e-11, 
    -1.6019039801841083e-11, -1.6230815661567661e-11, -1.638277086118356e-11, 
    -1.6467497921230956e-11, -1.6481684427284611e-11, 
    -1.6426056283815565e-11, -1.6305123685107048e-11, -1.612671492821729e-11, 
    -1.5901397147377875e-11, -1.5641765240087798e-11, -1.536170285011245e-11, 
    -1.507561760655712e-11, -1.4797715336737362e-11, -1.4541338246412042e-11, 
    -1.4318398220527414e-11, -1.4138925358434768e-11, 
    -1.4010752214983529e-11, -1.3939321778313961e-11, 
    -1.3927653242683859e-11, -1.397639076068565e-11, -1.4083973916934073e-11, 
    -1.4246886585404557e-11, -1.4459949660663401e-11, 
    -1.4716622055624013e-11, -1.5009327329170545e-11, 
    -1.5329744624883178e-11, -1.5669093656995458e-11, 
    -1.6018382765361567e-11, -1.6368655795535041e-11, 
    -1.6711219567538825e-11, -1.703788025102276e-11, -1.7341202847412966e-11, 
    -1.7614758418991338e-11, -1.7853391336737144e-11, 
    -1.8053457907675746e-11, -1.8213018438103369e-11, 
    -1.8331958761471885e-11, -1.8412005702852628e-11, 
    -1.8456615999436536e-11, -1.8470719225855146e-11, 
    -1.8460335801603102e-11, -1.8432067251891042e-11, 
    -1.8392534365605946e-11, -1.8347760253181916e-11, 
    -1.8302625598054421e-11, -1.8260394016170326e-11, 
    -1.8222431450761571e-11, -1.8188085450294155e-11, 
    -1.8154827778942694e-11, -1.8118592018361771e-11, -1.807433266901286e-11, 
    -1.801670218369824e-11, -1.7940837468037308e-11, -1.7843080146578748e-11, 
    -1.7721669123950593e-11, -1.7577188995463288e-11, 
    -1.7412832251783575e-11, -1.7234330853370934e-11, 
    -1.7049649830058118e-11, -1.6868375479796674e-11, 
    -1.6700931894100383e-11, -1.6557642010678771e-11, -1.64477886575707e-11, 
    -1.6378720639388296e-11, -1.6355159187336352e-11,
  // Sqw-F(3, 0-1999)
    0.057087479352590245, 0.057005779208843935, 0.05676222017799646, 
    0.056361352427440038, 0.055810518367261384, 0.055119509860033333, 
    0.054300124566273554, 0.053365653711247948, 0.052330337549663257, 
    0.051208825582646285, 0.050015676138979823, 0.048764924576258584, 
    0.047469741676870014, 0.046142194620777996, 0.04479311316233156, 
    0.043432054309131572, 0.042067350814888604, 0.040706222902308686, 
    0.039354929320693302, 0.038018933304735991, 0.036703061102578448, 
    0.035411635051258904, 0.034148569028998751, 0.032917420695251193, 
    0.031721401395884946, 0.030563350194420628, 0.029445682597255423, 
    0.028370326819873826, 0.027338660812511937, 0.026351461907654701, 
    0.025408878258040699, 0.024510427725136726, 0.023655026119294906, 
    0.022841043204047604, 0.02206638206310391, 0.021328575536286816, 
    0.020624892536686052, 0.019952447090029479, 0.019308303699966282, 
    0.018689573888875877, 0.018093500231808342, 0.017517525662462896, 
    0.016959347116344357, 0.016416953590645839, 0.015888649413923248, 
    0.015373063955380227, 0.014869149221013038, 0.014376166852956536, 
    0.013893666037432863, 0.013421453790848055, 0.012959559069777273, 
    0.012508192157274322, 0.012067700817457984, 0.011638524772523589, 
    0.011221150122404664, 0.010816065373422277, 0.010423720742828348, 
    0.010044492337245142, 0.009678652645721807, 0.0093263485319619727, 
    0.0089875875558627569, 0.0086622330153048564, 0.0083500076014053921, 
    0.008050505041328081, 0.0077632086064949009, 0.0074875149369301027, 
    0.0072227613170122874, 0.0069682543673725041, 0.006723298111471222, 
    0.0064872195362181287, 0.0062593900788952264, 0.0060392419062751685, 
    0.0058262783617332482, 0.0056200784897935605, 0.0054202960504004857, 
    0.0052266538573651402, 0.0050389345777303602, 0.0048569692876729662, 
    0.0046806250908295799, 0.0045097929800213613, 0.0043443768927662442, 
    0.0041842846154402404, 0.0040294208759027077, 0.0038796826729429316, 
    0.003734956657441761, 0.0035951182258318801, 0.0034600319171346709, 
    0.0033295527118615293, 0.0032035278944035307, 0.0030817992339016707, 
    0.0029642053350251996, 0.0028505840871642053, 0.0027407751841187185, 
    0.0026346226923405357, 0.0025319776196430096, 0.0024327003908276345, 
    0.0023366630884052702, 0.0022437512818506643, 0.0021538652602101321, 
    0.0020669205068067327, 0.0019828473104830211, 0.0019015894878695553, 
    0.0018231022832530491, 0.0017473496021512551, 0.0016743008076176599, 
    0.0016039273536030301, 0.0015361995412086903, 0.0014710836607962283, 
    0.0014085397303847196, 0.0013485199674313937, 0.0012909680481700877, 
    0.0012358191277679188, 0.0011830005257535147, 0.0011324329316962627, 
    0.0010840319595414359, 0.0010377098751912772, 0.00099337733754960755, 
    0.00095094502283580066, 0.00091032503906620494, 0.00087143207596460722, 
    0.00083418427012356357, 0.00079850379268660526, 0.00076431718576939415, 
    0.00073155548463076352, 0.00070015416681019004, 0.00067005296924159874, 
    0.00064119561187060703, 0.00061352946316495835, 0.00058700517993267903, 
    0.00056157635106061834, 0.00053719917155033148, 0.00051383216870601865, 
    0.00049143599580954824, 0.00046997329989052457, 0.00044940865973747059, 
    0.0004297085792708129, 0.00041084151147007837, 0.00039277788103991797, 
    0.00037549007147188995, 0.00035895234504647734, 0.00034314067265362738, 
    0.00032803246315611282, 0.00031360619757928471, 0.00029984098933181634, 
    0.00028671610543321073, 0.0002742104931293763, 0.00026230235976519188, 
    0.00025096885074027967, 0.00024018586119507911, 0.00022992800309201374, 
    0.00022016873257851694, 0.00021088062530691008, 0.00020203577205743801, 
    0.00019360625550915347, 0.00018556466261609981, 0.00017788458627587288, 
    0.00017054107451116841, 0.00016351099421641597, 0.00015677328814043536, 
    0.00015030911643897232, 0.00014410188612091782, 0.00013813718159340354, 
    0.00013240261629964914, 0.00012688762871401686, 0.00012158324584017948, 
    0.00011648183446369238, 0.00011157685567882458, 0.00010686263273391623, 
    0.00010233413706110894, 9.7986793312792485e-05, 9.3816301824540198e-05, 
    8.981847629888667e-05, 8.5989095431372961e-05, 8.2323769181956238e-05, 
    7.8817822770837559e-05, 7.5466203568610128e-05, 7.2263417276826965e-05, 
    6.9203499781050876e-05, 6.6280029677243772e-05, 6.3486183858016737e-05, 
    6.0814835044237903e-05, 5.8258686256457046e-05, 5.5810433486712565e-05, 
    5.3462944776525145e-05, 5.120944193936108e-05, 4.9043670543573938e-05, 
    4.696004456564944e-05, 4.4953754234179874e-05, 4.3020828758531763e-05, 
    4.1158149516995865e-05, 3.936341345079279e-05, 3.7635050456083066e-05, 
    3.597210210610081e-05, 3.4374071772600307e-05, 3.2840757950165959e-05, 
    3.1372083237310799e-05, 2.9967931018761037e-05, 2.86280005508072e-05, 
    2.7351689070476009e-05, 2.6138006975167784e-05, 2.498552930680508e-05, 
    2.3892383970475032e-05, 2.2856274529816383e-05, 2.1874533214406535e-05, 
    2.0944198055487556e-05, 2.0062106897871169e-05, 1.922500043314342e-05, 
    1.8429626351360286e-05, 1.7672837175216909e-05, 1.6951675270180285e-05, 
    1.6263439843237078e-05, 1.5605732366115761e-05, 1.4976478677375041e-05, 
    1.4373927908042381e-05, 1.379663019477887e-05, 1.3243396749042767e-05, 
    1.2713247100917395e-05, 1.220534912298951e-05, 1.1718957691130048e-05, 
    1.1253357543257224e-05, 1.0807815096202991e-05, 1.0381542778132569e-05, 
    9.9736779708015247e-06, 9.5832771022032163e-06, 9.2093239521652465e-06, 
    8.8507499803336787e-06, 8.5064635646352131e-06, 8.1753845099222445e-06, 
    7.8564800575728738e-06, 7.5487988627132195e-06, 7.251499932792784e-06, 
    6.9638742519787282e-06, 6.6853576513659964e-06, 6.4155343391188277e-06, 
    6.1541313004712507e-06, 5.9010044624441021e-06, 5.6561180543890333e-06, 
    5.4195189678593431e-06, 5.1913081230084488e-06, 4.9716108947222327e-06, 
    4.7605485553802132e-06, 4.5582124776352553e-06, 4.3646425346238864e-06, 
    4.1798107670860102e-06, 4.0036109824087894e-06, 3.8358545381746159e-06, 
    3.6762721628528778e-06, 3.5245213007007318e-06, 3.3801981508309369e-06, 
    3.2428533174894176e-06, 3.1120098092954281e-06, 2.9871820311690086e-06, 
    2.8678944084060728e-06, 2.7536983726974702e-06, 2.6441866186966537e-06, 
    2.5390037980018205e-06, 2.4378531324086627e-06, 2.3404987748984549e-06, 
    2.2467640894500306e-06, 2.1565263285428615e-06, 2.0697084275248496e-06, 
    1.9862687897158433e-06, 1.9061899935267733e-06, 1.8294673194313995e-06, 
    1.7560978841060707e-06, 1.6860710080340538e-06, 1.6193602572332776e-06, 
    1.5559174179472634e-06, 1.4956685037353708e-06, 1.4385117708328502e-06, 
    1.3843176304589159e-06, 1.3329302920223796e-06, 1.2841709363415581e-06, 
    1.237842193110039e-06, 1.193733669919792e-06, 1.1516282485473447e-06, 
    1.1113088265200919e-06, 1.0725651463663586e-06, 1.0352003291172034e-06, 
    9.990367245051604e-07, 9.6392071447969293e-07, 9.2972616455001979e-07, 
    8.9635630618639204e-07, 8.6374394755344969e-07, 8.3185003621103757e-07, 
    8.0066072451943263e-07, 7.7018320049414641e-07, 7.4044063408776389e-07, 
    7.1146664145273964e-07, 6.8329968568549138e-07, 6.5597781114545358e-07, 
    6.2953405595485235e-07, 6.0399280947154252e-07, 5.7936728946281768e-07, 
    5.5565821442268169e-07, 5.3285365104216257e-07, 5.1092993057276187e-07, 
    4.898534580399392e-07, 4.6958318717456594e-07, 4.5007350491626467e-07, 
    4.3127726071598339e-07, 4.1314868816477414e-07, 3.9564599517803918e-07, 
    3.7873344241135858e-07, 3.6238278206391544e-07, 3.4657398806262033e-07, 
    3.3129526783112672e-07, 3.1654240298750148e-07, 3.0231751586803678e-07, 
    2.8862739933286822e-07, 2.7548157413721973e-07, 2.6289025174414936e-07, 
    2.5086237768894532e-07, 2.3940391400447911e-07, 2.2851648845982621e-07, 
    2.1819649825389139e-07, 2.084347084237336e-07, 1.9921633747699748e-07, 
    1.9052157750945307e-07, 1.8232646013703007e-07, 1.7460395435914055e-07, 
    1.6732517252602076e-07, 1.6046056357999403e-07, 1.5398098958174646e-07, 
    1.4785860685995796e-07, 1.4206750474448841e-07, 1.3658408635980959e-07, 
    1.3138720506145739e-07, 1.2645809196550228e-07, 1.2178012455851399e-07, 
    1.173384915026899e-07, 1.1311980742267722e-07, 1.0911172366347299e-07, 
    1.0530257094369333e-07, 1.0168105804820816e-07, 9.8236040690335908e-08, 
    9.4956365923188893e-08, 9.1830791905801185e-08, 8.884797875805014e-08, 
    8.5996544425833029e-08, 8.326517769035028e-08, 8.0642799710556473e-08, 
    7.811876348965188e-08, 7.5683079275602166e-08, 7.3326651379848084e-08, 
    7.1041510366360349e-08, 6.8821022749862074e-08, 6.6660060318133077e-08, 
    6.4555111586803452e-08, 6.2504320426854655e-08, 6.0507440268900107e-08, 
    5.85656976515241e-08, 5.6681564687214874e-08, 5.485844744568829e-08, 
    5.3100304176123107e-08, 5.1411214807955789e-08, 4.9794928765592285e-08, 
    4.8254422910984364e-08, 4.6791502726355137e-08, 4.5406478975029806e-08, 
    4.4097947048746086e-08, 4.2862688727257722e-08, 4.1695705309365212e-08, 
    4.0590379582058423e-08, 3.9538751552926595e-08, 3.8531882724325388e-08, 
    3.7560275435881995e-08, 3.6614310295063714e-08, 3.5684664957561082e-08, 
    3.4762682776679102e-08, 3.3840667988175524e-08, 3.291209493008476e-08, 
    3.1971729658802705e-08, 3.1015672357425424e-08, 3.0041335744290003e-08, 
    2.9047378658463749e-08, 2.8033613324557899e-08, 2.700090169627622e-08, 
    2.5951050294634152e-08, 2.4886706719504668e-08, 2.3811254939627418e-08, 
    2.2728702860549994e-08, 2.1643554044046516e-08, 2.0560657330562791e-08, 
    1.9485031728346987e-08, 1.8421669805783093e-08, 1.7375328396671456e-08, 
    1.6350320958878834e-08, 1.5350329026382473e-08, 1.4378251400049249e-08, 
    1.3436107548288817e-08, 1.2525007593712986e-08, 1.1645194326932008e-08, 
    1.0796155220730393e-08, 9.9767942520399072e-09, 9.1856464647270568e-09, 
    8.4211128059443707e-09, 7.6816905183456297e-09, 6.9661745583619733e-09, 
    6.2738093038181003e-09, 5.6043756972289738e-09, 4.9582071532608596e-09, 
    4.3361358667510702e-09, 3.7393796397259203e-09, 3.169385466896321e-09, 
    2.6276505242879822e-09, 2.1155420038927857e-09, 1.6341356694137718e-09, 
    1.1840885941873536e-09, 7.6555597981991644e-10, 3.7815530291342629e-10, 
    2.0975523575975398e-11, -3.0737578847480307e-10, -6.0869711361956299e-10, 
    -8.8510023170648608e-10, -1.1389099467122316e-09, 
    -1.3725645416568877e-09, -1.5885226966846153e-09, 
    -1.7891806270942348e-09, -1.9768011075089744e-09, 
    -2.1534554289085855e-09, -2.3209784889705763e-09, 
    -2.4809375324782495e-09, -2.6346149346711234e-09, 
    -2.7830054701240028e-09, -2.9268278719452572e-09, 
    -3.0665498754953727e-09, -3.202424473084466e-09, -3.3345342056610133e-09, 
    -3.4628390008594081e-09, -3.5872227482065322e-09, -3.707533597414646e-09, 
    -3.8236138338997534e-09, -3.935316302732683e-09, -4.0425062127772819e-09, 
    -4.1450488791508886e-09, -4.2427860635721685e-09, 
    -4.3355049447814682e-09, -4.422905189418716e-09, -4.5045699244957675e-09, 
    -4.5799465547226725e-09, -4.6483423826006765e-09, 
    -4.7089388318202093e-09, -4.7608258534106529e-09, -4.803056057379407e-09, 
    -4.8347154193412109e-09, -4.8550053499591219e-09, 
    -4.8633287457814219e-09, -4.8593717053912746e-09, 
    -4.8431720642442331e-09, -4.8151667783923928e-09, -4.776211735483784e-09, 
    -4.7275702697693343e-09, -4.6708695900122407e-09, 
    -4.6080277380424718e-09, -4.541156685812564e-09, -4.4724496482055612e-09, 
    -4.4040621478105952e-09, -4.3379968899813575e-09, 
    -4.2760015937173451e-09, -4.219487445123649e-09, -4.1694731894509022e-09, 
    -4.1265572274668447e-09, -4.0909171272309653e-09, 
    -4.0623337559335087e-09, -4.0402351398568357e-09, 
    -4.0237544941605603e-09, -4.0117963823896137e-09, 
    -4.0031057495510685e-09, -3.9963354305833058e-09, 
    -3.9901092184786066e-09, -3.9830787669897516e-09, 
    -3.9739738418985481e-09, -3.9616460126274694e-09, 
    -3.9451063049577135e-09, -3.9235570395475228e-09, 
    -3.8964178018951037e-09, -3.8633447292509679e-09, 
    -3.8242419899925326e-09, -3.7792637566825159e-09, 
    -3.7288053941055546e-09, -3.6734827122396518e-09, 
    -3.6140992796890304e-09, -3.551602750606615e-09, -3.4870325601257426e-09, 
    -3.4214623213537355e-09, -3.3559412997256113e-09, 
    -3.2914395504841602e-09, -3.2288012801014775e-09, 
    -3.1687101709056528e-09, -3.1116693544546845e-09, 
    -3.0579970075098845e-09, -3.0078371349171041e-09, 
    -2.9611833948943689e-09, -2.9179127370071151e-09, -2.877824670348534e-09, 
    -2.8406818663145278e-09, -2.8062477987211006e-09, 
    -2.7743179677443643e-09, -2.7447420307620678e-09, 
    -2.7174354361255642e-09, -2.6923801585729216e-09, 
    -2.6696153824216563e-09, -2.6492196464070124e-09, 
    -2.6312869567713573e-09, -2.6158994281408869e-09, 
    -2.6030995469922515e-09, -2.5928648424770351e-09, 
    -2.5850876624110095e-09, -2.5795620795281049e-09, 
    -2.5759795167735237e-09, -2.5739336051457929e-09, -2.572934210998223e-09, 
    -2.5724293128990005e-09, -2.5718329831651312e-09, 
    -2.5705567263273321e-09, -2.5680414640745081e-09, 
    -2.5637871189536855e-09, -2.557377387455156e-09, -2.5484977362105709e-09, 
    -2.5369457761622234e-09, -2.5226338289240625e-09, 
    -2.5055847440310707e-09, -2.4859223700548144e-09, 
    -2.4638587231745685e-09, -2.4396796336330875e-09, 
    -2.4137305624302977e-09, -2.3864034456511077e-09, 
    -2.3581250011133078e-09, -2.329345964927808e-09, -2.3005305831983458e-09, 
    -2.2721452174314942e-09, -2.2446452936416643e-09, 
    -2.2184600405921513e-09, -2.1939752815480007e-09, 
    -2.1715150564753672e-09, -2.151323681730527e-09, -2.1335500012431155e-09, 
    -2.1182360373121759e-09, -2.1053116963238768e-09, 
    -2.0945969830735666e-09, -2.0858121676095401e-09, 
    -2.0785957062884587e-09, -2.0725286162284838e-09, 
    -2.0671634824240386e-09, -2.0620555022101906e-09, -2.056793025684109e-09, 
    -2.0510247491006484e-09, -2.0444813947016794e-09, 
    -2.0369900365584433e-09, -2.028480178512673e-09, -2.0189812277689726e-09, 
    -2.0086121278543646e-09, -1.9975642547564846e-09, 
    -1.9860794999828096e-09, -1.9744255511794466e-09, 
    -1.9628707251687193e-09, -1.9516603337217994e-09, 
    -1.9409965781857264e-09, -1.9310232467238921e-09, 
    -1.9218162729387304e-09, -1.9133803781580374e-09, 
    -1.9056517991132501e-09, -1.8985063508226898e-09, 
    -1.8917720386430813e-09, -1.8852448326774978e-09, 
    -1.8787064019867759e-09, -1.8719423179400378e-09, 
    -1.8647595461266051e-09, -1.8570018761397476e-09, 
    -1.8485625107433168e-09, -1.8393928633510947e-09, -1.829507280686432e-09, 
    -1.8189833159557824e-09, -1.8079577501882772e-09, 
    -1.7966186003310423e-09, -1.7851937647825473e-09, 
    -1.7739369599420821e-09, -1.7631120060772614e-09, -1.752976285511939e-09, 
    -1.74376459280117e-09, -1.7356741965110493e-09, -1.728852202381966e-09, 
    -1.7233858441583569e-09, -1.7192964753086785e-09, 
    -1.7165374995207739e-09, -1.714996571694239e-09, -1.7145018536287816e-09, 
    -1.7148321311234074e-09, -1.7157300563069615e-09, -1.71691784014192e-09, 
    -1.7181142213758652e-09, -1.7190516669912957e-09, 
    -1.7194924070939191e-09, -1.7192422260141197e-09, 
    -1.7181607587087891e-09, -1.7161675745054417e-09, 
    -1.7132433918135624e-09, -1.7094264610501667e-09, 
    -1.7048043057771689e-09, -1.699501714426433e-09, -1.6936659943669486e-09, 
    -1.6874509738040843e-09, -1.681001135781784e-09, -1.6744374334885176e-09, 
    -1.6678459393863847e-09, -1.6612703663019065e-09, 
    -1.6547088721853968e-09, -1.6481153676942902e-09, 
    -1.6414048654270119e-09, -1.6344623106842807e-09, 
    -1.6271538207186181e-09, -1.6193393672129876e-09, 
    -1.6108856316844625e-09, -1.6016781372594987e-09, 
    -1.5916315928566902e-09, -1.5806979475373294e-09, 
    -1.5688715017812328e-09, -1.5561910400732302e-09, 
    -1.5427388300828086e-09, -1.5286368088408682e-09, 
    -1.5140401861020149e-09, -1.4991290772643226e-09, -1.484098617845539e-09, 
    -1.4691483370697196e-09, -1.4544713491824846e-09, 
    -1.4402441896622277e-09, -1.4266177806727911e-09, -1.413710270340067e-09, 
    -1.4016019937313255e-09, -1.3903330321236379e-09, 
    -1.3799032782942058e-09, -1.3702751005934626e-09, 
    -1.3613781522796659e-09, -1.3531160184085227e-09, 
    -1.3453740235687705e-09, -1.3380276699013376e-09, 
    -1.3309509278987574e-09, -1.3240239214980843e-09, 
    -1.3171393431995934e-09, -1.3102073476360214e-09, 
    -1.3031585938691468e-09, -1.2959454629553018e-09, 
    -1.2885414459288817e-09, -1.2809390186285868e-09, -1.273146209609926e-09, 
    -1.2651823708969781e-09, -1.2570733985764616e-09, 
    -1.2488469958656319e-09, -1.240528165166832e-09, -1.2321354086649546e-09, 
    -1.2236777626378145e-09, -1.2151530223989091e-09, 
    -1.2065470889603494e-09, -1.1978346599434474e-09, 
    -1.1889810684441235e-09, -1.1799453039856734e-09, 
    -1.1706838456034063e-09, -1.1611551681981427e-09, 
    -1.1513244362102466e-09, -1.1411681187208959e-09, 
    -1.1306779671631356e-09, -1.119864117993026e-09, -1.1087568586812424e-09, 
    -1.097406998093074e-09, -1.0858846047975499e-09, -1.0742763676977559e-09, 
    -1.0626816275465762e-09, -1.0512075770637511e-09, 
    -1.0399639153486111e-09, -1.0290575144387457e-09, 
    -1.0185874124148654e-09, -1.008640575760692e-09, -9.9928857782169001e-10, 
    -9.9058540411930586e-10, -9.8256627130313266e-10, 
    -9.7524749315915197e-10, -9.6862708785266524e-10, 
    -9.6268605128919086e-10, -9.5739001052675914e-10, 
    -9.5269115283136138e-10, -9.4853025646294587e-10, 
    -9.4483883833733411e-10, -9.4154128755324689e-10, 
    -9.3855707460608626e-10, -9.3580300069832856e-10, 
    -9.3319553935314127e-10, -9.3065318795090191e-10, 
    -9.2809889126202362e-10, -9.2546233875729431e-10, 
    -9.2268215375135509e-10, -9.1970773622317913e-10, 
    -9.1650074138467489e-10, -9.1303597512477941e-10, 
    -9.0930167531934587e-10, -9.0529906708410589e-10, 
    -9.0104124820060755e-10, -8.9655135978701095e-10, 
    -8.9186025688027517e-10, -8.8700373387983298e-10, 
    -8.8201963274026742e-10, -8.7694496021996567e-10, 
    -8.7181339658700477e-10, -8.6665329100500426e-10, -8.614864619235826e-10, 
    -8.5632780712459316e-10, -8.5118584524658671e-10, -8.460640182144594e-10, 
    -8.409626709459633e-10, -8.3588136726747586e-10, -8.3082132020482204e-10, 
    -8.2578752717481493e-10, -8.207903825161137e-10, -8.1584645294054098e-10, 
    -8.1097835431719801e-10, -8.062136322748876e-10, -8.0158277575581818e-10, 
    -7.9711655093330734e-10, -7.9284298367974962e-10, 
    -7.8878426794522146e-10, -7.8495400159865102e-10, 
    -7.8135501611232394e-10, -7.7797809002884049e-10, 
    -7.7480162119680361e-10, -7.7179235972729607e-10, 
    -7.6890706644396167e-10, -7.6609500416527845e-10, 
    -7.6330095952234588e-10, -7.6046859913041845e-10, 
    -7.5754383759667605e-10, -7.5447801607309118e-10, 
    -7.5123063146038697e-10, -7.4777153312692685e-10, 
    -7.4408240557589352e-10, -7.4015758991013021e-10, -7.360041567046828e-10, 
    -7.3164135151847746e-10, -7.2709940560494731e-10, 
    -7.2241787475805062e-10, -7.1764350580935458e-10, 
    -7.1282782301745408e-10, -7.0802445702196763e-10, 
    -7.0328640422189877e-10, -6.9866326299373299e-10, -6.941986793242058e-10, 
    -6.899280245645438e-10, -6.8587655861980685e-10, -6.8205811306474375e-10, 
    -6.7847446779902572e-10, -6.7511542175094739e-10, -6.719596493464991e-10, 
    -6.6897620157867009e-10, -6.6612663025489884e-10, 
    -6.6336749501214711e-10, -6.6065312615958309e-10, 
    -6.5793832979405809e-10, -6.5518090747836412e-10, 
    -6.5234370743188588e-10, -6.4939615117697985e-10, 
    -6.4631509238516448e-10, -6.4308509112613469e-10, 
    -6.3969808062353971e-10, -6.361526550673247e-10, -6.3245304723619215e-10, 
    -6.2860804386794237e-10, -6.2462990134750453e-10, 
    -6.2053348703641397e-10, -6.163355882996354e-10, -6.1205447761121248e-10, 
    -6.0770963963879723e-10, -6.0332164264171513e-10, 
    -5.9891196033447606e-10, -5.9450274671085889e-10, 
    -5.9011641557221778e-10, -5.8577503432416855e-10, 
    -5.8149951417413194e-10, -5.7730869320682766e-10, 
    -5.7321833761410822e-10, -5.6924029700154181e-10, 
    -5.6538182036232548e-10, -5.6164525483921395e-10, 
    -5.5802814585118601e-10, -5.5452383091933449e-10, 
    -5.5112244605160473e-10, -5.4781233830325929e-10, 
    -5.4458167549671101e-10, -5.4142015602248203e-10, 
    -5.3832054749904633e-10, -5.352799649847415e-10, -5.3230063244356466e-10, 
    -5.2939008676137506e-10, -5.2656075389490029e-10, 
    -5.2382891876735818e-10, -5.212131758852434e-10, -5.1873254148557106e-10, 
    -5.1640436679633923e-10, -5.1424231924392049e-10, 
    -5.1225457646747763e-10, -5.1044247764359511e-10, 
    -5.0879970405400334e-10, -5.0731211316719637e-10, 
    -5.0595820058552995e-10, -5.0471018271577176e-10, 
    -5.0353552818922631e-10, -5.0239886152602625e-10, -5.012639986716954e-10, 
    -5.0009598469406835e-10, -4.9886291150871975e-10, -4.975374561339496e-10, 
    -4.9609795315523096e-10, -4.9452903048503821e-10, 
    -4.9282178501243744e-10, -4.9097356273521461e-10, 
    -4.8898741729306971e-10, -4.8687140162646893e-10, 
    -4.8463773944979343e-10, -4.8230203770460696e-10, -4.798825625306126e-10, 
    -4.7739965446664763e-10, -4.7487523499496194e-10, 
    -4.7233240730128669e-10, -4.6979505471837216e-10, 
    -4.6728740339227208e-10, -4.6483344681265276e-10, 
    -4.6245623622560849e-10, -4.6017698803745505e-10, -4.580140649091136e-10, 
    -4.5598189135578775e-10, -4.5408989345646177e-10, 
    -4.5234158154837206e-10, -4.5073389029340894e-10, 
    -4.4925685834354082e-10, -4.478937670069812e-10, -4.4662170990118291e-10, 
    -4.4541264004109003e-10, -4.4423480391599116e-10, -4.430544999882097e-10, 
    -4.4183801516625968e-10, -4.4055361688229122e-10, 
    -4.3917343962027076e-10, -4.3767513711859962e-10, 
    -4.3604317691371347e-10, -4.3426968244617145e-10, 
    -4.3235477968964835e-10, -4.3030643208703061e-10, 
    -4.2813978838439987e-10, -4.2587612051887434e-10, 
    -4.2354142163291733e-10, -4.2116483276367767e-10, 
    -4.1877695553677912e-10, -4.1640822984982292e-10, 
    -4.1408744994390095e-10, -4.1184054312874488e-10, 
    -4.0968960977319776e-10, -4.0765231150752574e-10, 
    -4.0574152906101562e-10, -4.0396532312215345e-10, 
    -4.0232704962997837e-10, -4.008256589800862e-10, -3.9945602195465559e-10, 
    -3.9820929802488667e-10, -3.9707325425912325e-10, 
    -3.9603259540135445e-10, -3.9506925738671783e-10, 
    -3.9416274551867594e-10, -3.9329053538357714e-10, 
    -3.9242862533522537e-10, -3.9155220214801758e-10, 
    -3.9063650759464643e-10, -3.896577964666702e-10, -3.8859441695896373e-10, 
    -3.8742784539236981e-10, -3.861436703422989e-10, -3.8473231800554669e-10, 
    -3.8318957112193334e-10, -3.8151669886197957e-10, 
    -3.7972025337409452e-10, -3.7781153159689973e-10, 
    -3.7580576878394854e-10, -3.7372112095945703e-10, 
    -3.7157759204788417e-10, -3.6939593355722012e-10, 
    -3.6719668430464091e-10, -3.6499934351462987e-10, 
    -3.6282176374357856e-10, -3.6067970449858981e-10, 
    -3.5858661607810395e-10, -3.5655348556964138e-10, 
    -3.5458881536632759e-10, -3.526985761739539e-10, -3.5088620674640127e-10, 
    -3.4915254817750197e-10, -3.4749580332766131e-10, 
    -3.4591146878513522e-10, -3.4439238218564454e-10, 
    -3.4292881097997493e-10, -3.4150877692954593e-10, 
    -3.4011849283996489e-10, -3.3874305781723378e-10, 
    -3.3736728723404024e-10, -3.3597672864140483e-10, 
    -3.3455867380910665e-10, -3.3310320336303581e-10, 
    -3.3160402730332005e-10, -3.3005913303587067e-10, -3.284710546333951e-10, 
    -3.2684678785391581e-10, -3.2519724827385467e-10, 
    -3.2353637788866295e-10, -3.2187987679526032e-10, 
    -3.2024374073638393e-10, -3.1864267772983367e-10, 
    -3.1708860735048058e-10, -3.1558932750844959e-10, 
    -3.1414756961470545e-10, -3.1276045721894588e-10, 
    -3.1141951008365907e-10, -3.1011114449991908e-10, 
    -3.0881770177741097e-10, -3.0751884002899722e-10, -3.061932577895921e-10, 
    -3.048204999465739e-10, -3.0338276780836804e-10, -3.0186648307888918e-10, 
    -3.0026355292564813e-10, -2.985721268625389e-10, -2.9679686449440942e-10, 
    -2.949486209349243e-10, -2.9304367281951363e-10, -2.9110245806949839e-10, 
    -2.8914808007664775e-10, -2.8720459948068843e-10, 
    -2.8529537075388315e-10, -2.8344148439389907e-10, 
    -2.8166053793660614e-10, -2.7996570781891889e-10, 
    -2.7836528504375721e-10, -2.7686257206978424e-10, 
    -2.7545619935427994e-10, -2.7414070590993014e-10, 
    -2.7290736010148376e-10, -2.7174505759729094e-10, 
    -2.7064129229746025e-10, -2.6958300425640672e-10, 
    -2.6855735270452299e-10, -2.6755228835218409e-10, 
    -2.6655700546242002e-10, -2.655621775598767e-10, -2.6456009667269798e-10, 
    -2.6354465309251769e-10, -2.6251130540374373e-10, 
    -2.6145691353541164e-10, -2.6037966417189521e-10, -2.592789065030797e-10, 
    -2.5815508165102455e-10, -2.5700962922119935e-10, 
    -2.5584498160607065e-10, -2.5466453420178256e-10, 
    -2.5347267293167456e-10, -2.5227475367770576e-10, -2.510770969349743e-10, 
    -2.4988688503318021e-10, -2.4871201377907076e-10, 
    -2.4756081377029379e-10, -2.4644170558564607e-10, 
    -2.4536271301016473e-10, -2.4433094558234026e-10, 
    -2.4335200436641386e-10, -2.424294366123261e-10, -2.4156423721173888e-10, 
    -2.407545128933338e-10, -2.3999529531974183e-10, -2.3927862974713468e-10, 
    -2.3859386020225071e-10, -2.3792815881989487e-10, 
    -2.3726723890047075e-10, -2.3659623180224312e-10, 
    -2.3590057619319894e-10, -2.351669418190841e-10, -2.3438399879942665e-10, 
    -2.3354307219619852e-10, -2.3263853055036095e-10, 
    -2.3166798641584125e-10, -2.3063221926253121e-10, 
    -2.2953490761760415e-10, -2.2838218079684574e-10, 
    -2.2718206817281578e-10, -2.2594387835487186e-10, 
    -2.2467761109219209e-10, -2.2339340216280055e-10, 
    -2.2210106641587477e-10, -2.2080974277723067e-10, 
    -2.1952768421457649e-10, -2.1826211484952682e-10, 
    -2.1701919781833207e-10, -2.158040533655299e-10, -2.146208181542257e-10, 
    -2.1347269790847371e-10, -2.1236203614567598e-10, -2.1129033869648174e-10, 
    -2.1025830697327172e-10, -2.0926583892443041e-10, 
    -2.0831206517607899e-10, -2.0739538629219327e-10, 
    -2.0651357455098757e-10, -2.0566391876871941e-10, -2.048434564926166e-10, 
    -2.0404923384223096e-10, -2.0327864125180495e-10, 
    -2.0252974358409571e-10, -2.0180158670172486e-10, 
    -2.0109444523546345e-10, -2.0040998470425082e-10, 
    -1.9975126708332332e-10, -1.9912263371402256e-10, 
    -1.9852941670134357e-10, -1.979775365278643e-10, -1.9747297359486099e-10, 
    -1.9702120447786072e-10, -1.9662660639970886e-10, 
    -1.9629192281326269e-10, -1.9601780092813546e-10, 
    -1.9580246827541885e-10, -1.9564154612264652e-10, 
    -1.9552803552693941e-10, -1.9545243857928009e-10, 
    -1.9540304958565262e-10, -1.9536634153412287e-10, 
    -1.9532746258397838e-10, -1.9527079227214062e-10, 
    -1.9518055304737612e-10, -1.9504141810243201e-10, 
    -1.9483913279196868e-10, -1.9456108870865507e-10, 
    -1.9419685629483468e-10, -1.93738631740525e-10, -1.9318160873079902e-10, 
    -1.9252421338768021e-10, -1.9176824733510762e-10, -1.909188657124583e-10, 
    -1.8998445417180797e-10, -1.8897635688941628e-10, 
    -1.8790851226952832e-10, -1.8679697455731347e-10, -1.856593863576129e-10, 
    -1.8451438074436232e-10, -1.8338097757722827e-10, 
    -1.8227795237512749e-10, -1.8122323553001263e-10, 
    -1.8023332442794402e-10, -1.7932274401506346e-10, 
    -1.7850354738714471e-10, -1.7778491649766711e-10, 
    -1.7717282125246164e-10, -1.7666978861023565e-10, 
    -1.7627480289558444e-10, -1.7598332476037658e-10, 
    -1.7578744103010796e-10, -1.7567615437983037e-10, 
    -1.7563576091540414e-10, -1.7565034162362412e-10, 
    -1.7570227724105694e-10, -1.7577280856859283e-10, 
    -1.7584256545272247e-10, -1.7589208135663396e-10, 
    -1.7590224070340436e-10, -1.7585470975017963e-10, 
    -1.7573231007109946e-10, -1.7551939593958885e-10, 
    -1.7520222453965203e-10, -1.7476934868341561e-10, 
    -1.7421203285174374e-10, -1.7352466535320352e-10, 
    -1.7270515978479766e-10, -1.7175528639311908e-10, 
    -1.7068088039858268e-10, -1.6949191855963091e-10, 
    -1.6820236203050146e-10, -1.6682978565227591e-10, 
    -1.6539477908364992e-10, -1.6392014094036362e-10, 
    -1.6242990647676027e-10, -1.6094829183563112e-10, -1.594986123096503e-10, 
    -1.5810227353506676e-10, -1.5677790843891848e-10, 
    -1.5554071419407216e-10, -1.5440203487971783e-10, 
    -1.5336924035415899e-10, -1.5244583772455686e-10, 
    -1.5163182970840139e-10, -1.509242514136719e-10, -1.5031782967625506e-10, 
    -1.4980569342308387e-10, -1.4938005696111536e-10, 
    -1.4903283618567947e-10, -1.4875612605414382e-10, -1.485425212271276e-10, 
    -1.4838527570155549e-10, -1.4827828148461228e-10, 
    -1.4821591218096853e-10, -1.4819276203063302e-10, 
    -1.4820331737418778e-10, -1.482416196883868e-10, -1.4830096042459673e-10, 
    -1.4837365619703315e-10, -1.4845093983594782e-10, 
    -1.4852297831256536e-10, -1.485790215376935e-10, -1.4860768436526714e-10, 
    -1.4859733951510952e-10, -1.485365658867314e-10, -1.4841465174966305e-10, 
    -1.4822208193619895e-10, -1.4795097277948353e-10, -1.475954363259625e-10, 
    -1.4715185977816277e-10, -1.4661906492179708e-10, 
    -1.4599836502173559e-10, -1.4529353849462364e-10, 
    -1.4451073646729861e-10, -1.4365833446799008e-10, 
    -1.4274676249589114e-10, -1.4178830802893577e-10, 
    -1.4079691972181836e-10, -1.3978797688867651e-10, 
    -1.3877801563016057e-10, -1.3778439949258518e-10, 
    -1.3682489608829771e-10, -1.3591715464760736e-10, 
    -1.3507807405538067e-10, -1.3432307206849937e-10, 
    -1.3366529844607594e-10, -1.3311482947008778e-10, 
    -1.3267790561081888e-10, -1.3235630144141989e-10, 
    -1.3214689064794371e-10, -1.3204144689376352e-10, 
    -1.3202679762032661e-10, -1.3208526221872806e-10, 
    -1.3219542547997021e-10, -1.3233319685327305e-10, 
    -1.3247307591764629e-10, -1.325895347072218e-10, -1.3265843144973568e-10, 
    -1.3265832063461058e-10, -1.3257156240178481e-10, 
    -1.3238516236429118e-10, -1.3209126833818495e-10, 
    -1.3168730839584062e-10, -1.3117576783784214e-10, 
    -1.3056364621918382e-10, -1.2986167938303593e-10, -1.290833698208212e-10, 
    -1.2824395734394549e-10, -1.2735939368570304e-10, 
    -1.2644539895028301e-10, -1.2551667914226323e-10, 
    -1.2458632015321161e-10, -1.2366539061221396e-10, -1.22762737707891e-10, 
    -1.2188496193290958e-10, -1.2103654722729724e-10, 
    -1.2022009613570599e-10, -1.1943664467430906e-10, 
    -1.1868601315075524e-10, -1.1796719793814781e-10, 
    -1.1727874405170484e-10, -1.1661909572517237e-10, 
    -1.1598692365426757e-10, -1.1538138831421246e-10, 
    -1.1480233917727683e-10, -1.1425043355783454e-10, -1.137271582581617e-10, 
    -1.1323472575391834e-10, -1.1277589256882779e-10, 
    -1.1235363812698039e-10, -1.1197079861828911e-10, 
    -1.1162962179089716e-10, -1.1133133226214177e-10, 
    -1.1107573724092214e-10, -1.1086092076686189e-10, 
    -1.1068307227816899e-10, -1.1053648218912299e-10, 
    -1.1041372530364056e-10, -1.1030602227764999e-10, 
    -1.1020375050671003e-10, -1.1009707224192709e-10, 
    -1.0997661079236216e-10, -1.09834128238025e-10, -1.0966309893594364e-10, 
    -1.0945917070495818e-10, -1.0922043526390289e-10, 
    -1.0894748642815858e-10, -1.0864329273981031e-10, 
    -1.0831286943706364e-10, -1.079628252645889e-10, -1.0760081209160341e-10, 
    -1.0723496887335648e-10, -1.0687339055768461e-10, 
    -1.0652369582637512e-10, -1.061927026027343e-10, -1.0588624706824608e-10, 
    -1.0560911006945223e-10, -1.0536505192068175e-10, 
    -1.0515688622778463e-10, -1.0498657289327028e-10, 
    -1.0485527375111468e-10, -1.0476334355333331e-10, 
    -1.0471024352279077e-10, -1.0469439095538467e-10, 
    -1.0471295690239058e-10, -1.047616602572137e-10, -1.0483460180693804e-10, 
    -1.0492420515491483e-10, -1.0502128106834334e-10, 
    -1.0511526252265522e-10, -1.0519459781874184e-10, 
    -1.0524729757045626e-10, -1.052615774789652e-10, -1.0522655643140722e-10, 
    -1.0513290672614406e-10, -1.0497343203949608e-10, 
    -1.0474345474580593e-10, -1.0444102274340128e-10, 
    -1.0406686467431988e-10, -1.0362415855396226e-10, 
    -1.0311807594277495e-10, -1.0255523145519388e-10, 
    -1.0194304218669354e-10, -1.0128912119751456e-10, -1.00600728518063e-10, 
    -9.9884369907685969e-11, -9.9145552066727658e-11, 
    -9.8388700510734276e-11, -9.7617229466535479e-11, 
    -9.6833755213789281e-11, -9.6040339068503461e-11, 
    -9.5238797543709664e-11, -9.44309347950813e-11, -9.3618758440595765e-11, 
    -9.2804566450177091e-11, -9.199098189622547e-11, -9.1180879696980974e-11, 
    -9.037729746671748e-11, -8.958328022875178e-11, -8.8801813867228794e-11, 
    -8.8035721514250541e-11, -8.7287692441616467e-11, 
    -8.6560330504582506e-11, -8.5856285575784704e-11, 
    -8.5178391449975453e-11, -8.4529842042860264e-11, 
    -8.3914288826795487e-11, -8.3335919114468235e-11, 
    -8.2799405900787939e-11, -8.2309793982175455e-11, 
    -8.1872260902858472e-11, -8.1491817293326817e-11, 
    -8.1172934608308406e-11, -8.0919192700994626e-11, 
    -8.0732902595945681e-11, -8.0614836854265058e-11, 
    -8.0564004956734211e-11, -8.0577570550819506e-11, 
    -8.0650846191179493e-11, -8.0777433239254653e-11, 
    -8.0949411311754852e-11, -8.1157643446743767e-11, 
    -8.1392086590866232e-11, -8.1642141432876775e-11, 
    -8.1896991697053313e-11, -8.2145934839895866e-11, 
    -8.2378659308258638e-11, -8.2585540285681397e-11, 
    -8.2757855010142077e-11, -8.2888020020270725e-11, 
    -8.2969777275190161e-11, -8.2998403380163162e-11, 
    -8.2970874516959435e-11, -8.2886035419174838e-11, 
    -8.2744714188520611e-11, -8.254980536842658e-11, -8.2306245409631583e-11, 
    -8.2020937219724357e-11, -8.1702515972164989e-11, 
    -8.1361028809156363e-11, -8.1007456929212273e-11, 
    -8.0653175165898896e-11, -8.0309284968865774e-11, 
    -7.9985951771478485e-11, -7.9691725669203894e-11, 
    -7.9432947733568278e-11, -7.9213248482175086e-11, 
    -7.9033263440137221e-11, -7.8890488205183e-11, -7.8779416940045049e-11, 
    -7.8691866394400265e-11, -7.8617526229101851e-11, 
    -7.8544670091600626e-11, -7.8461016720073995e-11, 
    -7.8354621296746035e-11, -7.8214775577333543e-11, 
    -7.8032810917287588e-11, -7.7802794570892506e-11, 
    -7.7521979357002654e-11, -7.7191050799437472e-11, 
    -7.6814080187870948e-11, -7.6398246106768891e-11, 
    -7.5953269852968563e-11, -7.5490687052156651e-11, 
    -7.5022932138192802e-11, -7.4562398940927421e-11, 
    -7.4120468056109881e-11, -7.3706650723284997e-11, 
    -7.3327878141555945e-11, -7.2988051545319508e-11, 
    -7.2687809620413834e-11, -7.2424621340030032e-11, 
    -7.2193110569615773e-11, -7.1985649681056912e-11, 
    -7.1793096808363994e-11, -7.1605683560516538e-11, 
    -7.1413891040825699e-11, -7.1209318812392083e-11, 
    -7.0985396183612069e-11, -7.0737978854825714e-11, 
    -7.0465669626474689e-11, -7.0169966896862096e-11, 
    -6.9855125783840292e-11, -6.952786786320705e-11, -6.9196854732265228e-11, 
    -6.8872077874212248e-11, -6.8564129916538277e-11, 
    -6.8283485827177418e-11, -6.8039801456879951e-11, 
    -6.7841300913974589e-11, -6.7694269708049922e-11, 
    -6.7602734214576447e-11, -6.756826754982307e-11, -6.7589995773055212e-11, 
    -6.7664725641345682e-11, -6.7787244658008947e-11, 
    -6.7950672355135917e-11, -6.8146920813991694e-11, 
    -6.8367151128095337e-11, -6.8602249477922999e-11, 
    -6.8843241706786705e-11, -6.9081701737776207e-11, 
    -6.9310051049958492e-11, -6.9521835931847771e-11, 
    -6.9711891760721262e-11, -6.9876493686571392e-11, 
    -7.0013421580708762e-11, -7.0121970344532356e-11, 
    -7.0202901427570306e-11, -7.0258376064889583e-11, 
    -7.0291783202876268e-11, -7.0307552444137656e-11, 
    -7.0310872861306983e-11, -7.0307423662714675e-11, 
    -7.0302996952814888e-11, -7.0303179064592594e-11, 
    -7.0312978208247657e-11, -7.0336519358245978e-11, 
    -7.0376768921130612e-11, -7.0435370201838216e-11, 
    -7.0512530927789541e-11, -7.0607051968102992e-11, 
    -7.0716419964321261e-11, -7.0837025515905458e-11, -7.096440370678509e-11, 
    -7.1093576821641636e-11, -7.1219347466752124e-11, 
    -7.1336639876225445e-11, -7.1440742458741937e-11, 
    -7.1527544815610205e-11, -7.1593657230464428e-11, 
    -7.1636493490803438e-11, -7.1654249958348733e-11, 
    -7.1645875416966983e-11, -7.1610954260994282e-11, 
    -7.1549629570170452e-11, -7.1462485896067243e-11, -7.135048251662882e-11, 
    -7.1214895748222844e-11, -7.1057321564545879e-11, 
    -7.0879671777608288e-11, -7.0684217615211865e-11, 
    -7.0473602917267976e-11, -7.0250868372443267e-11, 
    -7.0019405473814347e-11, -6.9782904269469322e-11, 
    -6.9545217274234342e-11, -6.931020304217061e-11, -6.9081503178425201e-11, 
    -6.8862350306928101e-11, -6.8655323959016058e-11, 
    -6.8462186136542132e-11, -6.8283714417080796e-11, 
    -6.8119649411403516e-11, -6.7968678326404189e-11, 
    -6.7828507824234632e-11, -6.7695994102040132e-11, 
    -6.7567353997117718e-11, -6.7438376858382791e-11, -6.730469118397681e-11, 
    -6.7162002939371102e-11, -6.7006331582048913e-11, 
    -6.6834178168146107e-11, -6.6642687965578949e-11, 
    -6.6429710566628915e-11, -6.619382503558682e-11, -6.5934289352157902e-11, 
    -6.5650956351904757e-11, -6.5344123351666815e-11, 
    -6.5014397754417646e-11, -6.4662511331971744e-11, 
    -6.4289194787982997e-11, -6.3895045501220305e-11, 
    -6.3480479243544702e-11, -6.304568644865613e-11, -6.2590709118290204e-11, 
    -6.2115515648501926e-11, -6.162013354902722e-11, -6.1104792450290179e-11, 
    -6.0570089014077409e-11, -6.0017102136262765e-11, 
    -5.9447482612439452e-11, -5.8863474930596923e-11, 
    -5.8267915516075181e-11, -5.7664121655773931e-11, 
    -5.7055795895230213e-11, -5.6446867370472848e-11, 
    -5.5841335625207554e-11, -5.5243120540962976e-11, 
    -5.4655983029140206e-11, -5.4083448788558647e-11, 
    -5.3528812887358604e-11, -5.299517102033457e-11, -5.2485522979452638e-11, 
    -5.2002871692569871e-11, -5.155033614107467e-11, -5.1131238472753074e-11, 
    -5.0749177044133003e-11, -5.0408016370567688e-11, 
    -5.0111840332567886e-11, -4.9864815561009062e-11, 
    -4.9671021271057163e-11, -4.9534194700083323e-11, 
    -4.9457463182749839e-11, -4.9443035996136414e-11, 
    -4.9491901778387562e-11, -4.9603532942164268e-11, 
    -4.9775662330133506e-11, -5.0004082177587799e-11, 
    -5.0282577635136391e-11, -5.0602928870694289e-11, 
    -5.0955065150605904e-11, -5.1327334698587513e-11, 
    -5.1706914102454284e-11, -5.2080317847153397e-11, 
    -5.2434030720331819e-11, -5.2755158426644176e-11, 
    -5.3032103328594929e-11, -5.3255161541165762e-11, 
    -5.3417064077396853e-11, -5.3513306040737889e-11, -5.354232811697984e-11, 
    -5.3505454129087174e-11, -5.3406660278532163e-11, 
    -5.3252128072539097e-11, -5.3049691155216141e-11, 
    -5.2808175823934022e-11, -5.2536772144612488e-11, 
    -5.2244420401682884e-11, -5.1939341713210942e-11, 
    -5.1628688397158278e-11, -5.1318398459534098e-11, 
    -5.1013168195698002e-11, -5.0716602109726029e-11, -5.043141137523411e-11, 
    -5.0159697157074339e-11, -4.9903182377675454e-11, 
    -4.9663429182004713e-11, -4.9441940099622009e-11, 
    -4.9240199945399503e-11, -4.9059596308323433e-11, 
    -4.8901316205245111e-11, -4.8766180335256039e-11, 
    -4.8654507925096546e-11, -4.8565999959997253e-11, 
    -4.8499714390057926e-11, -4.8454087369565549e-11, 
    -4.8427058537956125e-11, -4.8416223599965482e-11, 
    -4.8419040738010776e-11, -4.8432998400287439e-11, 
    -4.8455805592531246e-11, -4.8485480768284533e-11, 
    -4.8520396699577276e-11, -4.8559258438170957e-11, 
    -4.8601036198767219e-11, -4.8644851572970137e-11, 
    -4.8689887948660656e-11, -4.8735285594071736e-11, 
    -4.8780116780609447e-11, -4.8823370373431824e-11, -4.886402862780437e-11, 
    -4.890114343728562e-11, -4.8933968683404314e-11, -4.8962052618705223e-11, 
    -4.8985340281778321e-11, -4.9004180386025011e-11, 
    -4.9019317717675692e-11, -4.9031769753172412e-11, 
    -4.9042672052746785e-11, -4.9053054900137607e-11, 
    -4.9063600747935282e-11, -4.9074398782680348e-11, -4.908473804329214e-11, 
    -4.9092948097217359e-11, -4.909632386305143e-11, -4.9091135663817409e-11, 
    -4.907275040711658e-11, -4.90358261307206e-11, -4.8974589637152029e-11, 
    -4.8883153157712693e-11, -4.8755868720607639e-11, -4.858765145746114e-11, 
    -4.837427497672484e-11, -4.8112602606000038e-11, -4.7800732850010786e-11, 
    -4.7438079393707885e-11, -4.7025348934256578e-11, 
    -4.6564467789225765e-11, -4.6058470189231171e-11, 
    -4.5511345333409816e-11, -4.4927896741427374e-11, 
    -4.4313614234116281e-11, -4.3674570075108301e-11, 
    -4.3017356537345692e-11, -4.2349035801506115e-11, 
    -4.1677105441713401e-11, -4.1009471309576675e-11, -4.035439495470395e-11, 
    -3.9720384798677625e-11, -3.9116060497541969e-11, 
    -3.8549952647245277e-11, -3.8030244266759055e-11, 
    -3.7564482676339329e-11, -3.7159266190520821e-11, 
    -3.6819925854389424e-11, -3.6550243461924955e-11, 
    -3.6352230020224725e-11, -3.6225965940793551e-11, 
    -3.6169544563534006e-11, -3.6179110843920811e-11, 
    -3.6248988392617357e-11, -3.6371897835289686e-11, 
    -3.6539241040168426e-11, -3.6741417538224696e-11, 
    -3.6968178085567063e-11, -3.7208957215766229e-11, 
    -3.7453192399175726e-11, -3.7690604341565287e-11, 
    -3.7911449797593626e-11, -3.8106720444888215e-11, 
    -3.8268339506610823e-11, -3.838931499025489e-11, -3.8463913027642062e-11, 
    -3.8487803626425221e-11, -3.8458242736486568e-11, 
    -3.8374225537985347e-11, -3.8236625707490187e-11, 
    -3.8048283977025813e-11, -3.7814059104232105e-11, 
    -3.7540746466582041e-11, -3.7236903051212155e-11, 
    -3.6912548493989169e-11, -3.6578726148720643e-11, 
    -3.6246984932035269e-11, -3.5928772727881303e-11, 
    -3.5634817172558825e-11, -3.5374544712015877e-11, 
    -3.5155575748034578e-11, -3.4983373827015022e-11, 
    -3.4861050355838354e-11, -3.478938394099732e-11, -3.4767007305132715e-11, 
    -3.4790767697472153e-11, -3.4856189388478014e-11, 
    -3.4958025727310068e-11, -3.5090786676169622e-11, 
    -3.5249214834506279e-11, -3.5428683649765373e-11, 
    -3.5625417277869473e-11, -3.5836597456495708e-11, 
    -3.6060342830276976e-11, -3.6295542436931267e-11, 
    -3.6541643911269179e-11, -3.6798390078567249e-11, 
    -3.7065568969655515e-11, -3.7342801063248283e-11, 
    -3.7629389228124367e-11, -3.7924233872587598e-11, 
    -3.8225821901555864e-11, -3.8532259831705258e-11, 
    -3.8841329099331916e-11, -3.9150556060943313e-11, 
    -3.9457253025095616e-11, -3.9758533030549919e-11, 
    -4.0051296332225782e-11, -4.0332171001833327e-11, 
    -4.0597462708798985e-11, -4.0843106681394431e-11, 
    -4.1064646713920334e-11, -4.125726799794701e-11, -4.1415923835516586e-11, 
    -4.153550709984093e-11, -4.1611095177167351e-11, -4.1638251865978482e-11, 
    -4.1613333229038056e-11, -4.1533780228151931e-11, 
    -4.1398390124865481e-11, -4.1207480256658723e-11, 
    -4.0962973369237163e-11, -4.0668373577368259e-11, 
    -4.0328626268158125e-11, -3.9949886471740858e-11, 
    -3.9539215399865466e-11, -3.9104216017598852e-11, 
    -3.8652659795710966e-11, -3.8192105506767801e-11, 
    -3.7729598413318257e-11, -3.7271398809807723e-11, 
    -3.6822813794065701e-11, -3.6388127564225946e-11, 
    -3.5970627649713219e-11, -3.5572735363017926e-11, 
    -3.5196200420249946e-11, -3.4842365008878363e-11, 
    -3.4512462279259611e-11, -3.4207894890668886e-11, 
    -3.3930488392447709e-11, -3.3682673194379339e-11, 
    -3.3467566911170709e-11, -3.3288947858705333e-11, 
    -3.3151112039996831e-11, -3.3058633222788838e-11, 
    -3.3016025593247136e-11, -3.3027371839034591e-11, 
    -3.3095947377120166e-11, -3.3223868220214374e-11, 
    -3.3411840575872499e-11, -3.3659006143764428e-11, 
    -3.3962921071680982e-11, -3.4319660672843608e-11, 
    -3.4724055270960476e-11, -3.5169983041781529e-11, 
    -3.5650733956071609e-11, -3.6159339279990757e-11, 
    -3.6688876582454119e-11, -3.7232681209331916e-11, -3.778444315169831e-11, 
    -3.8338194166770906e-11, -3.8888212725965464e-11, 
    -3.9428835883954696e-11, -3.995425328806225e-11, -4.0458306028755835e-11, 
    -4.0934367232956267e-11, -4.1375292415937767e-11, 
    -4.1773518517598798e-11, -4.212127687278187e-11, -4.2410926603104826e-11, 
    -4.2635379297102444e-11, -4.2788579295491574e-11, 
    -4.2865960376569609e-11, -4.2864874987538548e-11, 
    -4.2784887775336438e-11, -4.2627940356843964e-11, 
    -4.2398340534840012e-11, -4.210257743853871e-11, -4.1748963889649926e-11, 
    -4.1347163432328043e-11, -4.0907607288917417e-11, 
    -4.0440902556867335e-11, -3.9957231295043325e-11, 
    -3.9465862715548579e-11, -3.8974756571163251e-11, 
    -3.8490334682286112e-11, -3.8017410164300791e-11, 
    -3.7559288912129638e-11, -3.7117987052848955e-11, 
    -3.6694581172818173e-11, -3.628958870658407e-11, -3.5903358959834979e-11, 
    -3.553640538927921e-11, -3.5189669357187497e-11, -3.4864620970349099e-11, 
    -3.4563244003107343e-11, -3.4287851636953363e-11, 
    -3.4040790926063214e-11, -3.3824039916678619e-11, 
    -3.3638768961815036e-11, -3.3484898452285564e-11, -3.336073783826104e-11, 
    -3.3262749361859103e-11, -3.3185458331658079e-11, 
    -3.3121565492092173e-11, -3.3062286292280381e-11, 
    -3.2997834972206667e-11, -3.2918085918147087e-11, 
    -3.2813313682838307e-11, -3.2674968981923733e-11, 
    -3.2496397458716872e-11, -3.227344465002166e-11, -3.200486966129332e-11, 
    -3.1692545723453829e-11, -3.1341407409637168e-11, 
    -3.0959156875049664e-11, -3.0555764601359601e-11, 
    -3.0142788755254414e-11, -2.9732609898250818e-11, 
    -2.9337613610032426e-11, -2.8969413930772827e-11, -2.863817338144029e-11, 
    -2.8352053246989507e-11, -2.8116845031358569e-11, 
    -2.7935772959111776e-11, -2.7809482210502338e-11, 
    -2.7736175687523058e-11, -2.7711888130670899e-11, 
    -2.7730843953853171e-11, -2.7785875887700334e-11, 
    -2.7868857477742392e-11, -2.7971147003274021e-11, 
    -2.8083985624979919e-11, -2.819885678391988e-11, -2.8307796232538372e-11, 
    -2.8403662084418752e-11, -2.8480333455174866e-11, -2.85328921303079e-11, 
    -2.8557741161493813e-11, -2.8552711937837215e-11, 
    -2.8517121216369724e-11, -2.8451809619562709e-11, 
    -2.8359137223830972e-11, -2.8242939668862012e-11, 
    -2.8108439624200656e-11, -2.7962099368456407e-11, 
    -2.7811415355294159e-11, -2.7664661915141687e-11, 
    -2.7530562071460284e-11, -2.7417924933024674e-11, 
    -2.7335231161838129e-11, -2.7290226734965534e-11, 
    -2.7289509449781094e-11, -2.733815069708186e-11, -2.7439370632167083e-11, 
    -2.7594339056023055e-11, -2.7802031980757782e-11, 
    -2.8059247388174988e-11, -2.8360722905581737e-11, 
    -2.8699395406350658e-11, -2.9066756775535104e-11, 
    -2.9453313977454591e-11, -2.9849096605738851e-11, 
    -3.0244212836857015e-11, -3.0629375082171188e-11, 
    -3.0996419410775169e-11, -3.1338722919859768e-11, 
    -3.1651538077785012e-11, -3.1932208940215678e-11, 
    -3.2180244296301276e-11, -3.2397262600729815e-11, 
    -3.2586817129124702e-11, -3.275408968504236e-11, -3.2905505749954438e-11, 
    -3.3048269262743175e-11, -3.3189884957311453e-11, 
    -3.3337638693184092e-11, -3.3498144036494099e-11, -3.367691563006069e-11, 
    -3.3878009398801924e-11, -3.4103751229701365e-11, 
    -3.4354580358921956e-11, -3.4628955928985665e-11, 
    -3.4923376426327923e-11, -3.5232472868632167e-11, 
    -3.5549200856342613e-11, -3.5865081032940838e-11, -3.617051572452228e-11, 
    -3.6455162227536456e-11, -3.6708330362413121e-11, 
    -3.6919426079886588e-11, -3.7078413680925145e-11, 
    -3.7176260662866626e-11, -3.7205381442751934e-11, 
    -3.7160030878456733e-11, -3.7036625554521267e-11, 
    -3.6833976451862097e-11, -3.655343929387413e-11, -3.6198908464985007e-11, 
    -3.5776711694030189e-11, -3.5295369391173672e-11, 
    -3.4765250932574846e-11, -3.4198138923458038e-11, 
    -3.3606735215474924e-11, -3.3004141928838449e-11, 
    -3.2403345049225704e-11, -3.1816737747648421e-11, 
    -3.1255719042979013e-11, -3.0730345096968418e-11, 
    -3.0249120949417572e-11, -2.9818840290426844e-11, 
    -2.9444518731639922e-11, -2.9129401087205087e-11, 
    -2.8874997632248055e-11, -2.8681155851230064e-11, 
    -2.8546131368525581e-11, -2.8466660441901701e-11, -2.843802551432001e-11, 
    -2.8454114903872216e-11, -2.8507516572868768e-11, 
    -2.8589632413183714e-11, -2.8690852416743296e-11, 
    -2.8800800948008209e-11, -2.8908680373379374e-11, 
    -2.9003682709769862e-11, -2.9075488135830489e-11, 
    -2.9114808295887177e-11, -2.9113929647817822e-11, 
    -2.9067228792830301e-11, -2.8971609569717166e-11, -2.882679924346139e-11, 
    -2.8635471228435391e-11, -2.8403183906795999e-11, 
    -2.8138107447164293e-11, -2.7850566757508152e-11, 
    -2.7552408834321199e-11, -2.7256271785306963e-11, 
    -2.6974778137861191e-11, -2.6719744417325663e-11, 
    -2.6501448107103838e-11, -2.6328025386853362e-11, 
    -2.6205027607823686e-11, -2.6135178079201017e-11, 
    -2.6118335902364436e-11, -2.615165698713892e-11, -2.6229932000111782e-11, 
    -2.6346067649918291e-11, -2.6491673330232104e-11, 
    -2.6657681510540831e-11, -2.6834976947062421e-11, 
    -2.7014980282991475e-11, -2.7190134451915395e-11, 
    -2.7354283558557698e-11, -2.7502907672977205e-11, 
    -2.7633229499936235e-11, -2.7744159510503245e-11, 
    -2.7836138239903349e-11, -2.7910872087269477e-11, 
    -2.7970995024295151e-11, -2.80197050169064e-11, -2.806037728096721e-11, 
    -2.8096213721520907e-11, -2.8129934508563625e-11, 
    -2.8163530559124513e-11, -2.8198094131893611e-11, 
    -2.8233724890871171e-11, -2.8269510341054242e-11, 
    -2.8303588977992142e-11, -2.8333278700159306e-11, 
    -2.8355245100957039e-11, -2.836574489825738e-11, -2.8360899505144519e-11, 
    -2.8337010944140134e-11, -2.8290881203046482e-11, 
    -2.8220138263069752e-11, -2.8123576002763357e-11, 
    -2.8001431010999301e-11, -2.7855605572294662e-11, 
    -2.7689832403194158e-11, -2.7509718304250651e-11, 
    -2.7322688286026089e-11, -2.7137811505169306e-11, 
    -2.6965484995319123e-11, -2.6817033578136299e-11, 
    -2.6704198611470316e-11, -2.6638544870404729e-11, 
    -2.6630834472692118e-11, -2.6690409605542247e-11, 
    -2.6824581662106952e-11, -2.7038100248834494e-11, 
    -2.7332722177872384e-11, -2.7706918353633886e-11, 
    -2.8155727476779074e-11, -2.8670791470776211e-11, 
    -2.9240553993430613e-11, -2.9850638460486864e-11, 
    -3.0484362918862784e-11, -3.1123395787104358e-11, 
    -3.1748486190599892e-11, -3.2340243824150488e-11, 
    -3.2879929074786968e-11, -3.3350214891587733e-11, 
    -3.3735873069485983e-11, -3.4024359795171565e-11, 
    -3.4206290551506241e-11, -3.427576397005267e-11, -3.4230552844336981e-11, 
    -3.4072130734039223e-11, -3.3805562499362513e-11, 
    -3.3439242572029539e-11, -3.2984503248485515e-11, 
    -3.2455108940812627e-11, -3.1866653263944831e-11, 
    -3.1235867857837289e-11, -3.0579922776361472e-11, 
    -2.9915692013679622e-11, -2.9259066368880459e-11, 
    -2.8624360304132895e-11, -2.8023800035279253e-11, 
    -2.7467165981058678e-11, -2.6961592240278669e-11, 
    -2.6511516697177728e-11, -2.6118785245176594e-11, 
    -2.5782885798962294e-11, -2.550126948810233e-11, -2.5269737563904776e-11, 
    -2.5082854540292842e-11, -2.4934336351631794e-11, 
    -2.4817420618997452e-11, -2.4725188437917206e-11, 
    -2.4650840706993099e-11, -2.4587929112061039e-11, 
    -2.4530573563256346e-11, -2.447365480487287e-11, -2.4413012814774987e-11, 
    -2.4345644970421642e-11, -2.4269896956339707e-11, -2.418563315509786e-11, 
    -2.4094370916696977e-11, -2.3999322261536164e-11, -2.390535793033819e-11, 
    -2.3818831803331724e-11, -2.3747287418585941e-11, 
    -2.3699023868067495e-11, -2.368256216693632e-11, -2.3706026077368214e-11, 
    -2.3776497114360287e-11, -2.3899398418734996e-11, 
    -2.4077959965665834e-11, -2.4312817405230837e-11, 
    -2.4601783478870078e-11, -2.4939843357189584e-11, 
    -2.5319353029958147e-11, -2.5730435969709112e-11, 
    -2.6161561235532955e-11, -2.6600251641179691e-11, 
    -2.7033853578060806e-11, -2.7450312424351611e-11, 
    -2.7838897509174591e-11, -2.8190800282716774e-11, 
    -2.8499575093974053e-11, -2.8761389695903682e-11, 
    -2.8975059017822867e-11, -2.914187970484769e-11, -2.9265283501974946e-11, 
    -2.9350332593101093e-11, -2.9403118562216019e-11, 
    -2.9430117086899626e-11, -2.9437541992549126e-11, 
    -2.9430767465839246e-11, -2.9413858444512821e-11, 
    -2.9389247902223109e-11, -2.9357590459724134e-11, 
    -2.9317791025385824e-11, -2.9267213257598324e-11, 
    -2.9202038288763737e-11, -2.911774899047893e-11, -2.9009672277649428e-11, 
    -2.8873561583451752e-11, -2.8706146293867453e-11, 
    -2.8505593974846736e-11, -2.8271873404999591e-11, 
    -2.8006976103393717e-11, -2.771495652650947e-11, -2.740184166141955e-11, 
    -2.7075387640357213e-11, -2.6744714425014142e-11, -2.64198484383266e-11, 
    -2.6111228255781696e-11, -2.5829174722844659e-11, -2.558338969102593e-11, 
    -2.5382489855477827e-11, -2.5233612254447575e-11, 
    -2.5142086650750095e-11, -2.5111208370571554e-11,
  // Sqw-F(4, 0-1999)
    0.041175817675317861, 0.041148391701459106, 0.041066465015250728, 
    0.040931070011790936, 0.040743858465159863, 0.040507005485607123, 
    0.040223088762058767, 0.039894954885272997, 0.039525585463922742, 
    0.039117975256691043, 0.038675032742294412, 0.038199510682650678, 
    0.037693970664936301, 0.037160781765890313, 0.036602149808201034, 
    0.036020170574308612, 0.035416898120844253, 0.034794418192264004, 
    0.034154916726646251, 0.033500734510150128, 0.032834400985021876, 
    0.032158642779934909, 0.031476365393229767, 0.030790609293049373, 
    0.030104484206117721, 0.029421087312207734, 0.028743412290216541, 
    0.0280742566141103, 0.027416134205694061, 0.026771199629874603, 
    0.026141188639746096, 0.025527378247922904, 0.024930567823133104, 
    0.024351081166922629, 0.023788788246072542, 0.023243144313141208, 
    0.022713243549367507, 0.022197884066979662, 0.021695641032190818, 
    0.021204944723242143, 0.020724160436620665, 0.020251667243617981, 
    0.019785932661353287, 0.019325580358681371, 0.018869448119569799, 
    0.018416633500420772, 0.017966525004533298, 0.017518817194590877, 
    0.017073508974675071, 0.016630885256907237, 0.01619148330564045, 
    0.015756046117416406, 0.015325466129370233, 0.01490072324131396, 
    0.014482821500966411, 0.014072728789422942, 0.013671323451862769, 
    0.013279351088892962, 0.012897393737856788, 0.012525852539114708, 
    0.012164943820375824, 0.011814707460196649, 0.011475025510159392, 
    0.011145648436377078, 0.010826226022720042, 0.010516339962341383, 
    0.010215535419573285, 0.0099233493139890706, 0.0096393336889040344, 
    0.0093630731985782038, 0.0090941964069317302, 0.0088323811732827495, 
    0.0085773548629180536, 0.0083288904377699351, 0.0080867996498115227, 
    0.0078509245876832671, 0.0076211287375123043, 0.0073972885402476454, 
    0.0071792861904970097, 0.0069670041550758954, 0.0067603216195783189, 
    0.0065591128209247672, 0.0063632470119869295, 0.0061725896462631264, 
    0.0059870042773110853, 0.0058063546453996692, 0.0056305064725625676, 
    0.0054593285995656327, 0.0052926932590934683, 0.0051304754665622114, 
    0.0049725516963455294, 0.0048187981684731981, 0.0046690891735890819, 
    0.004523295894033527, 0.0043812861290660528, 0.0042429252078828176, 
    0.0041080781929955512, 0.0039766132663581226, 0.0038484059844498294, 
    0.0037233439194945331, 0.0036013310997923226, 0.0034822916404498106, 
    0.0033661720214795497, 0.0032529416147523927, 0.0031425912642764672, 
    0.0030351299570709569, 0.0029305798521278331, 0.0028289701315223651, 
    0.0027303302752969883, 0.0026346834240408993, 0.0025420404746721737, 
    0.0024523954612603112, 0.0023657226186797552, 0.0022819753341426223, 
    0.0022010869853710687, 0.0021229734694944943, 0.0020475370656764086, 
    0.0019746711633272089, 0.0019042653356682456, 0.0018362102467776443, 
    0.0017704019431935378, 0.0017067451868593847, 0.0016451556188310402, 
    0.0015855606851568696, 0.0015278993906718448, 0.0014721210587018349, 
    0.0014181833545657242, 0.0013660498730058335, 0.0013156875941031268, 
    0.0012670644832476195, 0.0012201474561763998, 0.0011749008597981372, 
    0.0011312855437578526, 0.0010892585257674683, 0.0010487731929193188, 
    0.0010097799361923803, 0.00097222708811075338, 0.00093606202357903812, 
    0.00090123228904769709, 0.00086768664203060511, 0.00083537590789656215, 
    0.00080425359024650174, 0.00077427620201361283, 0.00074540331424535484, 
    0.0007175973464561867, 0.00069082314502285952, 0.00066504741316222957, 
    0.00064023806665330972, 0.00061636359296055238, 0.0005933924874865767, 
    0.00057129282955735027, 0.00055003204332562314, 0.00052957686669207436, 
    0.00050989352687381495, 0.00049094809712252753, 0.00047270698816347475, 
    0.00045513751276877594, 0.00043820845441477327, 0.00042189057214642281, 
    0.00040615698338006446, 0.0003909833830625331, 0.00037634807905049378, 
    0.00036223184681669681, 0.00034861762847417349, 0.00033549011873280432, 
    0.00032283529155153199, 0.00031063992468991451, 0.00029889117500685072, 
    0.00028757624622026493, 0.00027668217487414055, 0.00026619574199134987, 
    0.00025610350005580312, 0.00024639189007260806, 0.00023704741343578801, 
    0.00022805681928556753, 0.00021940727011895037, 0.00021108645586948542, 
    0.00020308263800648712, 0.0001953846184604155, 0.00018798164126526204, 
    0.00018086324579933731, 0.00017401909793660089, 0.00016743882844666558, 
    0.00016111190646415723, 0.00015502757030117149, 0.00014917482935014855, 
    0.00014354254069374802, 0.00013811955379562866, 0.00013289490766972499, 
    0.00012785805831835216, 0.00012299911068393887, 0.00011830902912272452, 
    0.00011377980328398678, 0.00010940455170846166, 0.00010517755262275387, 
    0.00010109419935723018, 9.7150885597278904e-05, 9.334483244919449e-05, 
    8.9673874404041476e-05, 8.6136224304098763e-05, 8.2730238199766432e-05, 
    7.9454199625317906e-05, 7.6306139623247613e-05, 7.3283704279224535e-05, 
    7.038407615830153e-05, 6.7603950466204557e-05, 6.4939561574370511e-05, 
    6.2386751246797215e-05, 5.9941066862256726e-05, 5.7597876357954904e-05, 
    5.5352486574238293e-05, 5.32002530359178e-05, 5.1136671693012767e-05, 
    4.9157446387707563e-05, 4.7258529374309356e-05, 4.5436135655128511e-05, 
    4.3686734811670409e-05, 4.200702611127624e-05, 4.0393903780557769e-05, 
    3.8844419429241599e-05, 3.735574778120112e-05, 3.592516033876005e-05, 
    3.4550009655024379e-05, 3.3227724834107956e-05, 3.1955817015950508e-05, 
    3.0731892174079441e-05, 2.9553667714796895e-05, 2.8418989171908992e-05, 
    2.7325843696259642e-05, 2.6272367917721308e-05, 2.5256848920718796e-05, 
    2.4277718313741704e-05, 2.3333540484535212e-05, 2.2422996955168803e-05, 
    2.1544869180285362e-05, 2.0698022138718295e-05, 1.988139068947261e-05, 
    1.9093969995325237e-05, 1.8334810491332144e-05, 1.7603017039079505e-05, 
    1.6897751192336393e-05, 1.6218235011756234e-05, 1.5563754662664374e-05, 
    1.4933662123254517e-05, 1.4327373683236708e-05, 1.3744364455194911e-05, 
    1.3184158756365323e-05, 1.2646316848729226e-05, 1.2130419056414089e-05, 
    1.1636048643512532e-05, 1.116277499002971e-05, 1.071013854375687e-05, 
    1.0277638773843858e-05, 9.8647259597229854e-06, 9.47079718100166e-06, 
    9.0951964039187042e-06, 8.7372181521812216e-06, 8.3961139580139921e-06, 
    8.0711006410543056e-06, 7.7613694661861752e-06, 7.4660953667365755e-06, 
    7.1844456524672956e-06, 6.9155879015655541e-06, 6.6586970133454263e-06, 
    6.4129616238631762e-06, 6.1775902278400705e-06, 5.95181738623033e-06, 
    5.7349103312249358e-06, 5.5261761246244267e-06, 5.3249693134449267e-06, 
    5.1306997950556027e-06, 4.9428403956819738e-06, 4.7609335149455351e-06, 
    4.5845961246869361e-06, 4.4135224443801084e-06, 4.2474837499948747e-06, 
    4.0863249910157344e-06, 3.9299581670976909e-06, 3.7783527144452284e-06, 
    3.6315234365374379e-06, 3.4895167462762037e-06, 3.3523961402907215e-06, 
    3.2202278813319098e-06, 3.0930678189809446e-06, 2.9709501396852654e-06, 
    2.8538786276535037e-06, 2.7418207659096926e-06, 2.6347047471674181e-06, 
    2.5324192267905767e-06, 2.4348154625691908e-06, 2.3417113624309249e-06, 
    2.2528969083881603e-06, 2.1681404350399675e-06, 2.0871953014995516e-06, 
    2.009806584795053e-06, 1.9357175219644197e-06, 1.8646755170443381e-06, 
    1.7964375970654102e-06, 1.7307752405573508e-06, 1.6674785162051219e-06, 
    1.6063594633051339e-06, 1.5472546325585663e-06, 1.4900266950537287e-06, 
    1.4345650311570214e-06, 1.3807852344448475e-06, 1.3286275121150651e-06, 
    1.2780540281742813e-06, 1.2290453133500975e-06, 1.181595944399225e-06, 
    1.1357097658334029e-06, 1.0913949763039538e-06, 1.0486594240354513e-06, 
    1.007506443749137e-06, 9.6793152319857351e-07, 9.2992001278004116e-07, 
    8.9344599641242265e-07, 8.5847233448993649e-07, 8.2495178432080594e-07, 
    7.9282900952796902e-07, 7.620432193202181e-07, 7.3253113628586118e-07, 
    7.0422998230983839e-07, 6.7708019355060909e-07, 6.51027624271982e-07, 
    6.2602506668060357e-07, 6.0203299244241711e-07, 5.7901950054304467e-07, 
    5.5695952924848259e-07, 5.3583344937206581e-07, 5.1562520020081819e-07, 
    4.9632015496046566e-07, 4.7790291289286144e-07, 4.6035520946113714e-07, 
    4.4365411992606789e-07, 4.2777070467301123e-07, 4.1266921119566466e-07, 
    3.9830690704590397e-07, 3.8463457327862904e-07, 3.7159763864159964e-07, 
    3.5913788495383705e-07, 3.4719560501660765e-07, 3.3571205219443388e-07, 
    3.2463198787461586e-07, 3.139061161050823e-07, 3.0349319520294478e-07, 
    2.9336163744600582e-07, 2.8349044789215311e-07, 2.7386941025696791e-07, 
    2.6449849450739953e-07, 2.5538653211544009e-07, 2.465492712798275e-07, 
    2.3800698026780003e-07, 2.2978180465327616e-07, 2.2189510160376512e-07, 
    2.143649683778405e-07, 2.0720415621375405e-07, 2.0041851662776969e-07, 
    1.9400607246022063e-07, 1.8795674530389085e-07, 1.8225271304107618e-07, 
    1.768693200670692e-07, 1.7177642478317838e-07, 1.6694004496997275e-07, 
    1.623241538864786e-07, 1.5789248535288037e-07, 1.5361022336370107e-07, 
    1.4944547569165757e-07, 1.4537045897563254e-07, 1.4136235028653864e-07, 
    1.3740378597453803e-07, 1.3348301017627612e-07, 1.2959369384640073e-07, 
    1.2573445980310879e-07, 1.2190816217895489e-07, 1.1812097901042366e-07, 
    1.1438138594519776e-07, 1.106990849738993e-07, 1.0708396494155474e-07, 
    1.0354516748762864e-07, 1.0009032335132681e-07, 9.6725007920730319e-08, 
    9.3452443926016626e-08, 9.0273453787879004e-08, 8.7186639064209186e-08, 
    8.4188741570960148e-08, 8.1275125050041907e-08, 7.8440308447007369e-08, 
    7.5678484706028253e-08, 7.2983969894387906e-08, 7.0351545886361651e-08, 
    6.7776680741393912e-08, 6.525563183307539e-08, 6.2785452794301918e-08, 
    6.0363935217692814e-08, 5.7989517649941192e-08, 5.5661189476881265e-08, 
    5.337840684589842e-08, 5.1141026037879958e-08, 4.894924857044712e-08, 
    4.6803565764346422e-08, 4.4704688903724739e-08, 4.2653455731676947e-08, 
    4.0650712297773988e-08, 3.8697180193661964e-08, 3.679332841580937e-08, 
    3.493927554492617e-08, 3.3134747909260296e-08, 3.1379113869004802e-08, 
    2.9671502527313399e-08, 2.8011000523312216e-08, 2.6396904410539546e-08, 
    2.4828993280426795e-08, 2.3307777879684814e-08, 2.1834681878050567e-08, 
    2.041211737128174e-08, 1.9043430400932354e-08, 1.7732710045579029e-08, 
    1.6484474584447909e-08, 1.5303265871401592e-08, 1.4193196966524932e-08, 
    1.3157504433426549e-08, 1.2198156514466214e-08, 1.1315560303105554e-08, 
    1.0508398023628189e-08, 9.7736058508541281e-09, 9.1064918588409058e-09, 
    8.5009744311776148e-09, 7.9499115163971119e-09, 7.4454846716919898e-09, 
    6.979601068081014e-09, 6.5442798287582951e-09, 6.1319960420966949e-09, 
    5.7359638942799238e-09, 5.350349189139138e-09, 4.9704087461485532e-09, 
    4.5925600688069163e-09, 4.2143879865916175e-09, 3.8345969275065064e-09, 
    3.4529175619185408e-09, 3.0699763812286368e-09, 2.687136155113939e-09, 
    2.3063152812550249e-09, 1.9297941816059821e-09, 1.5600180018279161e-09, 
    1.1994053759903927e-09, 8.5017387606131157e-10, 5.1419218910795167e-10, 
    1.9286805088897455e-10, -1.1292165228516371e-10, -4.0285527492045938e-10, 
    -6.7714599933190612e-10, -9.364808995705474e-10, -1.1819272929867273e-09, 
    -1.4148162026832278e-09, -1.6366141109618877e-09, 
    -1.8487936293355527e-09, -2.0527127424155256e-09, -2.249509895709891e-09, 
    -2.4400202765184357e-09, -2.6247161001131955e-09, 
    -2.8036723586721748e-09, -2.976558002195086e-09, -3.1426520990850761e-09, 
    -3.3008838693177418e-09, -3.4498952178360141e-09, 
    -3.5881234824687847e-09, -3.7139011243255584e-09, 
    -3.8255673947379179e-09, -3.9215855443122976e-09, 
    -4.0006574243400192e-09, -4.0618267296186548e-09, 
    -4.1045619493857642e-09, -4.1288115461959225e-09, 
    -4.1350259536277771e-09, -4.1241443484925973e-09, 
    -4.0975474705914812e-09, -4.0569813644776247e-09, 
    -4.0044594421100426e-09, -3.9421521679649984e-09, -3.872273913408421e-09, 
    -3.796976084401597e-09, -3.7182537307544283e-09, -3.6378709992982926e-09, 
    -3.5573082959791212e-09, -3.4777322851468832e-09, 
    -3.3999880897479712e-09, -3.3246122969968266e-09, -3.251864537249638e-09, 
    -3.1817752510527746e-09, -3.1142065957447657e-09, 
    -3.0489231378842988e-09, -2.9856679054026121e-09, 
    -2.9242387577684955e-09, -2.8645589663543065e-09, 
    -2.8067357501125111e-09, -2.751100448010537e-09, -2.6982253348843995e-09, 
    -2.6489135883725298e-09, -2.6041617338862929e-09, -2.56509649345694e-09, 
    -2.5328910939254398e-09, -2.5086682405406984e-09, 
    -2.4933988788704494e-09, -2.4878062075149433e-09, 
    -2.4922842122697327e-09, -2.5068381892058404e-09, 
    -2.5310527351003057e-09, -2.5640897727647565e-09, 
    -2.6047165568319533e-09, -2.6513608625770758e-09, 
    -2.7021887303193021e-09, -2.7551984188350366e-09, 
    -2.8083237642402059e-09, -2.8595396392883268e-09, 
    -2.9069628795242922e-09, -2.9489424659887026e-09, -2.98413401429574e-09, 
    -3.0115545106256451e-09, -3.0306147496841746e-09, 
    -3.0411280211149415e-09, -3.0432952623782816e-09, 
    -3.0376680148169444e-09, -3.0250922010942522e-09, 
    -3.0066367330157673e-09, -2.9835122753188823e-09, 
    -2.9569859218142616e-09, -2.9282981107941744e-09, 
    -2.8985875974785005e-09, -2.8688298331291095e-09, 
    -2.8397925800951527e-09, -2.8120112952297947e-09, 
    -2.7857847544269864e-09, -2.7611898066351722e-09, 
    -2.7381123106088235e-09, -2.7162902821300897e-09, 
    -2.6953642547074706e-09, -2.6749299404143361e-09, 
    -2.6545882689198713e-09, -2.6339889940780225e-09, -2.61286480994758e-09, 
    -2.5910544514981662e-09, -2.5685141645774552e-09, 
    -2.5453182626581265e-09, -2.521649985660247e-09, -2.4977846549065205e-09, 
    -2.4740670458950002e-09, -2.4508852034250597e-09, -2.42864244487615e-09, 
    -2.407729382513921e-09, -2.3884973376982296e-09, -2.3712345659366773e-09, 
    -2.356146310477688e-09, -2.3433398423813041e-09, -2.3328152423467479e-09, 
    -2.3244626518225383e-09, -2.3180662232960878e-09, 
    -2.3133147841811274e-09, -2.3098185370567627e-09, 
    -2.3071308728720939e-09, -2.3047737168924426e-09, 
    -2.3022647983033038e-09, -2.2991448260718489e-09, 
    -2.2950029052637594e-09, -2.2894985678828114e-09, 
    -2.2823794057051544e-09, -2.2734935104988039e-09, -2.262796609765293e-09, 
    -2.25035397270691e-09, -2.2363375316595445e-09, -2.2210185930467767e-09, 
    -2.2047566904125378e-09, -2.1879847829146734e-09, 
    -2.1711912187897011e-09, -2.1548985702282507e-09, 
    -2.1396398363463085e-09, -2.1259325519524861e-09, 
    -2.1142518782484218e-09, -2.1050039770900158e-09, 
    -2.0985015192707641e-09, -2.0949431609592394e-09, 
    -2.0943990255456011e-09, -2.0968037052955619e-09, 
    -2.1019579712527554e-09, -2.1095393780853117e-09, 
    -2.1191213062475649e-09, -2.1301988627556507e-09, 
    -2.1422196225725222e-09, -2.1546164342551546e-09, 
    -2.1668396064726732e-09, -2.1783857620236503e-09, 
    -2.1888213080741376e-09, -2.1977989731329563e-09, 
    -2.2050668534465716e-09, -2.2104699982721319e-09, 
    -2.2139454427292156e-09, -2.2155118847092356e-09, -2.215255633949537e-09, 
    -2.2133143630746366e-09, -2.2098601991923455e-09, 
    -2.2050832680872043e-09, -2.1991767055962516e-09, 
    -2.1923236303085396e-09, -2.1846865595148497e-09, 
    -2.1763993793235418e-09, -2.1675620646463426e-09, -2.158238135679659e-09, 
    -2.1484549660810424e-09, -2.1382068412729997e-09, 
    -2.1274607406044763e-09, -2.1161644875566948e-09, 
    -2.1042569041605143e-09, -2.0916791809198977e-09, 
    -2.0783867065519046e-09, -2.0643601811188508e-09, 
    -2.0496150750317702e-09, -2.0342082978006314e-09, 
    -2.0182413965939997e-09, -2.0018596536854997e-09, 
    -1.9852471197220313e-09, -1.9686177607820539e-09, 
    -1.9522035690352823e-09, -1.9362405187191974e-09, 
    -1.9209537351347587e-09, -1.906543008355765e-09, -1.8931699697220128e-09, 
    -1.8809478125650405e-09, -1.8699343801881208e-09, 
    -1.8601288699907168e-09, -1.8514723753520321e-09, 
    -1.8438518979901676e-09, -1.8371075431663238e-09, 
    -1.8310421652183833e-09, -1.825432920096254e-09, -1.8200438614069193e-09, 
    -1.8146389404463329e-09, -1.8089945837504246e-09, 
    -1.8029112395828169e-09, -1.7962231220289391e-09, 
    -1.7888057119210594e-09, -1.7805804229358938e-09, 
    -1.7715162732570692e-09, -1.7616283809918585e-09, 
    -1.7509735134208124e-09, -1.7396430156573376e-09, 
    -1.7277538133016353e-09, -1.7154381317642894e-09, 
    -1.7028329381719568e-09, -1.690069765620396e-09, -1.6772658384831818e-09, 
    -1.6645168999283169e-09, -1.6518922278533081e-09, 
    -1.6394318470922769e-09, -1.6271460278229289e-09, 
    -1.6150166865218509e-09, -1.6030005476554642e-09, 
    -1.5910336323924876e-09, -1.579036884841638e-09, -1.566922542611307e-09, 
    -1.5546011202446056e-09, -1.5419886370791393e-09, 
    -1.5290139239015981e-09, -1.5156255036998636e-09, 
    -1.5017977333820491e-09, -1.4875355966998079e-09, 
    -1.4728777326790312e-09, -1.4578971616969807e-09, 
    -1.4426994819477683e-09, -1.4274183517087048e-09, 
    -1.4122085358170121e-09, -1.397236852053837e-09, -1.3826718347134286e-09, 
    -1.3686729138974206e-09, -1.3553801603883597e-09, 
    -1.3429054663125839e-09, -1.3313260228936147e-09, -1.320680560881313e-09, 
    -1.3109686847702424e-09, -1.3021531049696762e-09, 
    -1.2941645115647468e-09, -1.2869083611749455e-09, 
    -1.2802729095816763e-09, -1.2741376231331137e-09, 
    -1.2683813152566265e-09, -1.2628892768615972e-09, -1.257559073821533e-09, 
    -1.2523046727136558e-09, -1.247058925989044e-09, -1.2417744098507354e-09, 
    -1.2364229414992204e-09, -1.2309939059668962e-09, 
    -1.2254918048492579e-09, -1.2199331907823634e-09, 
    -1.2143433254777047e-09, -1.208752673040436e-09, -1.2031934752343452e-09, 
    -1.1976964765116881e-09, -1.1922880174432487e-09, 
    -1.1869874908020869e-09, -1.1818054105488107e-09, 
    -1.1767420574396248e-09, -1.1717868991673242e-09, 
    -1.1669187471519152e-09, -1.162106736353146e-09, -1.1573120248726084e-09, 
    -1.1524902005427019e-09, -1.1475941818599906e-09, 
    -1.1425775163132979e-09, -1.1373977810252358e-09, -1.132019922767523e-09, 
    -1.1264192552195954e-09, -1.1205839315613764e-09, 
    -1.1145166452694093e-09, -1.1082354691189316e-09, 
    -1.1017736413610836e-09, -1.0951783454692036e-09, 
    -1.0885084195361308e-09, -1.0818311439492672e-09, 
    -1.0752182232714407e-09, -1.0687412700619867e-09, 
    -1.0624669887704181e-09, -1.0564524889539581e-09, 
    -1.0507410213042932e-09, -1.0453585636311537e-09, 
    -1.0403114937152167e-09, -1.0355856543029621e-09, 
    -1.0311468797254874e-09, -1.0269430590897917e-09, 
    -1.0229075211146303e-09, -1.0189635540212989e-09, 
    -1.0150296367412136e-09, -1.011024983118779e-09, -1.0068749128932648e-09, 
    -1.0025156648324248e-09, -9.9789822533761303e-10, 
    -9.9299100539821936e-10, -9.8778114070446546e-10, 
    -9.8227448977650956e-10, -9.7649436334736439e-10, 
    -9.7047923467801514e-10, -9.6427961681861918e-10, 
    -9.5795444249337023e-10, -9.5156715566198695e-10, 
    -9.4518183410054908e-10, -9.3885949615141135e-10, -9.326548652896546e-10, 
    -9.2661366464164081e-10, -9.2077061937434921e-10, 
    -9.1514819609507217e-10, -9.0975616827783371e-10, 
    -9.0459193707390704e-10, -8.9964162527989621e-10, 
    -8.9488174875392402e-10, -8.9028140011038175e-10, 
    -8.8580467976102498e-10, -8.8141322780843075e-10, 
    -8.7706859513491326e-10, -8.7273434302696896e-10, 
    -8.6837765402868622e-10, -8.639704704455144e-10, -8.5949006311142835e-10, 
    -8.5491917573160499e-10, -8.502457665651654e-10, -8.4546254268530272e-10, 
    -8.405663746451633e-10, -8.3555775963019382e-10, -8.3044036433653327e-10, 
    -8.2522074216060864e-10, -8.1990816921287316e-10, 
    -8.1451457962591857e-10, -8.0905449332461389e-10, 
    -8.0354492398344654e-10, -7.9800508690112196e-10, 
    -7.9245597316319875e-10, -7.8691969595566574e-10, 
    -7.8141868999664003e-10, -7.7597479866659699e-10, 
    -7.7060837677266365e-10, -7.6533744670714689e-10, 
    -7.6017710349096033e-10, -7.5513913422279538e-10, -7.502319965544255e-10, 
    -7.4546108975872364e-10, -7.40829363683614e-10, -7.3633811439194599e-10, 
    -7.3198794808882209e-10, -7.2777974510003203e-10, 
    -7.2371554853010893e-10, -7.1979920768767257e-10, 
    -7.1603676860395128e-10, -7.1243644952958288e-10, 
    -7.0900824274050493e-10, -7.05763097614867e-10, -7.0271177651129744e-10, 
    -6.9986340558575903e-10, -6.9722391655422157e-10, -6.947944249620289e-10, 
    -6.925698158985747e-10, -6.9053757998585175e-10, -6.8867716745110297e-10, 
    -6.8695987989568979e-10, -6.8534946648681312e-10, 
    -6.8380335882681628e-10, -6.8227459018097123e-10, 
    -6.8071418412637728e-10, -6.7907393139364097e-10, 
    -6.7730922647183687e-10, -6.7538181948730316e-10, 
    -6.7326211856600625e-10, -6.7093093207668065e-10, 
    -6.6838040052283703e-10, -6.6561409712941817e-10, 
    -6.6264627096731288e-10, -6.5950036678975355e-10, 
    -6.5620695242469851e-10, -6.5280134361866313e-10, 
    -6.4932109973947732e-10, -6.4580373179698004e-10, 
    -6.4228470898707864e-10, -6.3879602697418004e-10, 
    -6.3536528736518703e-10, -6.3201536887392771e-10, 
    -6.2876453623125477e-10, -6.2562691195001835e-10, 
    -6.2261308949417967e-10, -6.1973080306449462e-10, 
    -6.1698542470567957e-10, -6.1438026926146592e-10, 
    -6.1191659526740084e-10, -6.0959335749932582e-10, 
    -6.0740671786158679e-10, -6.0534947202059379e-10, 
    -6.0341043896521172e-10, -6.015740441307115e-10, -5.9982010610624969e-10, 
    -5.9812403417044091e-10, -5.9645739400369807e-10, 
    -5.9478894689905844e-10, -5.9308603474745781e-10, -5.913162978801056e-10, 
    -5.8944953085304039e-10, -5.8745958886003623e-10, 
    -5.8532609975608148e-10, -5.8303589529874031e-10, 
    -5.8058394725082914e-10, -5.7797378939621662e-10, 
    -5.7521728797264249e-10, -5.7233385306574778e-10, 
    -5.6934907556227139e-10, -5.6629299166447609e-10, 
    -5.6319804001594704e-10, -5.6009697296359748e-10, 
    -5.5702083184002882e-10, -5.5399723178957332e-10, 
    -5.5104900004065941e-10, -5.4819335588674827e-10, 
    -5.4544157002110923e-10, -5.4279917570166265e-10, 
    -5.4026656856827739e-10, -5.3783997071351943e-10, 
    -5.3551254517774106e-10, -5.3327557279508378e-10, 
    -5.3111950163474574e-10, -5.2903482230272736e-10, 
    -5.2701262408818292e-10, -5.2504486976529697e-10, 
    -5.2312434502622532e-10, -5.2124440546716631e-10, 
    -5.1939853442415478e-10, -5.1757988670416379e-10, 
    -5.1578084325965334e-10, -5.1399274490214611e-10, 
    -5.1220578739465569e-10, -5.1040916815986292e-10, 
    -5.0859141277914878e-10, -5.067409263764018e-10, -5.0484660515472139e-10, 
    -5.02898520374502e-10, -5.0088852999927341e-10, -4.9881083197419468e-10, 
    -4.9666231441282067e-10, -4.9444278270311641e-10, 
    -4.9215496427855612e-10, -4.898044002690815e-10, -4.8739916591511611e-10, 
    -4.8494951587960709e-10, -4.8246743379682231e-10, 
    -4.7996617477002091e-10, -4.7745973033679968e-10, 
    -4.7496231116914011e-10, -4.7248777639815351e-10, -4.700490959110759e-10, 
    -4.6765777739296189e-10, -4.6532335370340277e-10, 
    -4.6305289605192196e-10, -4.6085065438926064e-10, 
    -4.5871778802537039e-10, -4.5665233013067914e-10, 
    -4.5464929536573107e-10, -4.5270104011210834e-10, 
    -4.5079780997922758e-10, -4.489284802351698e-10, -4.4708140245755732e-10, 
    -4.4524532814896052e-10, -4.4341028204472867e-10, 
    -4.4156835405306707e-10, -4.3971426561956929e-10, 
    -4.3784572684382449e-10, -4.3596345315236109e-10, 
    -4.3407093102833221e-10, -4.321738555384685e-10, -4.3027937171250739e-10, 
    -4.2839513333041031e-10, -4.2652832177344901e-10, 
    -4.2468467532830521e-10, -4.22867693155192e-10, -4.2107802337508428e-10, 
    -4.1931315966135214e-10, -4.1756743503536046e-10, 
    -4.1583234854773024e-10, -4.1409714336719458e-10, 
    -4.1234965212243018e-10, -4.1057723977108004e-10, 
    -4.0876783610844378e-10, -4.0691090171533707e-10, 
    -4.0499830767271521e-10, -4.0302500238100327e-10, 
    -4.0098946958714288e-10, -3.9889391825854906e-10, 
    -3.9674425124309837e-10, -3.9454977479339404e-10, 
    -3.9232275900620881e-10, -3.9007781940731829e-10, 
    -3.8783122916990719e-10, -3.8560016110837025e-10, 
    -3.8340196132165417e-10, -3.8125341490400405e-10, 
    -3.7917008594855123e-10, -3.771657170946359e-10, -3.7525171768033093e-10, 
    -3.7343671606155263e-10, -3.7172621423399245e-10, 
    -3.7012230045042995e-10, -3.6862349712191997e-10, 
    -3.6722466460268018e-10, -3.6591705557934575e-10, 
    -3.6468847373084468e-10, -3.635235953443635e-10, -3.6240443528594162e-10, 
    -3.6131097199456401e-10, -3.6022189968987325e-10, 
    -3.5911553638102442e-10, -3.5797075023479236e-10, 
    -3.5676798947741251e-10, -3.5549020571272938e-10, 
    -3.5412374167800409e-10, -3.5265902444810685e-10, 
    -3.5109109495120771e-10, -3.4941986461238248e-10, 
    -3.4765015330466924e-10, -3.4579143829644165e-10, -3.438573818050573e-10, 
    -3.4186512181806798e-10, -3.3983439242880289e-10, 
    -3.3778648046750812e-10, -3.3574310749159947e-10, 
    -3.3372523747186157e-10, -3.3175191513543425e-10, 
    -3.2983915414079083e-10, -3.2799898213955173e-10, 
    -3.2623867222691969e-10, -3.2456027355841599e-10, 
    -3.2296044227511115e-10, -3.2143068044965153e-10, -3.199579393212244e-10, 
    -3.1852558331534185e-10, -3.1711466289254734e-10, 
    -3.1570542311999877e-10, -3.1427886552751731e-10, 
    -3.1281831996280425e-10, -3.1131078994300414e-10, 
    -3.0974804182134753e-10, -3.0812725348489553e-10, 
    -3.0645125830755278e-10, -3.0472828602308268e-10, -3.029713001428819e-10, 
    -3.0119696490826989e-10, -2.9942438292282704e-10, 
    -2.9767368846333341e-10, -2.9596468253214372e-10, 
    -2.9431556402664765e-10, -2.9274192383245815e-10, 
    -2.9125600714908122e-10, -2.8986634905284137e-10, -2.885777099190859e-10, 
    -2.8739132325658387e-10, -2.8630535397902178e-10, 
    -2.8531551816001986e-10, -2.8441573570790387e-10, 
    -2.8359876210818414e-10, -2.82856702362248e-10, -2.8218139362406608e-10, 
    -2.8156460103293954e-10, -2.8099809745092272e-10, 
    -2.8047360042748691e-10, -2.7998269531669309e-10, 
    -2.7951672662576417e-10, -2.7906680798047121e-10, 
    -2.7862388051050825e-10, -2.7817894049403693e-10, 
    -2.7772334088446911e-10, -2.7724917866889229e-10, 
    -2.7674968359244966e-10, -2.7621959225736094e-10, 
    -2.7565538853403769e-10, -2.7505543247900574e-10, 
    -2.7441990065329752e-10, -2.7375058445149615e-10, -2.730505427659337e-10, 
    -2.7232367183550433e-10, -2.7157422175602483e-10, 
    -2.7080633784666813e-10, -2.7002363732527866e-10, -2.692288813439683e-10, 
    -2.6842372709021364e-10, -2.676085891281416e-10, -2.6678256016914775e-10, 
    -2.6594343063971532e-10, -2.6508775069528829e-10, 
    -2.6421095836544892e-10, -2.6330755758351321e-10, 
    -2.6237139951628156e-10, -2.6139600646071668e-10, 
    -2.6037503007370998e-10, -2.5930275814871319e-10, 
    -2.5817471699119895e-10, -2.5698827677112969e-10, 
    -2.5574325245864914e-10, -2.5444239130071918e-10, -2.530917282841851e-10, 
    -2.5170070283236096e-10, -2.5028205125197464e-10, 
    -2.4885139618170281e-10, -2.4742661290903316e-10, 
    -2.4602695498149551e-10, -2.4467204902023783e-10, 
    -2.4338081155092103e-10, -2.4217040224428206e-10, 
    -2.4105527754935631e-10, -2.4004644167299474e-10, 
    -2.3915092176734615e-10, -2.3837152860138406e-10, -2.37706857814271e-10, 
    -2.3715157367946218e-10, -2.3669685797398295e-10, 
    -2.3633102743137795e-10, -2.3604021937580319e-10, 
    -2.3580911467759925e-10, -2.3562160303259561e-10, 
    -2.3546138824851451e-10, -2.3531246390869969e-10, 
    -2.3515948592103896e-10, -2.3498799370538287e-10, -2.347845618349731e-10, 
    -2.3453682817387156e-10, -2.342335149116044e-10, -2.3386440209770673e-10, 
    -2.3342036559647894e-10, -2.3289343624126129e-10, 
    -2.3227694360563985e-10, -2.3156572622268272e-10, 
    -2.3075640885402219e-10, -2.2984770223361368e-10, 
    -2.2884070621621016e-10, -2.277391558507006e-10, -2.2654958108052923e-10, 
    -2.2528131183529224e-10, -2.2394634309121905e-10, 
    -2.2255899142260849e-10, -2.2113539130502547e-10, -2.196928293630134e-10, 
    -2.1824896560204802e-10, -2.1682099046976546e-10, 
    -2.1542478831728181e-10, -2.1407415927317554e-10, 
    -2.1278017338595462e-10, -2.1155070716993194e-10, 
    -2.1039020941421922e-10, -2.0929969485233841e-10, 
    -2.0827703577865562e-10, -2.0731744592463762e-10, -2.064142035746794e-10, 
    -2.0555950563753866e-10, -2.0474540968869077e-10, 
    -2.0396477136554035e-10, -2.0321209846036755e-10, 
    -2.0248423249820044e-10, -2.0178079144748848e-10, 
    -2.0110430987719005e-10, -2.0046007704425541e-10, 
    -1.9985562150231574e-10, -1.9929993433293697e-10, 
    -1.9880245028410424e-10, -1.9837190090164759e-10, 
    -1.9801514033640734e-10, -1.977360604272489e-10, -1.975347067748137e-10, 
    -1.9740671038008545e-10, -1.973430794353674e-10, -1.9733040551692295e-10, 
    -1.9735147717263044e-10, -1.9738625052430786e-10, 
    -1.9741309595771584e-10, -1.9741021864605864e-10, 
    -1.9735710931849213e-10, -1.97235912162885e-10, -1.9703256484395082e-10, 
    -1.9673765707237318e-10, -1.9634689961760766e-10, -1.958611984816206e-10, 
    -1.9528635433545793e-10, -1.9463242552886509e-10, 
    -1.9391283401420822e-10, -1.931433036015824e-10, -1.9234073486858186e-10, 
    -1.9152211296505219e-10, -1.9070351149391571e-10, 
    -1.8989928167398224e-10, -1.891214345964323e-10, -1.8837925454608652e-10, 
    -1.876791244290856e-10, -1.8702454475281214e-10, -1.8641630981289851e-10, 
    -1.8585279699180374e-10, -1.8533034499052292e-10, 
    -1.8484363667006051e-10, -1.8438610997000631e-10, -1.839503265307284e-10, 
    -1.835282920254073e-10, -1.8311175207954632e-10, -1.8269241959195306e-10, 
    -1.8226217418446244e-10, -1.8181324714649701e-10, 
    -1.8133839668089439e-10, -1.8083109096842778e-10, 
    -1.8028572613726515e-10, -1.7969784807256246e-10, 
    -1.7906438243741699e-10, -1.7838386408492104e-10, 
    -1.7765661731501611e-10, -1.7688486821771221e-10, 
    -1.7607274225825694e-10, -1.7522612925899811e-10, 
    -1.7435239566127022e-10, -1.734599379194728e-10, -1.7255759967844649e-10, 
    -1.7165399286584138e-10, -1.7075676778222142e-10, 
    -1.6987191810291012e-10, -1.6900318267987319e-10, 
    -1.6815162636736635e-10, -1.6731545824512825e-10, 
    -1.6649011994645275e-10, -1.6566868685875964e-10, 
    -1.6484253873736573e-10, -1.6400225857024195e-10, 
    -1.6313869181478445e-10, -1.6224408372398852e-10, 
    -1.6131314712427047e-10, -1.6034398537760214e-10, -1.593387654257619e-10, 
    -1.5830405056159516e-10, -1.5725074597151943e-10, 
    -1.5619367450786475e-10, -1.5515075719435895e-10, 
    -1.5414190612966252e-10, -1.5318769316965396e-10, 
    -1.5230791400741613e-10, -1.5152017901529335e-10, 
    -1.5083863610421194e-10, -1.5027292850171702e-10, 
    -1.4982750507028423e-10, -1.495012738594182e-10, -1.4928766498735931e-10, 
    -1.4917505189066966e-10, -1.4914749527578088e-10, 
    -1.4918572635990497e-10, -1.4926827851532884e-10, 
    -1.4937268582948484e-10, -1.4947664693824153e-10, 
    -1.4955908392654469e-10, -1.4960104211898714e-10, 
    -1.4958639476632925e-10, -1.4950234163044413e-10, 
    -1.4933968709306548e-10, -1.4909295564862073e-10, 
    -1.4876031446085161e-10, -1.4834338971290443e-10, 
    -1.4784695254858376e-10, -1.4727855771144537e-10, 
    -1.4664809743021037e-10, -1.4596734057442216e-10, 
    -1.4524943618787937e-10, -1.4450841868507494e-10, 
    -1.4375870301798162e-10, -1.4301460216122245e-10, -1.422898519095342e-10, 
    -1.4159718617627754e-10, -1.4094792952262489e-10, 
    -1.4035165732376824e-10, -1.3981588779525178e-10, 
    -1.3934585759413211e-10, -1.3894434464241146e-10, 
    -1.3861156751267223e-10, -1.383451654513074e-10, -1.3814026738408431e-10, 
    -1.3798964170925601e-10, -1.3788395890399213e-10, 
    -1.3781212630012445e-10, -1.3776173446812253e-10, 
    -1.3771953743399241e-10, -1.3767201614012879e-10, 
    -1.3760590051656296e-10, -1.3750871019487588e-10, 
    -1.3736917903061301e-10, -1.3717762088632988e-10, 
    -1.3692612574711544e-10, -1.3660867216233855e-10, 
    -1.3622106632188297e-10, -1.3576082189189709e-10, 
    -1.3522693673118214e-10, -1.346196849762384e-10, -1.3394038428768767e-10, 
    -1.3319126549593462e-10, -1.3237537316538726e-10, 
    -1.3149659101100526e-10, -1.3055969560262007e-10, 
    -1.2957050120693523e-10, -1.2853596338097833e-10, 
    -1.2746428896181329e-10, -1.2636492000154015e-10, 
    -1.2524846534028232e-10, -1.241264483649334e-10, -1.2301099415805244e-10, 
    -1.2191436570762859e-10, -1.2084848580924209e-10, 
    -1.1982439406912316e-10, -1.188518032144872e-10, -1.1793866653494864e-10, 
    -1.1709093620610089e-10, -1.1631240749114718e-10, 
    -1.1560474949301068e-10, -1.1496763811108066e-10, 
    -1.1439904347430228e-10, -1.1389553656322118e-10, 
    -1.1345269624023172e-10, -1.1306544199845825e-10, 
    -1.1272841627456739e-10, -1.1243623866141427e-10, 
    -1.1218375403281121e-10, -1.1196617570094138e-10, 
    -1.1177921616341155e-10, -1.1161912921552909e-10, 
    -1.1148277014848549e-10, -1.1136758008693235e-10, 
    -1.1127159901365737e-10, -1.1119340305587282e-10, 
    -1.1113206165472664e-10, -1.110869830153743e-10, -1.110577809939268e-10, 
    -1.1104401861264606e-10, -1.1104495492422066e-10, 
    -1.1105922331204652e-10, -1.1108456258880639e-10, 
    -1.1111753211255448e-10, -1.1115339200107632e-10, 
    -1.1118603921591452e-10, -1.1120816502212888e-10, 
    -1.1121153468547758e-10, -1.1118749003058245e-10, 
    -1.1112754033066347e-10, -1.1102407664173643e-10, 
    -1.1087107323690829e-10, -1.1066476416758695e-10, 
    -1.1040412983541248e-10, -1.1009123773060155e-10, -1.09731271225127e-10, 
    -1.093323152866306e-10, -1.0890483956094934e-10, -1.0846097488076205e-10, 
    -1.0801357135000487e-10, -1.0757520948316962e-10, 
    -1.0715717137857438e-10, -1.0676853369809791e-10, 
    -1.0641540931408125e-10, -1.0610048685165418e-10, 
    -1.0582280643944971e-10, -1.0557789636204617e-10, 
    -1.0535816595304984e-10, -1.0515359447064444e-10, 
    -1.0495257299229958e-10, -1.0474292439707232e-10, 
    -1.0451289613923276e-10, -1.04252152461799e-10, -1.0395259335560685e-10, 
    -1.0360901382826635e-10, -1.0321948917113589e-10, 
    -1.0278551092487528e-10, -1.0231182441305922e-10, 
    -1.0180603981226383e-10, -1.0127798902071523e-10, 
    -1.0073895751273157e-10, -1.0020077752723696e-10, -9.967494401434149e-11, 
    -9.9171744636760137e-11, -9.8699536030758074e-11, 
    -9.8264171862629362e-11, -9.7868683819769374e-11, -9.75131681992283e-11, 
    -9.719494194496514e-11, -9.6908896545217128e-11, -9.6648064419848358e-11, 
    -9.6404291056153156e-11, -9.6169014175809499e-11, 
    -9.5934032562030491e-11, -9.569225089598352e-11, -9.5438296632477167e-11, 
    -9.516904072448625e-11, -9.4883895408544756e-11, -9.4584955341831195e-11, 
    -9.4276906262248573e-11, -9.3966775040004024e-11, 
    -9.3663464478147797e-11, -9.3377171760115297e-11, 
    -9.3118671385061195e-11, -9.2898559513914505e-11, 
    -9.2726475533025274e-11, -9.2610384519425435e-11, -9.2555942162544e-11, 
    -9.2566044302902348e-11, -9.2640517681375913e-11, 
    -9.2776063447268277e-11, -9.2966358923551685e-11, 
    -9.3202398144793443e-11, -9.3472945384247446e-11, 
    -9.3765141821952724e-11, -9.4065148246938133e-11, 
    -9.4358830282359919e-11, -9.4632387465995522e-11, -9.487296184663426e-11, 
    -9.5069132124290496e-11, -9.5211346359513569e-11, 
    -9.5292232443604255e-11, -9.5306864587322731e-11, -9.525291404783903e-11, 
    -9.5130723463867839e-11, -9.4943289099692934e-11, 
    -9.4696186718441765e-11, -9.439734494996381e-11, -9.4056750634930404e-11, 
    -9.3686017465803817e-11, -9.3297891213958428e-11, 
    -9.2905640240495637e-11, -9.2522439426413415e-11, -9.216072331578644e-11, 
    -9.1831604540733307e-11, -9.1544351305603414e-11, 
    -9.1306026894047204e-11, -9.1121234585551804e-11, 
    -9.0992057226732615e-11, -9.0918115128955634e-11, 
    -9.0896784761920801e-11, -9.0923490916773572e-11, 
    -9.0992099367299603e-11, -9.1095299695430821e-11, -9.12250252602351e-11, 
    -9.1372812277561564e-11, -9.1530143714918482e-11, 
    -9.1688718229777053e-11, -9.1840688061006314e-11, 
    -9.1978830988192739e-11, -9.2096702694159585e-11, 
    -9.2188727172138369e-11, -9.2250301415592992e-11, 
    -9.2277831352852074e-11, -9.2268772468794386e-11, 
    -9.2221622272257372e-11, -9.2135907581212112e-11, 
    -9.2012112224826545e-11, -9.1851611049043297e-11, 
    -9.1656546302373579e-11, -9.1429722188877305e-11, 
    -9.1174463504982447e-11, -9.089450782308473e-11, -9.05938890500361e-11, 
    -9.0276866417703899e-11, -8.9947847016411019e-11, 
    -8.9611373001893532e-11, -8.9272089349743133e-11, 
    -8.8934749993592451e-11, -8.8604190279709442e-11, -8.828532244058934e-11, 
    -8.7983068051842592e-11, -8.7702278461127137e-11, 
    -8.7447588634765538e-11, -8.722327080445867e-11, -8.7033008603601138e-11, 
    -8.6879682321598334e-11, -8.6765123979742247e-11, 
    -8.6689889229013658e-11, -8.6653034282674175e-11, -8.665198102008439e-11, 
    -8.6682390326206121e-11, -8.6738152920803766e-11, -8.681143552690383e-11, 
    -8.6892862187558623e-11, -8.6971752507344781e-11, 
    -8.7036497010030448e-11, -8.7074980394082539e-11, 
    -8.7075108631530314e-11, -8.7025344033800561e-11, 
    -8.6915276530184615e-11, -8.6736136757884443e-11, 
    -8.6481275965607454e-11, -8.6146510074420635e-11, 
    -8.5730353866301138e-11, -8.5234079706532192e-11, 
    -8.4661659523788551e-11, -8.4019523491974665e-11, 
    -8.3316220057091145e-11, -8.2561974934331275e-11, 
    -8.1768219989781695e-11, -8.0947079314954126e-11, 
    -8.0110933776723148e-11, -7.9271998922729167e-11, 
    -7.8441994744594283e-11, -7.7631877676141826e-11, 
    -7.6851679116980611e-11, -7.6110365812823827e-11, 
    -7.5415772472918413e-11, -7.4774538501909905e-11, 
    -7.4192100090148536e-11, -7.3672661881975946e-11, 
    -7.3219197387314154e-11, -7.2833455678029834e-11, 
    -7.2516010443878839e-11, -7.2266312705725467e-11, 
    -7.2082799574040771e-11, -7.1963010229788094e-11, 
    -7.1903749490431538e-11, -7.1901235002885413e-11, 
    -7.1951252746037303e-11, -7.2049279244414167e-11, 
    -7.2190554791910673e-11, -7.2370097348044814e-11, -7.258267358036603e-11, 
    -7.2822677531700093e-11, -7.3084012222621662e-11, 
    -7.3359911532842272e-11, -7.3642807292698947e-11, 
    -7.3924231157759338e-11, -7.4194804794789744e-11, 
    -7.4444323070858034e-11, -7.4661987329687135e-11, 
    -7.4836731129555228e-11, -7.4957674268195924e-11, 
    -7.5014625867321603e-11, -7.4998663235470943e-11, 
    -7.4902645809836034e-11, -7.4721693286602046e-11, -7.445352413310298e-11, 
    -7.4098675230788456e-11, -7.3660523408764669e-11, 
    -7.3145170121133871e-11, -7.2561152934345427e-11, 
    -7.1919073234406594e-11, -7.1231120716782176e-11, 
    -7.0510596663632626e-11, -6.9771422356676314e-11, 
    -6.9027720997819645e-11, -6.8293433122495692e-11, 
    -6.7582016896784528e-11, -6.6906188138012295e-11, 
    -6.6277722827186176e-11, -6.5707254505442344e-11, 
    -6.5204098702837859e-11, -6.4776044324807873e-11, 
    -6.4429155274902168e-11, -6.4167540635065148e-11, 
    -6.3993180532463919e-11, -6.3905758787525505e-11, 
    -6.3902588057772712e-11, -6.3978618622790718e-11, 
    -6.4126581907066446e-11, -6.4337229351579165e-11, 
    -6.4599709886236211e-11, -6.4902020998211403e-11, -6.523154246151113e-11, 
    -6.557555681557876e-11, -6.5921803893640818e-11, -6.6258926102857376e-11, 
    -6.6576852160491518e-11, -6.6867051887147557e-11, -6.712269537965943e-11, 
    -6.7338658288465717e-11, -6.7511468764609326e-11, 
    -6.7639130877341401e-11, -6.7720935076989697e-11, 
    -6.7757200439174634e-11, -6.7749063809827301e-11, 
    -6.7698240451818628e-11, -6.7606850871395475e-11, -6.747726042242522e-11, 
    -6.731197416966962e-11, -6.7113543343890127e-11, -6.6884522205483883e-11, 
    -6.6627410033483636e-11, -6.6344627568707689e-11, 
    -6.6038470249036883e-11, -6.5711078144670542e-11, 
    -6.5364372952137512e-11, -6.5000033341430994e-11, 
    -6.4619433095106766e-11, -6.4223614263694844e-11, 
    -6.3813254950044413e-11, -6.3388676703044725e-11, 
    -6.2949857497621156e-11, -6.2496481474202232e-11, 
    -6.2027998792036615e-11, -6.1543725199813943e-11, 
    -6.1042934568093767e-11, -6.0524977515313203e-11, 
    -5.9989387675939187e-11, -5.943599778201606e-11, -5.8865045554935454e-11, 
    -5.8277253026118566e-11, -5.7673907319215254e-11, 
    -5.7056922484775138e-11, -5.642886804650585e-11, -5.5792988589267876e-11, 
    -5.5153183675270948e-11, -5.451396875067717e-11, -5.3880394124637591e-11, 
    -5.3257943502999122e-11, -5.2652391435958037e-11, 
    -5.2069656393072915e-11, -5.1515631177819829e-11, 
    -5.0996012798301589e-11, -5.0516146105312818e-11, 
    -5.0080895254552364e-11, -4.9694527265826168e-11, 
    -4.9360654343699555e-11, -4.908218107786737e-11, -4.8861289276436194e-11, 
    -4.8699424045968612e-11, -4.8597295635676806e-11, 
    -4.8554851134907192e-11, -4.8571231951048596e-11, 
    -4.8644711072628363e-11, -4.8772589057061392e-11, 
    -4.8951092154407543e-11, -4.9175263247591724e-11, 
    -4.9438871113543516e-11, -4.9734376050520235e-11, -5.005294987262779e-11, 
    -5.0384583769957402e-11, -5.0718293941973472e-11, 
    -5.1042433020273914e-11, -5.1345089743755407e-11, 
    -5.1614570904001979e-11, -5.1839944574076579e-11, 
    -5.2011587504718999e-11, -5.212172945170536e-11, -5.2164938107716575e-11, 
    -5.2138502080029086e-11, -5.2042686551424027e-11, 
    -5.1880822393050962e-11, -5.1659245944131501e-11, 
    -5.1387042025235033e-11, -5.1075625857622644e-11, 
    -5.0738199833198789e-11, -5.0389076989977231e-11, 
    -5.0042962791762309e-11, -4.9714201160300343e-11, 
    -4.9416057240057372e-11, -4.9160078020200605e-11, 
    -4.8955558238554817e-11, -4.8809154731191473e-11, 
    -4.8724662538203803e-11, -4.8702965223940807e-11, 
    -4.8742150334239902e-11, -4.8837775655724468e-11, 
    -4.8983266518900215e-11, -4.9170428091651371e-11, 
    -4.9390010719829691e-11, -4.9632315136117907e-11, 
    -4.9887809016134388e-11, -5.0147678786580094e-11, -5.040433535158149e-11, 
    -5.0651825923237505e-11, -5.0886114668248615e-11, 
    -5.1105235621108765e-11, -5.1309301436359899e-11, 
    -5.1500373632821537e-11, -5.1682185914614764e-11, 
    -5.1859763699750539e-11, -5.203893293804761e-11, -5.2225780867782344e-11, 
    -5.2426079291939663e-11, -5.2644723592524354e-11, 
    -5.2885222770933047e-11, -5.3149276275047074e-11, -5.343646722017661e-11, 
    -5.3744108225200891e-11, -5.4067219704748684e-11, 
    -5.4398688301375281e-11, -5.4729563496320253e-11, 
    -5.5049472094136448e-11, -5.534712663817572e-11, -5.5610915420798307e-11, 
    -5.5829484062601134e-11, -5.5992298587282784e-11, 
    -5.6090159515056447e-11, -5.611561306323188e-11, -5.6063256210689665e-11, 
    -5.5929948858764162e-11, -5.5714883018395206e-11, 
    -5.5419580478705399e-11, -5.5047801797509932e-11, -5.460540426443975e-11, 
    -5.4100156824137957e-11, -5.3541551297577857e-11, 
    -5.2940586522313158e-11, -5.2309539506745426e-11, 
    -5.1661707429670021e-11, -5.1011135539469886e-11, 
    -5.0372262970380437e-11, -4.9759527277501928e-11, 
    -4.9186896219347301e-11, -4.8667362526475768e-11, 
    -4.8212402517660469e-11, -4.7831450617815307e-11, 
    -4.7531427943091098e-11, -4.7316395987163073e-11, 
    -4.7187339321504989e-11, -4.7142163146874764e-11, 
    -4.7175887848687285e-11, -4.7281060015543805e-11, 
    -4.7448352873790534e-11, -4.7667298130515755e-11, 
    -4.7927108977655068e-11, -4.8217501582160662e-11, 
    -4.8529438926656685e-11, -4.8855749174566686e-11, 
    -4.9191515891031565e-11, -4.953425077006659e-11, -4.9883809411558106e-11, 
    -5.0242051019631711e-11, -5.0612305942262134e-11, 
    -5.0998692762464993e-11, -5.1405333136641094e-11, 
    -5.1835589075310322e-11, -5.2291330190828422e-11, 
    -5.2772364715769197e-11, -5.3276041508653177e-11, -5.379706698213742e-11, 
    -5.4327569518334779e-11, -5.4857396210888793e-11, 
    -5.5374608860261836e-11, -5.5866144151439697e-11, 
    -5.6318573846221647e-11, -5.6718925493084902e-11, 
    -5.7055451729879291e-11, -5.7318333835586631e-11, 
    -5.7500225992060601e-11, -5.7596616073313649e-11, 
    -5.7605974640442377e-11, -5.75296923659947e-11, -5.737180714110995e-11, 
    -5.7138571359734636e-11, -5.6837880416173971e-11, 
    -5.6478645855478786e-11, -5.6070139464004227e-11, -5.562139172454452e-11, 
    -5.5140670994078443e-11, -5.4635093767424874e-11, 
    -5.4110367266456239e-11, -5.3570700121518421e-11, -5.301883521964304e-11, 
    -5.2456227872735483e-11, -5.1883303495829766e-11, 
    -5.1299797256918685e-11, -5.0705115192748285e-11, -5.009871974711944e-11, 
    -4.9480479188334697e-11, -4.8850994316891985e-11, 
    -4.8211856515116754e-11, -4.7565841143648922e-11, 
    -4.6917009566380566e-11, -4.6270738440587354e-11, 
    -4.5633621890457827e-11, -4.5013296062167015e-11, 
    -4.4418133990901371e-11, -4.3856856255081587e-11, 
    -4.3338048453320095e-11, -4.2869619766748894e-11, 
    -4.2458224411156021e-11, -4.2108714345834415e-11, 
    -4.1823651605820197e-11, -4.1602923553991754e-11, 
    -4.1443531049510951e-11, -4.1339591866369508e-11, 
    -4.1282540515634019e-11, -4.1261567942850966e-11, 
    -4.1264255291485209e-11, -4.127737669343141e-11, -4.1287790394866379e-11, 
    -4.1283362925943762e-11, -4.1253822337053135e-11, 
    -4.1191493541080343e-11, -4.109181739455538e-11, -4.0953631313678754e-11, 
    -4.0779161816453457e-11, -4.0573747293146935e-11, -4.034530474733646e-11, 
    -4.0103585737106987e-11, -3.9859291456410974e-11, 
    -3.9623124512081275e-11, -3.9404842971111588e-11, 
    -3.9212419425303475e-11, -3.905134544958406e-11, -3.8924169405427845e-11, 
    -3.8830274429461285e-11, -3.8765939550484058e-11, 
    -3.8724639846479026e-11, -3.8697610519155247e-11, 
    -3.8674556400857173e-11, -3.8644519893262333e-11, 
    -3.8596762067679465e-11, -3.8521634733665304e-11, 
    -3.8411342493775959e-11, -3.8260570294688113e-11, 
    -3.8066880958668835e-11, -3.7830938965091439e-11, 
    -3.7556481762196969e-11, -3.725012079307072e-11, -3.6920956637435962e-11, 
    -3.6580099086580397e-11, -3.6240095594711523e-11, 
    -3.5914326895965377e-11, -3.5616421795214719e-11, 
    -3.5359686251897946e-11, -3.5156577675522921e-11, 
    -3.5018247846076295e-11, -3.4954117821648187e-11, 
    -3.4971522562231318e-11, -3.5075396174757163e-11, 
    -3.5268045065136674e-11, -3.5548980484290282e-11, 
    -3.5914854087836176e-11, -3.6359496732493653e-11, 
    -3.6874124982607902e-11, -3.7447648906402443e-11, 
    -3.8067153409704156e-11, -3.8718480925892803e-11, 
    -3.9386927584848555e-11, -4.0057970004636088e-11, 
    -4.0718004541347577e-11, -4.135500945280124e-11, -4.1959103838370223e-11, 
    -4.252292877724924e-11, -4.3041856917157383e-11, -4.3513982816216726e-11, 
    -4.3939927544549769e-11, -4.4322479006063413e-11, 
    -4.4666095128900247e-11, -4.4976336548415667e-11, 
    -4.5259292463540376e-11, -4.552101051979144e-11, -4.5767024682525382e-11, 
    -4.6001969982561116e-11, -4.6229335185281732e-11, 
    -4.6451323172520627e-11, -4.6668846907527985e-11, 
    -4.6881611983769809e-11, -4.7088256539155429e-11, 
    -4.7286538791307021e-11, -4.7473546273074031e-11, 
    -4.7645866603421216e-11, -4.7799745358308741e-11, -4.793119029682545e-11, 
    -4.8036050811882157e-11, -4.811005761203846e-11, -4.8148856713291893e-11, 
    -4.8148051092178897e-11, -4.8103262844712373e-11, 
    -4.8010238903176855e-11, -4.7865028489837971e-11, 
    -4.7664193980883324e-11, -4.7405091782777568e-11, 
    -4.7086182795582154e-11, -4.6707347202550159e-11, 
    -4.6270167073130442e-11, -4.5778187646614306e-11, -4.523703959297988e-11, 
    -4.4654473392467758e-11, -4.4040232970562002e-11, 
    -4.3405789560232156e-11, -4.2763925446946559e-11, 
    -4.2128191866216936e-11, -4.1512276446846892e-11, 
    -4.0929328518582921e-11, -4.0391278972795223e-11, 
    -3.9908241802264621e-11, -3.9488001069382618e-11, 
    -3.9135684577029889e-11, -3.8853600237008272e-11, 
    -3.8641263434793628e-11, -3.8495617214695341e-11, 
    -3.8411403023617656e-11, -3.8381633035537159e-11, 
    -3.8398129307049318e-11, -3.8452048658685169e-11, 
    -3.8534363555320621e-11, -3.8636233926568003e-11, 
    -3.8749284490032279e-11, -3.8865748398120373e-11, -3.89785092107716e-11, 
    -3.9081083592117887e-11, -3.9167582413338287e-11, 
    -3.9232681959990179e-11, -3.9271669949226444e-11, 
    -3.9280565372362554e-11, -3.9256324099330361e-11, 
    -3.9197117282863639e-11, -3.9102647613989876e-11, 
    -3.8974442691164888e-11, -3.8816075410977983e-11, -3.863325754327996e-11, 
    -3.8433775387719236e-11, -3.8227222617388053e-11, 
    -3.8024545131253234e-11, -3.7837427638686019e-11, -3.767754919322499e-11, 
    -3.7555790044187727e-11, -3.7481441520679248e-11, 
    -3.7461511266589932e-11, -3.7500165715407023e-11, 
    -3.7598388562532368e-11, -3.7753853356939711e-11, 
    -3.7961050913353396e-11, -3.8211638077001188e-11, 
    -3.8494988885520587e-11, -3.8798888343458369e-11, 
    -3.9110322565790724e-11, -3.9416288923034852e-11, 
    -3.9704574016366679e-11, -3.9964435296937766e-11, 
    -4.0187144215452126e-11, -4.0366367318434707e-11, 
    -4.0498363101083617e-11, -4.0581990555094364e-11, 
    -4.0618554997124969e-11, -4.0611521253814511e-11, 
    -4.0566099999718965e-11, -4.0488778758460728e-11, 
    -4.0386802972928606e-11, -4.0267652578198933e-11, 
    -4.0138538144506707e-11, -4.0005948166810231e-11, -3.987524567395209e-11, 
    -3.9750363347908432e-11, -3.9633570321599262e-11, 
    -3.9525371375159484e-11, -3.9424510812044019e-11, 
    -3.9328100285225165e-11, -3.923188187081946e-11, -3.9130610567501103e-11, 
    -3.9018552745592282e-11, -3.8890032593073474e-11, 
    -3.8740034932720904e-11, -3.8564807887428619e-11, 
    -3.8362381117269268e-11, -3.8132978493723423e-11, 
    -3.7879286647730083e-11, -3.7606528584006617e-11, 
    -3.7322340313759791e-11, -3.703645801029456e-11, -3.676022763503464e-11, 
    -3.6505985380846673e-11, -3.6286354531388109e-11, 
    -3.6113495603249631e-11, -3.5998388295212255e-11, 
    -3.5950188416170885e-11, -3.59756862733414e-11, -3.6078896899814963e-11, 
    -3.6260813353447746e-11, -3.6519312180472447e-11, 
    -3.6849215211564373e-11, -3.7242470229641852e-11, 
    -3.7688464453197756e-11, -3.8174432044048966e-11, 
    -3.8685922237970901e-11, -3.9207326382663542e-11, 
    -3.9722440434697958e-11, -4.0215026743413307e-11, 
    -4.0669389803515728e-11, -4.1070933990408307e-11, 
    -4.1406690274689981e-11, -4.1665796357868085e-11, 
    -4.1839914447078348e-11, -4.1923562584888177e-11, 
    -4.1914337900305172e-11, -4.1813000976770852e-11, 
    -4.1623422989613726e-11, -4.1352357838755236e-11, 
    -4.1009064860375912e-11, -4.0604782847202437e-11, 
    -4.0152101457488487e-11, -3.9664235592995219e-11, 
    -3.9154321128949433e-11, -3.8634726153433888e-11, 
    -3.8116479387764109e-11, -3.7608848273906747e-11, 
    -3.7119096721487783e-11, -3.6652431401544138e-11, 
    -3.6212137383342472e-11, -3.5799852088112061e-11, 
    -3.5415948108847817e-11, -3.5059948170143855e-11, 
    -3.4730931294431366e-11, -3.4427859761595506e-11, 
    -3.4149820871214835e-11, -3.3896125034052783e-11, 
    -3.3666303730550992e-11, -3.3460021496129683e-11, 
    -3.3276919807237468e-11, -3.311647142186945e-11, -3.2977868915195921e-11, 
    -3.2859984102089242e-11, -3.2761441482136053e-11, 
    -3.2680788408139987e-11, -3.2616755437014556e-11, 
    -3.2568579639667541e-11, -3.253633553959793e-11, -3.252121587540208e-11, 
    -3.2525727225975505e-11, -3.2553733728896566e-11, 
    -3.2610333166336182e-11, -3.2701549204929347e-11, -3.283385355862743e-11, 
    -3.3013551675576681e-11, -3.3246084584431327e-11, -3.35353249041183e-11, 
    -3.388292950793531e-11, -3.428782530799989e-11, -3.4745888768766004e-11, 
    -3.5249882031426405e-11, -3.5789636338526978e-11, 
    -3.6352488676814762e-11, -3.69239532891877e-11, -3.7488555533235084e-11, 
    -3.8030763568379255e-11, -3.8535933012026406e-11, -3.899118766863407e-11, 
    -3.9386148714034272e-11, -3.9713466248541487e-11, 
    -3.9969106683320462e-11, -4.0152374465358913e-11, 
    -4.0265688507266435e-11, -4.0314129192157953e-11, 
    -4.0304818370490922e-11, -4.0246180633941194e-11, 
    -4.0147165033415896e-11, -4.0016487746901244e-11, 
    -3.9861952724273361e-11, -3.9689915584376274e-11, 
    -3.9504909346871905e-11, -3.9309463579480155e-11, 
    -3.9104119432028484e-11, -3.8887623329323936e-11, 
    -3.8657280046185292e-11, -3.8409429784667128e-11, 
    -3.8140009672225323e-11, -3.7845139876191157e-11, 
    -3.7521715127174235e-11, -3.7167931921461787e-11, 
    -3.6783727424136569e-11, -3.6371106624306908e-11, 
    -3.5934300295912839e-11, -3.5479788021419677e-11, 
    -3.5016148209661778e-11, -3.4553756202989518e-11, 
    -3.4104347658320407e-11, -3.368046398630555e-11, -3.3294832311687148e-11, 
    -3.2959698730303173e-11, -3.2686174716094348e-11, 
    -3.2483623490007531e-11, -3.2359137609644614e-11, -3.2317142228265973e-11,
  // Sqw-F(5, 0-1999)
    0.032332496205479962, 0.032322570206769402, 0.032292799253829642, 
    0.032243205956153285, 0.032173832660284403, 0.032084747554795678, 
    0.031976051608887911, 0.031847885114634607, 0.031700432724760842, 
    0.031533926244583191, 0.031348644996289976, 0.031144914232563145, 
    0.030923102711660082, 0.030683621024134373, 0.030426922462446417, 
    0.030153508066901317, 0.029863936941385564, 0.029558842057281931, 
    0.029238950670220355, 0.028905107333100113, 0.028558296498734294, 
    0.028199661057588084, 0.027830512997576929, 0.027452332776929305, 
    0.027066754949430623, 0.026675538963794907, 0.02628052569040315, 
    0.025883581880726619, 0.025486536205119984, 0.025091111547045714, 
    0.024698858727936038, 0.02431109675477048, 0.023928864067410113, 
    0.023552884232576683, 0.02318354824927089, 0.022820914272191017, 
    0.022464724282608029, 0.022114436155576372, 0.021769268750314895, 
    0.021428257097126851, 0.021090314439680131, 0.020754297765288039, 
    0.020419073466594172, 0.020083579889375369, 0.019746883719977106, 
    0.019408227461611745, 0.019067065664440767, 0.01872308813288593, 
    0.018376229042981314, 0.018026661744770009, 0.017674779950975508, 
    0.017321166947177714, 0.016966555307135131, 0.016611780264589288, 
    0.016257730299533837, 0.015905298591228974, 0.015555338758958258, 
    0.015208627781538295, 0.014865838220186786, 0.014527520954007049, 
    0.014194098672486381, 0.013865869452825093, 0.013543018966077057, 
    0.01322563926797766, 0.012913751775283469, 0.012607331917728663, 
    0.012306333076910378, 0.012010707744689667, 0.011720424308646173, 
    0.011435478445084853, 0.011155898711155623, 0.010881746517697705, 
    0.010613111179914954, 0.010350101140507939, 0.010092832709999647, 
    0.0098414177589734465, 0.0095959517317770957, 0.0093565031525734074, 
    0.0091231054974897884, 0.0088957519545556918, 0.0086743932320460376, 
    0.0084589382480065173, 0.008249257272469843, 0.0080451869201361922, 
    0.0078465363123276372, 0.0076530937372026675, 0.0074646332206315209, 
    0.0072809205543839855, 0.0071017184885007155, 0.0069267909572990607, 
    0.0067559063538100714, 0.0065888399816210422, 0.0064253758882896967, 
    0.0062653083185687996, 0.0061084430211114545, 0.0059545986049400462, 
    0.0058036080796506871, 0.0056553206350586291, 0.0055096036310636146, 
    0.0053663446860788373, 0.0052254536810798849, 0.0050868644440420704, 
    0.0049505358528689264, 0.0048164520987396637, 0.0046846218885576571, 
    0.0045550764342362224, 0.0044278661736723464, 0.0043030562854287236, 
    0.0041807211848994214, 0.0040609383100760222, 0.0039437816049329973, 
    0.0038293151738308419, 0.0037175876001848563, 0.0036086273909881447, 
    0.0035024399260304732, 0.0033990061641163754, 0.0032982832017877097, 
    0.0032002066110695744, 0.0031046943216181556, 0.0030116516783823496, 
    0.0029209772136308391, 0.0028325686309671008, 0.0027463285105072876, 
    0.0026621693033433095, 0.0025800172785626664, 0.00249981520272836, 
    0.002421523654253232, 0.0023451209896575048, 0.002270602074996212, 
    0.0021979759680800896, 0.0021272627842469404, 0.0020584900026449117, 
    0.0019916884755349197, 0.001926888394710757, 0.0018641154506280511, 
    0.0018033873935996848, 0.0017447111733630205, 0.0016880807935235696, 
    0.0016334759709651899, 0.0015808616383921695, 0.0015301882733382162, 
    0.001481392983385954, 0.0014344012301159882, 0.0013891290386165572, 
    0.0013454855193019398, 0.0013033755263088993, 0.0012627022912030746, 
    0.0012233698988228414, 0.0011852855084352454, 0.0011483612615937866, 
    0.0011125158520425094, 0.0010776757580529784, 0.0010437761513819228, 
    0.0010107614999463213, 0.0009785858760906947, 0.00094721297339198064, 
    0.00091661582728808978, 0.00088677623279803002, 0.00085768385898083702, 
    0.0008293350751002247, 0.00080173152593011562, 0.00077487851953586952, 
    0.00074878331533598892, 0.00072345341831867092, 0.00069889499287892798, 
    0.00067511150450303065, 0.00065210267927334861, 0.00062986384192240184, 
    0.00060838565676064849, 0.00058765425718005184, 0.00056765171375893148, 
    0.0005483567627966267, 0.00052974569957408386, 0.00051179333520138767, 
    0.00049447392215766278, 0.00047776196953515696, 0.00046163289142230713, 
    0.00044606345716001055, 0.00043103203686105314, 0.0004165186567317071, 
    0.00040250489449386747, 0.00038897365480342343, 0.00037590886822665669, 
    0.00036329515606820287, 0.0003511174985538549, 0.00033936093705963196, 
    0.00032801033353967076, 0.00031705020296777516, 0.00030646462796385496, 
    0.00029623725895008818, 0.00028635139803664093, 0.0002767901601471339, 
    0.00026753670047529796, 0.00025857449318709725, 0.00024988764250313952, 
    0.00024146120424770534, 0.00023328149406193444, 0.00022533635818452639, 
    0.00021761538432641493, 0.00021011003383569261, 0.000202813681930994, 
    0.00019572155987397142, 0.00018883060090564875, 0.00018213919977853537, 
    0.00017564690290228322, 0.00016935405168088771, 0.00016326140492431006, 
    0.00015736976692078396, 0.00015167964583700562, 0.00014619096289370559, 
    0.00014090282684828519, 0.00013581338150997989, 0.00013091972718739397, 
    0.00012621791093945793, 0.00012170297589892722, 0.00011736905713387396, 
    0.00011320951057254439, 0.00010921706222652899, 0.0001053839668674175, 
    0.00010170216788480973, 9.8163452703842121e-05, 9.4759600386794959e-05, 
    9.1482519567544617e-05, 8.8324375559537953e-05, 8.5277705423513728e-05, 
    8.2335519228559227e-05, 7.9491385021113436e-05, 7.6739494476851729e-05, 
    7.4074706125127346e-05, 7.1492563565776917e-05, 6.8989287254004505e-05, 
    6.656174008697524e-05, 6.4207368950453092e-05, 6.1924126288675859e-05, 
    5.9710377356740415e-05, 5.756479987148369e-05, 5.5486283150336731e-05, 
    5.3473833487156959e-05, 5.152649152883627e-05, 4.9643265942718665e-05, 
    4.7823085904281355e-05, 4.6064773106366561e-05, 4.436703229139714e-05, 
    4.2728457893322679e-05, 4.1147553343880229e-05, 3.9622758993311676e-05, 
    3.8152484410537199e-05, 3.673514102060331e-05, 3.5369171539171979e-05, 
    3.4053073397480978e-05, 3.2785414231940434e-05, 3.1564838461158723e-05, 
    3.0390064910843375e-05, 2.9259876306307597e-05, 2.8173102170040582e-05, 
    2.7128597192207702e-05, 2.6125217450314192e-05, 2.516179692996951e-05, 
    2.4237126647766169e-05, 2.3349938330421954e-05, 2.2498894105497909e-05, 
    2.1682583067495097e-05, 2.0899524958986109e-05, 2.0148180610338867e-05, 
    1.9426968261650918e-05, 1.8734284485090877e-05, 1.8068528154509592e-05, 
    1.7428125780575699e-05, 1.6811556535782901e-05, 1.6217375420958603e-05, 
    1.5644233249024361e-05, 1.5090892419040592e-05, 1.4556237794475375e-05, 
    1.4039282359354148e-05, 1.3539167676360756e-05, 1.3055159491391178e-05, 
    1.2586639097357012e-05, 1.2133091273362487e-05, 1.1694089741985693e-05, 
    1.126928113589428e-05, 1.0858368436701553e-05, 1.0461094755368645e-05, 
    1.0077228177725619e-05, 9.7065482218634523e-06, 9.3488342650698068e-06, 
    9.0038561191390092e-06, 8.6713667792963527e-06, 8.3510972579717671e-06, 
    8.0427533433706262e-06, 7.7460140943236933e-06, 7.4605318867267795e-06, 
    7.1859338512566088e-06, 6.9218245694973371e-06, 6.6677899130454163e-06, 
    6.4234019047911486e-06, 6.1882244509802296e-06, 5.9618197375324747e-06, 
    5.7437550163166568e-06, 5.5336094394977469e-06, 5.3309805511964326e-06, 
    5.1354900284764688e-06, 4.9467882900606021e-06, 4.7645576615560963e-06, 
    4.5885138969881569e-06, 4.418405993292206e-06, 4.2540143817802417e-06, 
    4.0951477174433609e-06, 3.9416385984291434e-06, 3.7933386199351178e-06, 
    3.6501131953231949e-06, 3.5118365617173212e-06, 3.3783873360113959e-06, 
    3.2496449086316312e-06, 3.1254868695912316e-06, 3.0057875629191863e-06, 
    2.8904177711890312e-06, 2.7792454449494559e-06, 2.6721373168729204e-06, 
    2.5689611772438709e-06, 2.4695885392188891e-06, 2.3738973897796583e-06, 
    2.2817747106625715e-06, 2.1931184650459106e-06, 2.1078387851719646e-06, 
    2.0258581627417557e-06, 1.9471105366855851e-06, 1.8715392831049966e-06, 
    1.7990942304115317e-06, 1.7297279335946569e-06, 1.6633915323412527e-06, 
    1.6000305741096604e-06, 1.5395811986948807e-06, 1.481967050590676e-06, 
    1.4270972153281236e-06, 1.3748653731252292e-06, 1.3251502429781775e-06, 
    1.2778172663381214e-06, 1.2327213676635565e-06, 1.1897105398783251e-06, 
    1.1486299451308215e-06, 1.1093261965081815e-06, 1.0716514947286354e-06, 
    1.035467328700323e-06, 1.000647504999819e-06, 9.67080339574146e-07, 
    9.3466991977011755e-07, 9.033364184019279e-07, 8.7301551104217439e-07, 
    8.4365700756473229e-07, 8.1522285834952874e-07, 7.8768473053256336e-07, 
    7.6102137002920793e-07, 7.3521596784180619e-07, 7.1025373516376354e-07, 
    6.8611986002098537e-07, 6.6279797206146037e-07, 6.40269184033174e-07, 
    6.1851171568153597e-07, 5.9750104339805982e-07, 5.7721046639670175e-07, 
    5.5761194232424641e-07, 5.3867702896716352e-07, 5.2037777467201262e-07, 
    5.0268742856437625e-07, 4.8558088652768286e-07, 4.6903484416825924e-07, 
    4.5302768291232159e-07, 4.3753916229109475e-07, 4.2255002118974169e-07, 
    4.0804160026669444e-07, 3.9399558462339717e-07, 3.8039393496064596e-07, 
    3.6721903187837339e-07, 3.5445401201062359e-07, 3.4208323348175293e-07, 
    3.3009278107904277e-07, 3.1847091142269352e-07, 3.0720834807170584e-07, 
    2.9629836167008391e-07, 2.857366068743174e-07, 2.7552072709829639e-07, 
    2.6564977407232716e-07, 2.5612351431489586e-07, 2.4694170645002152e-07, 
    2.3810342981855728e-07, 2.2960652948265185e-07, 2.2144721831566346e-07, 
    2.1361985023884247e-07, 2.0611685362231173e-07, 1.9892879586862492e-07, 
    1.9204454037621714e-07, 1.8545145676109931e-07, 1.7913565172548372e-07, 
    1.730821996695342e-07, 1.6727536446470262e-07, 1.6169881497144847e-07, 
    1.5633584347498928e-07, 1.5116959853541839e-07, 1.4618334069969574e-07, 
    1.4136072370422295e-07, 1.3668609578392048e-07, 1.3214480857695066e-07, 
    1.2772351540104038e-07, 1.2341043861400968e-07, 1.191955863871552e-07, 
    1.1507090343471742e-07, 1.1103034583534604e-07, 1.0706987706835675e-07, 
    1.0318738841691377e-07, 9.9382552139868499e-08, 9.5656618494614882e-08, 
    9.2012169162580028e-08, 8.8452838786308308e-08, 8.4983015279316899e-08, 
    8.1607527814809581e-08, 7.8331330883209467e-08, 7.5159192572605919e-08, 
    7.2095396709780965e-08, 6.9143469736905383e-08, 6.6305945199893751e-08, 
    6.3584178818018938e-08, 6.0978226491447197e-08, 5.8486794160488252e-08, 
    5.6107263747628954e-08, 5.3835792730360736e-08, 5.1667478309224527e-08, 
    4.9596570694718436e-08, 4.7616715908861072e-08, 4.5721206368539141e-08, 
    4.3903218926455226e-08, 4.2156023558702735e-08, 4.0473152071928016e-08, 
    3.8848522697423277e-08, 3.7276523302671673e-08, 3.5752060770539348e-08, 
    3.4270587339769195e-08, 3.2828114716638073e-08, 3.1421224991841871e-08, 
    3.004708333320074e-08, 2.8703452919355407e-08, 2.7388708018979015e-08, 
    2.6101838122664508e-08, 2.4842434492261477e-08, 2.3610651641108527e-08, 
    2.2407138780876472e-08, 2.1232940818465821e-08, 2.0089372947686403e-08, 
    1.8977877600031999e-08, 1.7899875503970844e-08, 1.6856624380402532e-08, 
    1.5849098130946661e-08, 1.4877897429480915e-08, 1.3943198731143959e-08, 
    1.304474469261922e-08, 1.2181874229822391e-08, 1.1353586831023517e-08, 
    1.0558632449157955e-08, 9.7956167875568535e-09, 9.0631108000942014e-09, 
    8.3597539717917674e-09, 7.6843418430006741e-09, 7.0358903351566491e-09, 
    6.4136714498872171e-09, 5.8172176319495376e-09, 5.2462945758843771e-09, 
    4.7008453727943148e-09, 4.1809114402119224e-09, 3.6865386664697801e-09, 
    3.2176791230935519e-09, 2.7741003748032574e-09, 2.3553143934306602e-09, 
    1.9605371053839282e-09, 1.5886865136194834e-09, 1.2384233237415807e-09, 
    9.0823238061276447e-10, 5.965376853873444e-10, 3.0183815327259244e-10, 
    2.2847434562311499e-11, -2.4138117117772279e-10, -4.9136289895822479e-10, 
    -7.2713808822404271e-10, -9.482866084818401e-10, -1.1540027420813475e-09, 
    -1.3432250190867914e-09, -1.5148085349998942e-09, 
    -1.6677212476441777e-09, -1.8012427314659744e-09, 
    -1.9151431382008069e-09, -2.0098226873792025e-09, 
    -2.0863965260772103e-09, -2.1467164460331395e-09, -2.1933276419436e-09, 
    -2.2293657995401807e-09, -2.2584050452199796e-09, 
    -2.2842714753712284e-09, -2.3108386303556469e-09, 
    -2.3418215680001704e-09, -2.3805843514021574e-09, 
    -2.4299733671923777e-09, -2.4921854396880679e-09, 
    -2.5686765938351226e-09, -2.6601140165915799e-09, 
    -2.7663713675937344e-09, -2.8865651594072488e-09, 
    -3.0191284496801876e-09, -3.1619163157762966e-09, 
    -3.3123365947831476e-09, -3.4674980528488556e-09, 
    -3.6243675149829511e-09, -3.7799267222835264e-09, 
    -3.9313199492365586e-09, -4.0759837385198839e-09, 
    -4.2117516390003402e-09, -4.3369285160678004e-09, -4.450331545932116e-09, 
    -4.5512974542474196e-09, -4.6396582754833195e-09, 
    -4.7156898611542967e-09, -4.7800392732626512e-09, 
    -4.8336378596944898e-09, -4.8776072808976828e-09, 
    -4.9131651171187141e-09, -4.9415360683127306e-09, 
    -4.9638733758988289e-09, -4.9811941350214763e-09, 
    -4.9943307368438134e-09, -5.0038999012998168e-09, 
    -5.0102895903075686e-09, -5.0136635264124367e-09, 
    -5.0139820108538962e-09, -5.0110371522514686e-09, 
    -5.0044996095028404e-09, -4.9939733308559144e-09, 
    -4.9790538898613135e-09, -4.9593857962923446e-09, 
    -4.9347138684904809e-09, -4.9049243633498156e-09, 
    -4.8700722441461965e-09, -4.8303925280797927e-09, 
    -4.7862950671558529e-09, -4.7383441127523652e-09, 
    -4.6872254412199749e-09, -4.6337052661334298e-09, 
    -4.5785856995729848e-09, -4.5226617558247055e-09, 
    -4.4666841065212593e-09, -4.4113308695735287e-09, 
    -4.3571899189610351e-09, -4.3047518297094976e-09, 
    -4.2544118947371132e-09, -4.2064786707174276e-09, 
    -4.1611857709485927e-09, -4.118703780485453e-09, -4.079149546501429e-09, 
    -4.0425912305683873e-09, -4.0090484881011676e-09, 
    -3.9784885735904618e-09, -3.9508198725445311e-09, 
    -3.9258852703572876e-09, -3.9034576660921426e-09, 
    -3.8832399277386237e-09, -3.8648706831811595e-09, 
    -3.8479366914355999e-09, -3.8319913424425691e-09, 
    -3.8165781795124046e-09, -3.8012573832034009e-09, 
    -3.7856329840813529e-09, -3.7693782699159477e-09, 
    -3.7522572093666652e-09, -3.7341399100456847e-09, 
    -3.7150108937079757e-09, -3.6949693663635457e-09, 
    -3.6742215226078828e-09, -3.6530652672088051e-09, 
    -3.6318685015119039e-09, -3.6110423934981709e-09, 
    -3.5910115421998726e-09, -3.5721830927181882e-09, 
    -3.5549171479099084e-09, -3.5395005837635867e-09, 
    -3.5261264430457187e-09, -3.5148804423906964e-09, 
    -3.5057358216008289e-09, -3.4985568023154888e-09, 
    -3.4931104241619092e-09, -3.4890854373427683e-09, 
    -3.4861165249518209e-09, -3.4838113670458277e-09, 
    -3.4817780251297116e-09, -3.479649955400783e-09, -3.4771065199485345e-09, 
    -3.473887226414707e-09, -3.4697989462666004e-09, -3.4647159751712561e-09, 
    -3.4585738268305047e-09, -3.4513581008190988e-09, 
    -3.4430904110036508e-09, -3.4338133114738615e-09, 
    -3.4235762631708994e-09, -3.4124241019074179e-09, 
    -3.4003892153910372e-09, -3.3874877771193881e-09, -3.37372008510622e-09, 
    -3.3590743151209296e-09, -3.3435329080265963e-09, 
    -3.3270804026946271e-09, -3.3097117702917081e-09, 
    -3.2914401654014173e-09, -3.2723034866912217e-09, 
    -3.2523691011080789e-09, -3.2317365613688836e-09, 
    -3.2105381019229205e-09, -3.1889370509023323e-09, 
    -3.1671241453948934e-09, -3.1453120501448592e-09, 
    -3.1237281626473349e-09, -3.1026061248695692e-09, 
    -3.0821762637279732e-09, -3.0626555348257249e-09, 
    -3.0442373889117041e-09, -3.0270823025486177e-09, 
    -3.0113094713423433e-09, -2.9969904061371356e-09, 
    -2.9841448161244822e-09, -2.9727392055478313e-09, 
    -2.9626882578481682e-09, -2.9538590125231729e-09, 
    -2.9460774417186766e-09, -2.9391371018514095e-09, 
    -2.9328091708935281e-09, -2.9268533746881077e-09, 
    -2.9210290578603565e-09, -2.9151059341958614e-09, 
    -2.9088738835923548e-09, -2.9021514587656495e-09, -2.894792632204553e-09, 
    -2.8866915887435697e-09, -2.8777852434489595e-09, 
    -2.8680534590866643e-09, -2.8575168119768028e-09, 
    -2.8462321081071069e-09, -2.8342857563134275e-09, 
    -2.8217854867933918e-09, -2.8088508167015716e-09, 
    -2.7956030207642569e-09, -2.7821552074578343e-09, -2.768603343648207e-09, 
    -2.7550188042382289e-09, -2.7414431200887762e-09, -2.727885181057233e-09, 
    -2.7143211681282096e-09, -2.7006970290765701e-09, 
    -2.6869333273917669e-09, -2.67293185180571e-09, -2.6585835232483032e-09, 
    -2.6437768320172581e-09, -2.6284062954074205e-09, 
    -2.6123802431933612e-09, -2.5956275839107143e-09, 
    -2.5781031224995473e-09, -2.5597913261532845e-09, 
    -2.5407083148772907e-09, -2.5209021901295455e-09, 
    -2.5004516459784825e-09, -2.4794630775367774e-09, 
    -2.4580662269020563e-09, -2.4364086990911587e-09, 
    -2.4146494947488655e-09, -2.3929519957540496e-09, 
    -2.3714767070608666e-09, -2.350374312103146e-09, -2.329779376507095e-09, 
    -2.309805283463607e-09, -2.2905406465753031e-09, -2.2720475412996282e-09, 
    -2.2543615412090848e-09, -2.2374935496074203e-09, 
    -2.2214330270692651e-09, -2.2061523070723469e-09, 
    -2.1916113649628487e-09, -2.1777625943418668e-09, 
    -2.1645550290035239e-09, -2.1519377341304841e-09, 
    -2.1398620397452872e-09, -2.1282827075918004e-09, 
    -2.1171580468379193e-09, -2.1064493345290008e-09, 
    -2.0961197628475752e-09, -2.0861333524067522e-09, 
    -2.0764540089505076e-09, -2.0670450124629403e-09, 
    -2.0578689249737719e-09, -2.0488879699906808e-09, 
    -2.0400646509957637e-09, -2.0313625173762422e-09, 
    -2.0227467663202322e-09, -2.014184632009737e-09, -2.0056453162646325e-09, 
    -1.9970995812565745e-09, -1.9885189597397053e-09, -1.979874836115778e-09, 
    -1.9711375284990558e-09, -1.9622756710619964e-09, 
    -1.9532560160586072e-09, -1.944043901698348e-09, -1.9346043470552342e-09, 
    -1.9249038577226494e-09, -1.9149127234115762e-09, 
    -1.9046077050942114e-09, -1.8939747852561157e-09, 
    -1.8830117792620761e-09, -1.871730453189538e-09, -1.860157991792993e-09, 
    -1.8483375160154064e-09, -1.8363276230511615e-09, 
    -1.8242007868908003e-09, -1.8120407217800722e-09, 
    -1.7999387356941496e-09, -1.7879893335509549e-09, 
    -1.7762852176342706e-09, -1.7649120836772438e-09, 
    -1.7539434766778826e-09, -1.743436174469382e-09, -1.7334263462607075e-09, 
    -1.7239269348501028e-09, -1.7149264188356347e-09, 
    -1.7063892194212579e-09, -1.6982576963673772e-09, 
    -1.6904557288021169e-09, -1.6828935686870387e-09, -1.675473684652281e-09, 
    -1.6680970761553736e-09, -1.6606696232515816e-09, 
    -1.6531078841724638e-09, -1.6453439687257344e-09, 
    -1.6373290099397791e-09, -1.6290350936014929e-09, 
    -1.6204554659871892e-09, -1.6116031593379028e-09, 
    -1.6025081750944989e-09, -1.5932136262615346e-09, 
    -1.5837711591117364e-09, -1.5742361806649058e-09, -1.564663229885293e-09, 
    -1.5551019532144567e-09, -1.5455938880945402e-09, 
    -1.5361703117055478e-09, -1.5268511628078829e-09, 
    -1.5176450708016005e-09, -1.5085502903614758e-09, 
    -1.4995564207414215e-09, -1.4906465977659136e-09, 
    -1.4817999708223237e-09, -1.4729941531725848e-09, 
    -1.4642074904550892e-09, -1.4554209189897752e-09, -1.446619371214188e-09, 
    -1.4377926018237005e-09, -1.4289355255507168e-09, 
    -1.4200480438774795e-09, -1.4111345400478789e-09, 
    -1.4022030712665523e-09, -1.3932644722495372e-09, 
    -1.3843313922349263e-09, -1.3754174289750386e-09, 
    -1.3665363513393857e-09, -1.3577015022528103e-09, 
    -1.3489253067197845e-09, -1.3402189155677412e-09, 
    -1.3315918962267277e-09, -1.3230520135010822e-09, 
    -1.3146049778479447e-09, -1.3062542623850035e-09, 
    -1.2980009288786639e-09, -1.2898435670733673e-09, 
    -1.2817783459942523e-09, -1.273799277976952e-09, -1.2658986601865424e-09, 
    -1.2580677958342488e-09, -1.2502978698218244e-09, 
    -1.2425810051551386e-09, -1.2349113491078086e-09, 
    -1.2272861409901447e-09, -1.2197065781996327e-09, 
    -1.2121784503794418e-09, -1.2047123928938283e-09, 
    -1.1973237570493193e-09, -1.1900320501053544e-09, 
    -1.1828600394092158e-09, -1.1758325094136676e-09, 
    -1.1689748535143435e-09, -1.162311548141332e-09, -1.1558646900698984e-09, 
    -1.1496526466298729e-09, -1.143688971128823e-09, -1.1379815801234123e-09, 
    -1.1325323071411366e-09, -1.1273367512329093e-09, 
    -1.1223844912129939e-09, -1.1176595370669336e-09, 
    -1.1131410503726718e-09, -1.1088041937779477e-09, 
    -1.1046211253754676e-09, -1.1005619982704514e-09, -1.096595998594127e-09, 
    -1.0926922959237559e-09, -1.0888209584549318e-09, 
    -1.0849537278757375e-09, -1.0810647274505464e-09, 
    -1.0771310285068354e-09, -1.0731331272777611e-09, 
    -1.0690553188371721e-09, -1.0648859991084668e-09, 
    -1.0606178688086399e-09, -1.0562481090085262e-09, 
    -1.0517784432722487e-09, -1.0472151808087174e-09, 
    -1.0425691242037092e-09, -1.037855415325852e-09, -1.0330932064030213e-09, 
    -1.0283052147187408e-09, -1.0235170522628649e-09, 
    -1.0187564005208192e-09, -1.0140519547814919e-09, 
    -1.0094322379771384e-09, -1.0049242466953775e-09, 
    -1.0005520662987509e-09, -9.9633548507550437e-10, 
    -9.9228874471091691e-10, -9.8841949204743703e-10, 
    -9.8472808136637612e-10, -9.8120723615845854e-10, 
    -9.7784222187701278e-10, -9.7461145746937854e-10, 
    -9.7148763483154181e-10, -9.684392162569046e-10, -9.6543229287611455e-10, 
    -9.6243259509152261e-10, -9.5940757881334e-10, -9.5632836415618747e-10, 
    -9.5317144356954132e-10, -9.4991994520011508e-10, 
    -9.4656442028713396e-10, -9.4310303665110188e-10, 
    -9.3954122648988962e-10, -9.3589075983465966e-10, 
    -9.3216839014383199e-10, -9.2839414582088638e-10, 
    -9.2458946715665807e-10, -9.2077529193190814e-10, 
    -9.1697030741531414e-10, -9.1318945246099866e-10, 
    -9.0944285073853393e-10, -9.0573515850539989e-10, 
    -9.0206546623901485e-10, -8.9842763949357046e-10, 
    -8.9481113055476926e-10, -8.9120211473716253e-10, 
    -8.8758490647267522e-10, -8.8394347181303504e-10, -8.802629639879777e-10, 
    -8.7653111264525676e-10, -8.7273942307783869e-10, 
    -8.6888401156771238e-10, -8.6496610715307708e-10, 
    -8.6099209564286664e-10, -8.5697318888197827e-10, 
    -8.5292466802936235e-10, -8.4886483335527743e-10, 
    -8.4481367592923013e-10, -8.4079144917912953e-10, 
    -8.3681718231437377e-10, -8.3290732310116663e-10, 
    -8.2907455638892066e-10, -8.2532695879316643e-10, 
    -8.2166748617553344e-10, -8.1809387869431053e-10, 
    -8.1459894350876801e-10, -8.1117122143389708e-10, 
    -8.0779591068707113e-10, -8.0445603407104293e-10, 
    -8.0113366176316481e-10, -7.9781117360605893e-10, 
    -7.9447238635605293e-10, -7.9110351555760042e-10, 
    -7.8769386745227117e-10, -7.8423629371640109e-10, 
    -7.8072730372062336e-10, -7.771669460452109e-10, -7.7355841263142533e-10, 
    -7.6990749042865633e-10, -7.6622184433808926e-10, 
    -7.6251025983542963e-10, -7.587818487297825e-10, -7.5504532714277927e-10, 
    -7.513083436274975e-10, -7.4757699917656268e-10, -7.4385546367578891e-10, 
    -7.4014583080205201e-10, -7.3644812628709624e-10, 
    -7.3276054732729955e-10, -7.2907985505216967e-10, 
    -7.2540194687575216e-10, -7.2172252084061798e-10, 
    -7.1803782412347389e-10, -7.1434536664379373e-10, 
    -7.1064458341415652e-10, -7.0693731629427666e-10, 
    -7.0322812169085939e-10, -6.9952429227887593e-10, 
    -6.9583563397705577e-10, -6.921739647458049e-10, -6.8855241223590368e-10, 
    -6.8498452884738468e-10, -6.8148336889210513e-10, 
    -6.7806053506777488e-10, -6.7472536051687716e-10, 
    -6.7148422587529682e-10, -6.6834012221264962e-10, 
    -6.6529242338564116e-10, -6.6233693199035763e-10, -6.59466109045147e-10, 
    -6.5666950758016745e-10, -6.5393431203505322e-10, 
    -6.5124599431050396e-10, -6.485889698930901e-10, -6.4594729457378565e-10, 
    -6.4330529243996602e-10, -6.4064818698056118e-10, -6.379626112130346e-10, 
    -6.3523710476758975e-10, -6.3246247724705937e-10, 
    -6.2963210940536862e-10, -6.2674214034284979e-10, 
    -6.2379157744309175e-10, -6.2078228419684479e-10, 
    -6.1771889655826254e-10, -6.1460863236724244e-10, -6.114610554738555e-10, 
    -6.0828774111924737e-10, -6.0510191590048428e-10, 
    -6.0191801230556811e-10, -5.9875122230590584e-10, 
    -5.9561696417175324e-10, -5.9253034974221353e-10, 
    -5.8950560941265239e-10, -5.8655553267951431e-10, 
    -5.8369093164301353e-10, -5.8092016608402299e-10, 
    -5.7824876244934404e-10, -5.756791979834237e-10, -5.732107821981604e-10, 
    -5.7083979105275603e-10, -5.685596935590571e-10, -5.6636157038258381e-10, 
    -5.6423460827112974e-10, -5.6216668091610618e-10, 
    -5.6014490994521856e-10, -5.5815621527394367e-10, 
    -5.5618775833797419e-10, -5.5422731719211671e-10, 
    -5.5226352533308433e-10, -5.5028604659747511e-10, 
    -5.4828563854740259e-10, -5.4625420500644691e-10, 
    -5.4418479831593674e-10, -5.4207165212997982e-10, 
    -5.3991020629571032e-10, -5.3769719783086593e-10, 
    -5.3543073350634099e-10, -5.3311040829679148e-10, 
    -5.3073737515258531e-10, -5.2831442606036363e-10, 
    -5.2584598076906133e-10, -5.2333801912790384e-10, 
    -5.2079792141111495e-10, -5.1823424046576973e-10, 
    -5.1565636443795383e-10, -5.1307414865429403e-10, 
    -5.1049747647864528e-10, -5.0793583836432839e-10, 
    -5.0539790119229812e-10, -5.0289117184072186e-10, 
    -5.0042171182238185e-10, -4.979939810914976e-10, -4.9561078704600239e-10, 
    -4.932733720133174e-10, -4.9098159291049996e-10, -4.8873421988979432e-10, 
    -4.8652928187510448e-10, -4.8436446898064137e-10, 
    -4.8223751705230818e-10, -4.8014659850490361e-10, 
    -4.7809063056888144e-10, -4.7606952875979701e-10, 
    -4.7408434713058854e-10, -4.7213733239276973e-10, 
    -4.7023183863555076e-10, -4.6837215376039395e-10, -4.6656319466124488e-10, 
    -4.6481013659508598e-10, -4.6311795601855049e-10, 
    -4.6149097338280904e-10, -4.5993239194333137e-10, 
    -4.5844392667420573e-10, -4.5702551700353484e-10, 
    -4.5567523161110161e-10, -4.5438930444666133e-10, 
    -4.5316238041056336e-10, -4.5198790247604704e-10, 
    -4.5085859130879185e-10, -4.4976698896312509e-10, -4.487059725485085e-10, 
    -4.4766915232456705e-10, -4.4665112441221326e-10, 
    -4.4564750533333172e-10, -4.4465477448110348e-10, 
    -4.4366990366514542e-10, -4.4268986635406506e-10, 
    -4.4171105230062378e-10, -4.4072870287116095e-10, 
    -4.3973642651951245e-10, -4.3872587906807867e-10, 
    -4.3768664149256996e-10, -4.3660634721561822e-10, -4.35471032473793e-10, 
    -4.3426572743266996e-10, -4.3297520663501257e-10, 
    -4.3158488334472316e-10, -4.3008177296200184e-10, 
    -4.2845547381761593e-10, -4.2669908600381696e-10, 
    -4.2481004208150471e-10, -4.2279074841730201e-10, 
    -4.2064902287711084e-10, -4.1839824207131639e-10, 
    -4.1605719015502187e-10, -4.1364954881058456e-10, 
    -4.1120305605276429e-10, -4.0874831308896365e-10, 
    -4.0631732349018127e-10, -4.0394180704588094e-10, 
    -4.0165143205777567e-10, -3.9947204628468049e-10, 
    -3.9742409017715653e-10, -3.9552128676331149e-10, 
    -3.9376975004964676e-10, -3.9216759177432099e-10, 
    -3.9070507928724886e-10, -3.8936533021277717e-10, 
    -3.8812553059967991e-10, -3.8695854333308807e-10, 
    -3.8583482932865816e-10, -3.8472448607045868e-10, 
    -3.8359926956929213e-10, -3.8243443534744109e-10, 
    -3.8121027106287754e-10, -3.7991319381277682e-10, 
    -3.7853636840149381e-10, -3.7707979808190831e-10, 
    -3.7554993550263912e-10, -3.7395883045784936e-10, 
    -3.7232296003778066e-10, -3.7066179491726893e-10, 
    -3.6899627283814121e-10, -3.6734726754305357e-10, -3.657341999084983e-10, 
    -3.6417384524864554e-10, -3.6267943488499025e-10, 
    -3.6126006169834858e-10, -3.5992041733863747e-10, 
    -3.5866082921046583e-10, -3.5747755723546151e-10, 
    -3.5636330442032706e-10, -3.5530788281437218e-10, -3.542989569563338e-10, 
    -3.5332285001044812e-10, -3.5236532325426272e-10, 
    -3.5141232847586344e-10, -3.5045068522167274e-10, 
    -3.4946869173247379e-10, -3.4845662595454421e-10, 
    -3.4740716236066072e-10, -3.46315669503114e-10, -3.4518040789444118e-10, 
    -3.4400261330195239e-10, -3.4278646893217952e-10, 
    -3.4153895737843097e-10, -3.4026963536696305e-10, 
    -3.3899028717791109e-10, -3.3771450628206514e-10, 
    -3.3645719768754156e-10, -3.3523402530603866e-10, 
    -3.3406080301522748e-10, -3.3295284852081774e-10, 
    -3.3192431088553127e-10, -3.3098748393650348e-10, 
    -3.3015212156171594e-10, -3.2942480126385842e-10, 
    -3.2880833370903008e-10, -3.2830130203171548e-10, 
    -3.2789773414091396e-10, -3.2758698526957575e-10, 
    -3.2735385079022353e-10, -3.2717893872482238e-10, 
    -3.2703931463170878e-10, -3.2690940286338937e-10, 
    -3.2676210368288919e-10, -3.2657006783803365e-10, 
    -3.2630705245824722e-10, -3.2594925762863889e-10, 
    -3.2547656248615107e-10, -3.2487356459885669e-10, 
    -3.2413035145928764e-10, -3.2324295220306727e-10, 
    -3.2221343070199923e-10, -3.2104965949847298e-10, 
    -3.1976475269678923e-10, -3.1837624063771395e-10, 
    -3.1690503913978068e-10, -3.1537428382002466e-10, 
    -3.1380811976857676e-10, -3.122304935588895e-10, -3.1066402728687205e-10, 
    -3.0912902796053142e-10, -3.0764265792044172e-10, 
    -3.0621830947981116e-10, -3.0486519106173536e-10, 
    -3.0358814255061159e-10, -3.0238767125424609e-10, 
    -3.0126021141993385e-10, -3.0019858330614774e-10, 
    -2.9919263496812778e-10, -2.9823003540345229e-10, 
    -2.9729715920453966e-10, -2.9638003282179389e-10, 
    -2.9546527183455672e-10, -2.9454093420979201e-10, 
    -2.9359726443657442e-10, -2.9262722856734351e-10, 
    -2.9162683252190613e-10, -2.9059519164519553e-10, 
    -2.8953435027945007e-10, -2.8844887120047353e-10, -2.873452588302743e-10, 
    -2.8623124907048638e-10, -2.8511505512837051e-10, 
    -2.8400463045478561e-10, -2.8290702158331341e-10, 
    -2.8182785239628106e-10, -2.8077096300346172e-10, 
    -2.7973822223794313e-10, -2.7872950356092933e-10, -2.777427798803814e-10, 
    -2.7677432281732503e-10, -2.7581896325087616e-10, -2.748703686920509e-10, 
    -2.7392134022536954e-10, -2.7296410425060837e-10, 
    -2.7199060253643307e-10, -2.7099279109256883e-10, 
    -2.6996296414378549e-10, -2.6889410911686806e-10, 
    -2.6778030068905212e-10, -2.6661711447604615e-10, 
    -2.6540204347577966e-10, -2.6413490531071512e-10, 
    -2.6281815916894369e-10, -2.6145711905149147e-10, 
    -2.6006001954677225e-10, -2.586378912341252e-10, -2.5720423571143338e-10, 
    -2.5577451283372987e-10, -2.5436543744462663e-10, 
    -2.5299414501930281e-10, -2.516772722536209e-10, -2.5043001097679119e-10, 
    -2.4926522232477934e-10, -2.481926553151893e-10, -2.4721833257019653e-10, 
    -2.4634417117967646e-10, -2.4556781729154894e-10, 
    -2.4488275110518974e-10, -2.4427861321276611e-10, 
    -2.4374175211158641e-10, -2.432559379537858e-10, -2.4280320415064706e-10, 
    -2.4236475165962979e-10, -2.4192189653745997e-10, 
    -2.4145697718787362e-10, -2.4095420610388798e-10, 
    -2.4040042082591743e-10, -2.397857188871135e-10, -2.3910392508899268e-10, 
    -2.3835291837186132e-10, -2.3753474793896341e-10, 
    -2.3665558209556969e-10, -2.3572543478614786e-10, 
    -2.3475771303434892e-10, -2.3376855527224916e-10, 
    -2.3277601102453309e-10, -2.3179906426683406e-10, 
    -2.3085658229423889e-10, -2.2996619774540637e-10, 
    -2.2914323991444438e-10, -2.2839973670522336e-10, 
    -2.2774360768915532e-10, -2.2717805945037982e-10, 
    -2.2670127635331571e-10, -2.2630639866301467e-10, 
    -2.2598183986852585e-10, -2.2571188103448718e-10, -2.254775491051882e-10, 
    -2.2525767668915804e-10, -2.2503011890290781e-10, 
    -2.2477299536268307e-10, -2.2446590908918678e-10, 
    -2.2409102870357514e-10, -2.2363399322208396e-10, 
    -2.2308454552469904e-10, -2.2243689713603561e-10, 
    -2.2168976036294499e-10, -2.2084610927162118e-10, 
    -2.1991264299369776e-10, -2.1889905493349462e-10, 
    -2.1781711669344031e-10, -2.1667972564670013e-10, 
    -2.1549991597634107e-10, -2.1428999898579066e-10, 
    -2.1306082308437398e-10, -2.118212809985474e-10, -2.1057803486301612e-10, 
    -2.0933552046797045e-10, -2.0809616722441276e-10, 
    -2.0686083102893764e-10, -2.0562933705797243e-10, 
    -2.0440111816765715e-10, -2.0317579944059649e-10, -2.019537305618858e-10, 
    -2.0073634759233844e-10, -1.9952638505364425e-10, 
    -1.9832786684597165e-10, -1.9714595093384962e-10, 
    -1.9598660445798906e-10, -1.9485620914136808e-10, 
    -1.9376109944775073e-10, -1.9270716748885555e-10, 
    -1.9169948904325806e-10, -1.9074210862772364e-10, 
    -1.8983791132798505e-10, -1.8898864619101052e-10, 
    -1.8819503754440688e-10, -1.8745700473082223e-10, 
    -1.8677388061302617e-10, -1.8614467758249756e-10, 
    -1.8556826747505657e-10, -1.8504354247769466e-10, 
    -1.8456945505644721e-10, -1.8414500406689773e-10, 
    -1.8376910569378548e-10, -1.8344044810721369e-10, 
    -1.8315725949323706e-10, -1.8291712294829635e-10, 
    -1.8271676370456162e-10, -1.8255193375149269e-10, 
    -1.8241732031151043e-10, -1.8230657922075045e-10, 
    -1.8221240412626132e-10, -1.8212671518152193e-10, 
    -1.8204086902365892e-10, -1.819459362128958e-10, -1.8183297170250823e-10, 
    -1.8169332266624212e-10, -1.8151887606164841e-10, 
    -1.8130235117030328e-10, -1.8103751033018716e-10, 
    -1.8071941064952285e-10, -1.8034460113136032e-10, 
    -1.7991136442369064e-10, -1.7941991037566252e-10, 
    -1.7887259899974743e-10, -1.7827408692810718e-10, 
    -1.7763146225731926e-10, -1.769542328426331e-10, -1.7625424789280697e-10, 
    -1.7554540743858126e-10, -1.7484324144955727e-10, 
    -1.7416428132434169e-10, -1.735253102308913e-10, -1.7294245183842998e-10, 
    -1.724302456760704e-10, -1.7200068809591142e-10, -1.7166239365130786e-10, 
    -1.714198835161422e-10, -1.7127314721318296e-10, -1.7121742862394308e-10, 
    -1.7124336270351366e-10, -1.7133737501273405e-10, 
    -1.7148238975658368e-10, -1.7165872703849127e-10, 
    -1.7184520555351064e-10, -1.7202027727147048e-10, 
    -1.7216318994823945e-10, -1.7225503432591996e-10, 
    -1.7227967677597153e-10, -1.7222443802264166e-10, 
    -1.7208057704441056e-10, -1.7184346942481282e-10, 
    -1.7151259729626511e-10, -1.7109126014145929e-10, 
    -1.7058614793442528e-10, -1.70006736115332e-10, -1.6936463424983421e-10, 
    -1.6867286151921953e-10, -1.6794515753800547e-10, 
    -1.6719529938516022e-10, -1.6643653467514942e-10, 
    -1.6568104698613827e-10, -1.6493955114577133e-10, 
    -1.6422094865109985e-10, -1.6353211186222915e-10, 
    -1.6287771775352287e-10, -1.6226022657479406e-10, 
    -1.6167991424150649e-10, -1.6113504046956689e-10, 
    -1.6062208891262103e-10, -1.6013615328949538e-10, 
    -1.5967136089165496e-10, -1.5922141120254664e-10, 
    -1.5878009625021735e-10, -1.5834186924338417e-10, 
    -1.5790230398213631e-10, -1.5745849499613705e-10, 
    -1.5700928254552582e-10, -1.5655535193726306e-10, 
    -1.5609911721994914e-10, -1.5564448409551806e-10, 
    -1.5519643074474435e-10, -1.5476053913891728e-10, 
    -1.5434243607773571e-10, -1.5394728055122631e-10, 
    -1.5357926511949607e-10, -1.5324126026345481e-10, 
    -1.5293453511345904e-10, -1.5265867097856391e-10, 
    -1.5241157937556154e-10, -1.521896920905374e-10, -1.519882391798947e-10, 
    -1.5180166384592914e-10, -1.5162404865962655e-10, -1.514496166981184e-10, 
    -1.5127315923245849e-10, -1.5109047602563056e-10, 
    -1.5089867406740675e-10, -1.506963731395106e-10, -1.504837490637658e-10, 
    -1.5026248106568363e-10, -1.5003550566794425e-10, 
    -1.4980669538683823e-10, -1.4958042075435633e-10, 
    -1.4936111268010995e-10, -1.4915279007161861e-10, 
    -1.4895867824263655e-10, -1.4878087766322474e-10, 
    -1.4862018673078402e-10, -1.4847600569104607e-10, 
    -1.4834641899865171e-10, -1.4822832473832612e-10, 
    -1.4811769334308159e-10, -1.480098355828288e-10, -1.478997242140862e-10, 
    -1.4778226403656179e-10, -1.4765257827463263e-10, 
    -1.4750620683864728e-10, -1.4733930023118058e-10, 
    -1.4714873293883327e-10, -1.4693222176154919e-10, -1.466883707594541e-10, 
    -1.4641673846364242e-10, -1.4611784462975967e-10, 
    -1.4579318716304886e-10, -1.4544518900977033e-10, 
    -1.4507715202815254e-10, -1.4469312167378863e-10, 
    -1.4429771891540529e-10, -1.4389589618037348e-10, 
    -1.4349267273742033e-10, -1.4309279244274165e-10, 
    -1.4270041272607372e-10, -1.4231876321993675e-10, 
    -1.4194989962493512e-10, -1.415944852961092e-10, -1.412517403086962e-10, 
    -1.4091947115181856e-10, -1.4059428600930359e-10, 
    -1.4027190438395683e-10, -1.3994762956760039e-10, 
    -1.3961686653899941e-10, -1.3927571147149674e-10, 
    -1.3892148195078876e-10, -1.3855322703045223e-10, 
    -1.3817204939130742e-10, -1.3778129255121789e-10, 
    -1.3738647740051752e-10, -1.3699506204182623e-10, 
    -1.3661593429486521e-10, -1.3625876926349348e-10, 
    -1.3593321044464543e-10, -1.3564803371686099e-10, 
    -1.3541027144846751e-10, -1.3522450400362123e-10, 
    -1.3509226501057212e-10, -1.3501172446830956e-10, 
    -1.3497760583054361e-10, -1.3498143714233698e-10, 
    -1.3501201765638012e-10, -1.3505615166260936e-10, -1.350994883513918e-10, 
    -1.3512746530885865e-10, -1.3512618763370672e-10, 
    -1.3508323401274647e-10, -1.3498823484815201e-10, 
    -1.3483327368372545e-10, -1.3461301088634828e-10, -1.343246078632305e-10, 
    -1.3396744523857416e-10, -1.3354276108198926e-10, 
    -1.3305320633993928e-10, -1.3250245566725704e-10, 
    -1.3189487371231238e-10, -1.3123533619386112e-10, 
    -1.3052913641240504e-10, -1.2978206701770813e-10, 
    -1.2900053589035493e-10, -1.2819174237805603e-10, 
    -1.2736379812884454e-10, -1.2652582294147245e-10, 
    -1.2568786589491206e-10, -1.2486073673806514e-10, 
    -1.2405566244611921e-10, -1.2328387860514028e-10, 
    -1.2255610233529259e-10, -1.2188201795613051e-10, 
    -1.2126975862433586e-10, -1.2072551221983258e-10, 
    -1.2025319971945196e-10, -1.1985433505814905e-10, 
    -1.1952800586607987e-10, -1.1927103971223459e-10, 
    -1.1907825525104957e-10, -1.1894284524671821e-10, 
    -1.1885679021433592e-10, -1.1881131201511234e-10, 
    -1.1879727123908852e-10, -1.1880555152086715e-10, 
    -1.1882730665417307e-10, -1.1885415304389346e-10, 
    -1.1887821292549409e-10, -1.1889210203505325e-10, 
    -1.1888880816564783e-10, -1.188615689344809e-10, -1.1880371286663376e-10, 
    -1.1870859328539352e-10, -1.185695649157924e-10, -1.1838009872673292e-10, 
    -1.1813398893255002e-10, -1.1782571169282077e-10, -1.174508203727274e-10, 
    -1.1700642399141386e-10, -1.1649160489400962e-10, 
    -1.1590781443866187e-10, -1.1525909649222537e-10, 
    -1.1455218792002216e-10, -1.1379640339961598e-10, 
    -1.1300337039672124e-10, -1.1218657020030636e-10, 
    -1.1136078129526237e-10, -1.1054142211633227e-10, 
    -1.0974389322804056e-10, -1.0898291115447677e-10, 
    -1.0827193894602095e-10, -1.076226741322344e-10, -1.0704468624346306e-10, 
    -1.0654512839464924e-10, -1.0612861276278142e-10, 
    -1.0579715381012064e-10, -1.0555024635969999e-10, 
    -1.0538499946893969e-10, -1.0529639487306883e-10, 
    -1.0527756945932499e-10, -1.0532018355791429e-10, 
    -1.0541480347992635e-10, -1.0555133163585786e-10, 
    -1.0571940088774485e-10, -1.0590877171938274e-10, 
    -1.0610965586505645e-10, -1.0631300250169813e-10, -1.065106741843272e-10, 
    -1.0669559329376715e-10, -1.0686178510526915e-10, 
    -1.0700438264037755e-10, -1.0711959453645355e-10, 
    -1.0720466891064389e-10, -1.0725783713189212e-10, 
    -1.0727828599524059e-10, -1.0726612020026136e-10, 
    -1.0722233617978874e-10, -1.0714875930102906e-10, 
    -1.0704797260403669e-10, -1.0692316428247328e-10, 
    -1.0677794084292525e-10, -1.0661605497860528e-10, 
    -1.0644110146144302e-10, -1.0625616192944755e-10, 
    -1.0606347869001147e-10, -1.0586412315669128e-10, 
    -1.0565776452201267e-10, -1.0544251894258884e-10, 
    -1.0521492494853459e-10, -1.0497004207049277e-10, -1.047017008380057e-10, 
    -1.0440285045412448e-10, -1.040660169069308e-10, -1.0368381333964524e-10, 
    -1.0324948421354416e-10, -1.0275742633487351e-10, 
    -1.0220365891125703e-10, -1.0158618640499985e-10, 
    -1.0090525701411342e-10, -1.0016345929583941e-10, -9.93656776457636e-11, 
    -9.8518877910153591e-11, -9.7631775474270273e-11, 
    -9.6714376052014384e-11, -9.5777433553645027e-11, 
    -9.4831871766344566e-11, -9.3888216089980671e-11, 
    -9.2956051776403636e-11, -9.2043580730489802e-11, 
    -9.1157273438147031e-11, -9.0301674435437889e-11, 
    -8.9479331005429903e-11, -8.8690883411027564e-11, 
    -8.7935279732442122e-11, -8.7210119895028383e-11, 
    -8.6512084399478173e-11, -8.5837426517399662e-11, 
    -8.5182494592296282e-11, -8.4544248137545101e-11, 
    -8.3920716166106959e-11, -8.3311394896579151e-11, 
    -8.2717510173616018e-11, -8.2142149898234917e-11, 
    -8.1590232414559999e-11, -8.1068314302529477e-11, 
    -8.0584225473463872e-11, -8.014657203638124e-11, -7.9764128441009362e-11, 
    -7.9445156675693291e-11, -7.9196730717876263e-11, 
    -7.9024105677551046e-11, -7.89301988274856e-11, -7.8915236292402492e-11, 
    -7.89765935243269e-11, -7.910886101802793e-11, -7.9304123522273744e-11, 
    -7.9552439609784163e-11, -7.984246944122662e-11, -8.0162197512034679e-11, 
    -8.0499688133995705e-11, -8.0843782829251215e-11, 
    -8.1184704242001665e-11, -8.1514497450191965e-11, 
    -8.1827284156879882e-11, -8.2119304248249279e-11, 
    -8.2388773608365655e-11, -8.2635588251094007e-11, 
    -8.2860901149301107e-11, -8.3066642699489314e-11, 
    -8.3255041482821645e-11, -8.3428191247640749e-11, 
    -8.3587711155642119e-11, -8.3734518756243259e-11, 
    -8.3868735870493034e-11, -8.3989718794096817e-11, 
    -8.4096191279412089e-11, -8.4186452785979744e-11, 
    -8.4258633632067726e-11, -8.4310961838338306e-11, 
    -8.4342012679749576e-11, -8.4350920859233059e-11, 
    -8.4337535965188248e-11, -8.4302534931555243e-11, 
    -8.4247464129879457e-11, -8.4174738014259069e-11, 
    -8.4087604816329532e-11, -8.399005751735687e-11, -8.388673214280483e-11, 
    -8.3782786088060174e-11, -8.3683742835517925e-11, 
    -8.3595322963568054e-11, -8.3523259767445804e-11, 
    -8.3473089354802157e-11, -8.3449930281192105e-11, 
    -8.3458259669026586e-11, -8.3501676206457102e-11, 
    -8.3582685932347816e-11, -8.3702496193328057e-11, 
    -8.3860846198284181e-11, -8.405588519482788e-11, -8.4284101787173519e-11, 
    -8.4540323510714944e-11, -8.4817793823785692e-11, 
    -8.5108318069285335e-11, -8.5402509310296558e-11, 
    -8.5690093450317112e-11, -8.5960282251873395e-11, 
    -8.6202186258243556e-11, -8.6405270170522403e-11, 
    -8.6559789755366069e-11, -8.665719453778943e-11, -8.6690490151498683e-11, 
    -8.6654499806506266e-11, -8.6546037405204874e-11, 
    -8.6363994093986993e-11, -8.6109295482578333e-11, 
    -8.5784796838283628e-11, -8.5395101669199216e-11, 
    -8.4946335815050757e-11, -8.4445901490512141e-11, 
    -8.3902240448892103e-11, -8.3324606203493022e-11, 
    -8.2722847165403586e-11, -8.2107206653841662e-11, 
    -8.1488147797980676e-11, -8.0876145348863799e-11, 
    -8.0281470978429374e-11, -7.9713946877873709e-11, 
    -7.9182683332443742e-11, -7.8695793673922119e-11, 
    -7.8260127754044197e-11, -7.7881034045539481e-11, 
    -7.7562203362105112e-11, -7.7305598986240731e-11, 
    -7.7111509247718303e-11, -7.6978716272876774e-11, 
    -7.6904780728077015e-11, -7.688640349586296e-11, -7.6919829013855239e-11, 
    -7.7001238646116679e-11, -7.7127088801464661e-11, 
    -7.7294333290270213e-11, -7.7500527388076648e-11, 
    -7.7743764761237047e-11, -7.8022498677654133e-11, 
    -7.8335244688617319e-11, -7.8680228666745478e-11, 
    -7.9055028078271457e-11, -7.9456283321816242e-11, 
    -7.9879487449101526e-11, -8.0318954293135714e-11, 
    -8.0767903594741161e-11, -8.1218724934132059e-11, -8.166335591495034e-11, 
    -8.2093731769794867e-11, -8.2502259006687941e-11, 
    -8.2882276546105297e-11, -8.3228403891390968e-11, -8.353678659850954e-11, 
    -8.3805171326527883e-11, -8.4032860487397089e-11, 
    -8.4220484835315213e-11, -8.4369708404762546e-11, 
    -8.4482833961400389e-11, -8.4562400127083654e-11, 
    -8.4610793859939722e-11, -8.4629941569428453e-11, 
    -8.4621070150032467e-11, -8.4584617324160763e-11, 
    -8.4520222236189683e-11, -8.4426850453624223e-11, 
    -8.4302988093309969e-11, -8.4146896816083526e-11, 
    -8.3956880647962623e-11, -8.3731547206303833e-11, 
    -8.3469991697556834e-11, -8.3171935041391156e-11, 
    -8.2837734433609995e-11, -8.246833333474844e-11, -8.2065098054644477e-11, 
    -8.1629619109783398e-11, -8.1163458555606929e-11, 
    -8.0667937264282677e-11, -8.0143938321474535e-11, 
    -7.9591820833167136e-11, -7.9011410102094993e-11, 
    -7.8402125282754594e-11, -7.7763190161453562e-11, 
    -7.7093958788294774e-11, -7.6394262700002238e-11, -7.5664800523723e-11, 
    -7.4907458792435792e-11, -7.4125587211825444e-11, 
    -7.3324132917993973e-11, -7.2509658560381558e-11, 
    -7.1690196191265054e-11, -7.0874992015269789e-11, 
    -7.0074117937409811e-11, -6.9298005328901721e-11, 
    -6.8556931257867868e-11, -6.7860526046952612e-11, 
    -6.7217288158864379e-11, -6.6634190286375598e-11, 
    -6.6116360461886661e-11, -6.5666899902763496e-11, 
    -6.5286786011828173e-11, -6.4974922843752111e-11, 
    -6.4728270486001298e-11, -6.4542094659425035e-11, 
    -6.4410265354572667e-11, -6.4325633476363704e-11, 
    -6.4280415819766926e-11, -6.4266595019209157e-11, 
    -6.4276292860418928e-11, -6.4302103244830849e-11, 
    -6.4337344428772469e-11, -6.4376258500143371e-11, 
    -6.4414095283554973e-11, -6.4447134513456941e-11, 
    -6.4472609679035523e-11, -6.4488584550015122e-11, 
    -6.4493775884468198e-11, -6.4487365268930478e-11, 
    -6.4468800158409834e-11, -6.4437638654458288e-11, 
    -6.4393405379265805e-11, -6.4335530769141691e-11, 
    -6.4263315364324528e-11, -6.4175961751804651e-11, 
    -6.4072647511235618e-11, -6.3952653562039237e-11, 
    -6.3815498521681918e-11, -6.3661127773527094e-11, 
    -6.3490077844749015e-11, -6.3303671210619348e-11, 
    -6.3104172196668819e-11, -6.2894937580637611e-11, 
    -6.2680508189028987e-11, -6.246664725769353e-11, -6.2260302445601e-11, 
    -6.2069479045819681e-11, -6.1903008669082919e-11, 
    -6.1770229533565519e-11, -6.1680564173789228e-11, 
    -6.1643034987138292e-11, -6.1665728099442808e-11, -6.175527172332543e-11, 
    -6.1916349658150749e-11, -6.215130189125173e-11, -6.2459856880481796e-11, 
    -6.2839053415004296e-11, -6.3283316227340447e-11, 
    -6.3784741730252831e-11, -6.433354767901483e-11, -6.4918658232931341e-11, 
    -6.5528382693589575e-11, -6.6151123316413833e-11, 
    -6.6776044181549089e-11, -6.7393662156850162e-11, 
    -6.7996273324920614e-11, -6.8578226030356179e-11, 
    -6.9135979671494964e-11, -6.9667979390969741e-11, 
    -7.0174364276340881e-11, -7.0656536750918045e-11, -7.111665550521772e-11, 
    -7.155712153363945e-11, -7.1980075917957188e-11, -7.2387001413225574e-11, 
    -7.2778428352591181e-11, -7.3153804936609382e-11, 
    -7.3511491772589175e-11, -7.3848906660211657e-11, 
    -7.4162782865618464e-11, -7.4449471741151487e-11, 
    -7.4705295870864781e-11, -7.4926884800216015e-11, 
    -7.5111447961402998e-11, -7.525696204295055e-11, -7.5362260116532207e-11, 
    -7.5427011312391277e-11, -7.5451591749792311e-11, 
    -7.5436884506498597e-11, -7.5384022207739545e-11, 
    -7.5294105023138262e-11, -7.5167950264105305e-11, 
    -7.5005884460956397e-11, -7.4807625476957967e-11, 
    -7.4572255903048905e-11, -7.4298320904997219e-11, 
    -7.3984017574703878e-11, -7.3627479748120752e-11, 
    -7.3227150589926858e-11, -7.2782168639150262e-11, 
    -7.2292766243100599e-11, -7.1760628156875107e-11, 
    -7.1189178302924842e-11, -7.0583759421442068e-11, 
    -6.9951683276921506e-11, -6.9302138356284502e-11, 
    -6.8645942563572058e-11, -6.7995160109123135e-11, 
    -6.7362601123186628e-11, -6.6761213197996995e-11, 
    -6.6203441539426751e-11, -6.5700571396353404e-11, 
    -6.5262092182799854e-11, -6.4895167122158006e-11, 
    -6.4604200601793951e-11, -6.4390557461996245e-11, 
    -6.4252447147126746e-11, -6.4184969516589826e-11, 
    -6.4180320115865963e-11, -6.4228140172992514e-11, 
    -6.4315997175448847e-11, -6.4429954863417421e-11, 
    -6.4555203527922472e-11, -6.4676740098928393e-11, 
    -6.4780060274071953e-11, -6.485182843278172e-11, -6.4880510407199079e-11, 
    -6.4856934326851912e-11, -6.4774744664685787e-11, 
    -6.4630731975766164e-11, -6.4425004374162822e-11, 
    -6.4160985321989535e-11, -6.38452153746841e-11, -6.3486975231046651e-11, 
    -6.3097731766197713e-11, -6.2690450635872122e-11, 
    -6.2278808216371333e-11, -6.187637029048043e-11, -6.1495786913591032e-11, 
    -6.1148069496442222e-11, -6.0841994637667919e-11, 
    -6.0583681581181323e-11, -6.0376364868389339e-11, 
    -6.0220361395578017e-11, -6.0113232699018054e-11, 
    -6.0050112513693871e-11, -6.0024162881342695e-11, 
    -6.0027122968306871e-11, -6.0049895667027227e-11, 
    -6.0083142093760527e-11, -6.0117832824901934e-11, 
    -6.0145735149056428e-11, -6.0159795378419175e-11, 
    -6.0154416741163054e-11, -6.0125621019613269e-11, 
    -6.0071101459411823e-11, -5.9990151302806066e-11, 
    -5.9883529116034537e-11, -5.9753238249407436e-11, 
    -5.9602270793806729e-11, -5.9434333060307072e-11, 
    -5.9253565700600574e-11, -5.9064280483695611e-11, 
    -5.8870737523330127e-11, -5.867694691019017e-11, -5.8486523857164668e-11, 
    -5.8302577520788186e-11, -5.8127641054848368e-11, 
    -5.7963645346785103e-11, -5.7811927114432702e-11, 
    -5.7673256245293546e-11, -5.7547916944826256e-11, -5.743580348938573e-11, 
    -5.733655531656555e-11, -5.7249691424033505e-11, -5.7174762233689829e-11, 
    -5.7111506985805194e-11, -5.7059979577407819e-11, -5.702064185333898e-11, 
    -5.699443156715399e-11, -5.6982766570424501e-11, -5.6987515451770354e-11, 
    -5.7010918648218335e-11, -5.7055478189219757e-11, -5.712382873652508e-11, 
    -5.7218604374061709e-11, -5.7342288381723408e-11, 
    -5.7497093412801089e-11, -5.7684851332147121e-11, 
    -5.7906925220047503e-11, -5.8164124400660916e-11, 
    -5.8456653868116422e-11, -5.878407567717903e-11, -5.9145290927300388e-11, 
    -5.9538519674789077e-11, -5.9961321243726117e-11, 
    -6.0410615250535017e-11, -6.0882715632404663e-11, 
    -6.1373375911643088e-11, -6.1877838225584977e-11, 
    -6.2390868816700248e-11, -6.2906794460928305e-11, 
    -6.3419526548446877e-11, -6.3922582862172344e-11, 
    -6.4409099932487093e-11, -6.4871871789258846e-11, -6.530340829354559e-11, 
    -6.5696040088598687e-11, -6.6042065731458983e-11, 
    -6.6333962470011939e-11, -6.6564640201187648e-11, 
    -6.6727732869784364e-11, -6.681790264572792e-11, -6.6831144432985641e-11, 
    -6.6765025328780354e-11, -6.661888442371819e-11, -6.6393924497157242e-11, 
    -6.6093211452041681e-11, -6.5721573868688914e-11, 
    -6.5285400905007059e-11, -6.4792361725945689e-11, 
    -6.4251083588220331e-11, -6.3670788788825799e-11, 
    -6.3060952098217882e-11, -6.2430976853982084e-11, 
    -6.1789931858614891e-11, -6.1146336771951425e-11, 
    -6.0508036350738109e-11, -5.9882110428897717e-11, -5.927485456533848e-11, 
    -5.8691798425087171e-11, -5.8137735257369638e-11, 
    -5.7616776648178118e-11, -5.7132400462657843e-11, -5.668749446011585e-11, 
    -5.6284413417692269e-11, -5.5925026957323464e-11, -5.561078929763309e-11, 
    -5.5342830757841136e-11, -5.5122073703142295e-11, 
    -5.4949353667484984e-11, -5.4825569072529549e-11, 
    -5.4751801634540456e-11, -5.4729411639563684e-11, 
    -5.4760070523441225e-11, -5.4845709627064182e-11, 
    -5.4988365585417926e-11, -5.5189928628360944e-11, 
    -5.5451791876185545e-11, -5.5774436606143174e-11, 
    -5.6156979102258773e-11, -5.6596742868501842e-11, 
    -5.7088912423779199e-11, -5.7626307926746365e-11, 
    -5.8199336632674851e-11, -5.879615860945278e-11, -5.9403065778391098e-11, 
    -6.0005074574366411e-11, -6.0586680506596495e-11, 
    -6.1132736720903868e-11, -6.1629350902574375e-11, 
    -6.2064751898560134e-11, -6.243001007104033e-11, -6.271955497077735e-11, 
    -6.293142032534204e-11, -6.3067205810933561e-11, -6.3131726938982648e-11, 
    -6.3132412700865663e-11, -6.3078499645940335e-11, 
    -6.2980101473378842e-11, -6.2847255176234041e-11, 
    -6.2689042122183154e-11, -6.2512861946813162e-11, -6.23239473393766e-11, 
    -6.2125133005430878e-11, -6.1916919272331797e-11, -6.169778754417466e-11, 
    -6.1464735280714895e-11, -6.1213950262126693e-11, 
    -6.0941553765062512e-11, -6.0644326874776132e-11, 
    -6.0320353612462176e-11, -5.9969503668350113e-11, 
    -5.9593755520348033e-11, -5.9197287867024278e-11, 
    -5.8786399869309988e-11, -5.8369247647912802e-11, 
    -5.7955447459254665e-11, -5.7555576788036356e-11, 
    -5.7180631437699189e-11, -5.6841466214273196e-11, -5.654826198971764e-11, 
    -5.6310045911673995e-11, -5.613427807612428e-11, -5.6026524573998265e-11, 
    -5.5990220076141371e-11,
  // Sqw-F(6, 0-1999)
    0.026152068924167011, 0.026147953913105718, 0.02613560876565215, 
    0.026115031694899263, 0.026086215183419151, 0.026049140090693892, 
    0.026003769084629577, 0.025950040750577687, 0.025887865711692139, 
    0.025817125866854369, 0.025737677456958107, 0.025649358173829882, 
    0.025551998009821591, 0.02544543309157796, 0.025329521415786573, 
    0.025204159249012884, 0.025069296976511567, 0.024924953361543097, 
    0.024771227455390583, 0.024608307711159905, 0.024436478132122789, 
    0.024256121471448941, 0.02406771956335696, 0.023871850806676385, 
    0.023669184673509602, 0.023460472936786863, 0.023246537173149191, 
    0.023028252071771456, 0.022806524217377722, 0.022582266337676998, 
    0.022356367494100828, 0.02212966029380779, 0.021902886822943914, 
    0.02167666554139942, 0.021451461733736393, 0.021227564195133893, 
    0.021005070596518089, 0.020783883417500287, 0.020563717506920907, 
    0.020344119320443787, 0.020124496815665222, 0.019904157992968491, 
    0.019682355281762067, 0.019458332485360861, 0.019231370868684546, 
    0.019000831204840623, 0.018766189142495133, 0.018527062027056704, 
    0.018283226190625678, 0.018034624597619547, 0.01778136548764252, 
    0.01752371321695927, 0.017262072827127897, 0.0169969699683486, 
    0.016729027716755655, 0.016458941614685082, 0.016187454005282546, 
    0.015915328495186065, 0.01564332520897211, 0.01537217741663289, 
    0.015102570111887276, 0.014835121162606515, 0.014570365699554957, 
    0.014308744409360511, 0.014050596315998186, 0.013796156455181396, 
    0.013545558574145774, 0.013298842653456856, 0.01305596669157234, 
    0.012816821867529905, 0.012581249949453893, 0.012349061681267112, 
    0.012120054873252416, 0.011894031039510441, 0.01167080964389453, 
    0.011450239299506799, 0.011232205573449732, 0.011016635338626866, 
    0.010803497857211903, 0.01059280295829524, 0.010384596781657814, 
    0.010178955609307322, 0.0099759783129450309, 0.0097757779279778346, 
    0.0095784728393406206, 0.0093841780409528366, 0.0091929969106333033, 
    0.0090050139199854638, 0.0088202886640203204, 0.0086388515377108666, 
    0.0084607012996443, 0.0082858046465480503, 0.008114097784505921, 
    0.0079454898374973805, 0.0077798677993758366, 0.0076171026290051125, 
    0.0074570560230921889, 0.0072995873832474951, 0.0071445605208161744, 
    0.0069918497058472596, 0.0068413447516289276, 0.0066929549191328324, 
    0.0065466115146545949, 0.0064022691319734005, 0.0062599055560590665, 
    0.0061195204017777749, 0.0059811326132917222, 0.005844777002196563, 
    0.0057105000558372978, 0.0055783552980096102, 0.0054483985243902293, 
    0.0053206832541503072, 0.0051952567274605108, 0.0050721567299957682, 
    0.0049514094404851678, 0.0048330283838086494, 0.0047170144449912412, 
    0.0046033567780389088, 0.0044920343479652319, 0.0043830177912065017, 
    0.0042762712784014034, 0.0041717541142824634, 0.0040694219024294256, 
    0.0039692272200038126, 0.00387111986677157, 0.003775046850986531, 
    0.0036809523336617106, 0.0035887777620465036, 0.0034984623824325344, 
    0.0034099442413667823, 0.0033231616803859384, 0.0032380552240016125, 
    0.0031545696748879288, 0.0030726561803075701, 0.0029922740280188698, 
    0.0029133919671163709, 0.002835988919604111, 0.0027600540359061696, 
    0.0026855861334585808, 0.0026125926252050249, 0.0025410880827626274, 
    0.0024710925833485459, 0.0024026299643808303, 0.002335726065703717, 
    0.0022704069910480821, 0.0022066973821111835, 0.0021446186815679905, 
    0.0020841873704414496, 0.0020254131984864072, 0.0019682974750212644, 
    0.0019128315390218411, 0.0018589955670045518, 0.001806757892967087, 
    0.0017560749988803001, 0.0017068922858105042, 0.0016591456602637533, 
    0.0016127638788778435, 0.0015676715015544951, 0.0015237922234388249, 
    0.0014810523025131858, 0.0014393837802678946, 0.0013987272106357567, 
    0.0013590336640867131, 0.0013202658515898541, 0.0012823983059368916, 
    0.0012454166532946814, 0.0012093160940877421, 0.0011740992799400343, 
    0.0011397738162465748, 0.0011063496355239891, 0.0010738364760477998, 
    0.0010422416673827491, 0.0010115683752152291, 0.00098181439939551136, 
    0.00095297155834915895, 0.00092502563637256294, 0.00089795682284303784, 
    0.00087174053749499759, 0.00084634851535358155, 0.000821750018762787, 
    0.00079791305088204047, 0.00077480546269129505, 0.00075239587090193314, 
    0.00073065433390488862, 0.00070955276373815433, 0.00068906508111012154, 
    0.00066916714538622912, 0.00064983651040199377, 0.00063105206895245779, 
    0.0006127936534486056, 0.0005950416577562319, 0.00057777673641692983, 
    0.00056097962351238037, 0.0005446310959498446, 0.0005287120867326525, 
    0.00051320393477319206, 0.0004980887409101409, 0.00048334978672108704, 
    0.00046897196481841098, 0.00045494216740223623, 0.0004412495840874338, 
    0.00042788586989387159, 0.00041484515858267943, 0.00040212391349014166, 
    0.00038972062556964446, 0.00037763538436429519, 0.0003658693601915901, 
    0.00035442424352803936, 0.00034330168972158053, 0.00033250281379823549, 
    0.00032202777205496733, 0.00031187545571170885, 0.00030204330882824829, 
    0.00029252726973518281, 0.00028332182392913668, 0.00027442014788067086, 
    0.00026581431810535148, 0.00025749555822257201, 0.00024945449816637748, 
    0.00024168142348880429, 0.0002341664979151596, 0.0002268999480899336, 
    0.00021987220503891485, 0.00021307400173284279, 0.00020649642996438026, 
    0.0002001309624511678, 0.00019396944770760021, 0.00018800408593203359, 
    0.00018222739410036768, 0.00017663216779922539, 0.00017121144619575336, 
    0.00016595848503361485, 0.00016086674076570438, 0.00015592986700925586, 
    0.00015114172259390426, 0.00014649638876261382, 0.0001419881917833972, 
    0.00013761172652545901, 0.00013336187656989184, 0.00012923382718996729, 
    0.00012522306894913532, 0.00012132539150664172, 0.00011753686916997137, 
    0.00011385384142761938, 0.00011027289278959099, 0.00010679083650763857, 
    0.00010340470603836739, 0.00010011175653105073, 9.6909476421517515e-05, 
    9.3795606787007595e-05, 9.0768163918117885e-05, 8.7825459028216052e-05, 
    8.4966108471312742e-05, 8.2189028429684451e-05, 7.9493409706102208e-05, 
    7.6878670763826418e-05, 7.4344390097648281e-05, 7.1890221920039004e-05, 
    6.9515801546868674e-05, 6.7220648406541279e-05, 6.5004075067206591e-05, 
    6.286511005815408e-05, 6.0802440703789195e-05, 5.8814379980657721e-05, 
    5.6898858907643674e-05, 5.5053443555064602e-05, 5.3275373717450128e-05, 
    5.1561618849555371e-05, 4.9908946103297713e-05, 4.8313995199196662e-05, 
    4.6773355296919518e-05, 4.5283639819009982e-05, 4.3841556132489028e-05, 
    4.2443967929843495e-05, 4.1087948941153996e-05, 3.9770827183740422e-05, 
    3.8490219302058161e-05, 3.7244054711632981e-05, 3.6030589308909945e-05, 
    3.4848408534324265e-05, 3.3696419658203144e-05, 3.2573833359896412e-05, 
    3.1480135014021051e-05, 3.0415046576278068e-05, 2.9378480528791456e-05, 
    2.8370487934701498e-05, 2.7391203178896107e-05, 2.644078835678011e-05, 
    2.5519380445359058e-05, 2.4627044309287623e-05, 2.3763734244456393e-05, 
    2.2929266166113313e-05, 2.2123301756681601e-05, 2.1345344976714573e-05, 
    2.0594750396852247e-05, 1.9870741921413436e-05, 1.9172439726369705e-05, 
    1.8498892693283916e-05, 1.7849113328667829e-05, 1.7222112134714144e-05, 
    1.661692863362548e-05, 1.603265671528018e-05, 1.5468462625353582e-05, 
    1.4923594676889079e-05, 1.439738457933135e-05, 1.388924106368543e-05, 
    1.3398637169167035e-05, 1.2925093087188318e-05, 1.2468156785385701e-05, 
    1.2027384732404284e-05, 1.1602324906259657e-05, 1.1192503914319357e-05, 
    1.079741951865732e-05, 1.041653920620467e-05, 1.004930473780249e-05, 
    9.6951419323491637e-06, 9.3534743641881142e-06, 9.0237392379282715e-06, 
    8.7054034974685939e-06, 8.3979782460005243e-06, 8.1010297919788264e-06, 
    7.8141860606092974e-06, 7.537137664510248e-06, 7.2696335435150164e-06, 
    7.0114716863784811e-06, 6.7624859688770831e-06, 6.5225305260003962e-06, 
    6.2914632859959341e-06, 6.0691303161245972e-06, 5.8553524753295809e-06, 
    5.6499155652397827e-06, 5.4525647632613625e-06, 5.2630036596920362e-06, 
    5.0808977585164915e-06, 4.9058818845530624e-06, 4.7375706069446565e-06, 
    4.5755705646292508e-06, 4.419493476864538e-06, 4.2689686390551626e-06, 
    4.1236538308825647e-06, 3.983243777898442e-06, 3.8474755846870093e-06, 
    3.7161308660321176e-06, 3.5890346139937953e-06, 3.4660511238192591e-06, 
    3.3470775381961594e-06, 3.2320357381786452e-06, 3.1208634011608462e-06, 
    3.0135050569325775e-06, 2.9099039081384895e-06, 2.8099950509774725e-06, 
    2.7137005535003302e-06, 2.6209266412020548e-06, 2.5315630253347653e-06, 
    2.4454842082267122e-06, 2.3625524314594404e-06, 2.2826218096720145e-06, 
    2.205543125116727e-06, 2.1311687467593989e-06, 2.0593571808881304e-06, 
    1.9899768473280084e-06, 1.9229087951833234e-06, 1.8580482077688085e-06, 
    1.7953046837309044e-06, 1.7346014043627309e-06, 1.6758733956841787e-06, 
    1.6190651587502943e-06, 1.5641279709365404e-06, 1.5110171544875655e-06, 
    1.4596895723133182e-06, 1.4101015514933777e-06, 1.362207362722837e-06, 
    1.3159583077247693e-06, 1.2713023969056851e-06, 1.2281845423878549e-06, 
    1.1865471535617326e-06, 1.1463310041090379e-06, 1.1074762416302688e-06, 
    1.0699234287031042e-06, 1.0336145329941542e-06, 9.9849381596178131e-07, 
    9.6450859935868457e-07, 9.3160990943119202e-07, 8.9975300851207107e-07, 
    8.688978209173264e-07, 8.3900924841582014e-07, 8.1005735342350395e-07, 
    7.8201737288711222e-07, 7.5486951708747969e-07, 7.2859851114603938e-07, 
    7.0319285357444029e-07, 6.7864379580531964e-07, 6.5494408388091215e-07, 
    6.3208654314760242e-07, 6.1006262011833836e-07, 5.8886101689838837e-07, 
    5.684665564446787e-07, 5.4885940063863346e-07, 5.300147080194969e-07, 
    5.1190276997361102e-07, 4.9448960942639891e-07, 4.7773797382836899e-07, 
    4.6160861143741274e-07, 4.4606169361713985e-07, 4.3105823805264946e-07, 
    4.1656139963460641e-07, 4.0253752278596337e-07, 3.8895688699690716e-07, 
    3.7579411844909244e-07, 3.6302827965460902e-07, 3.5064267934196811e-07, 
    3.3862446474208566e-07, 3.2696406567491542e-07, 3.1565455708012414e-07, 
    3.0469099572246772e-07, 2.9406977267953568e-07, 2.8378800836274313e-07, 
    2.738430053606938e-07, 2.6423176681592501e-07, 2.5495058553791017e-07, 
    2.4599470953403e-07, 2.3735809243206543e-07, 2.2903323898034137e-07, 
    2.2101115601793447e-07, 2.1328141565853914e-07, 2.0583233103707775e-07, 
    1.9865123555195947e-07, 1.9172484665994402e-07, 1.8503968574525793e-07, 
    1.7858251927968767e-07, 1.7234078347283039e-07, 1.6630295671016458e-07, 
    1.6045884976091193e-07, 1.5479979320898942e-07, 1.493187120631299e-07, 
    1.4401008877646518e-07, 1.3886982484554256e-07, 1.3389501840168111e-07, 
    1.2908367873194324e-07, 1.2443440009272688e-07, 1.1994601597332665e-07, 
    1.1561725321754746e-07, 1.1144640299297829e-07, 1.0743102425611519e-07, 
    1.0356769430176612e-07, 9.9851820961034048e-08, 9.6277530424964185e-08, 
    9.2837643642705548e-08, 8.9523751007738915e-08, 8.6326390102498901e-08, 
    8.323532361045115e-08, 8.0239905702419762e-08, 7.7329515306122385e-08, 
    7.4494026129230937e-08, 7.1724276554145335e-08, 6.9012499923547068e-08, 
    6.6352676963670431e-08, 6.3740778431094894e-08, 6.1174875690678262e-08, 
    5.8655109879038421e-08, 5.6183523563054728e-08, 5.376377180900678e-08, 
    5.1400739555377968e-08, 4.9100098913852479e-08, 4.686784211106823e-08, 
    4.4709824383745549e-08, 4.263134594538289e-08, 4.0636795655386878e-08, 
    3.8729371283769595e-08, 3.6910884774023156e-08, 3.5181655121400537e-08, 
    3.354048791968121e-08, 3.1984737837277831e-08, 3.0510448654944176e-08, 
    2.9112563353023454e-08, 2.7785194302391509e-08, 2.6521939733414642e-08, 
    2.5316228536158634e-08, 2.4161670692879071e-08, 2.3052387441624808e-08, 
    2.1983293580327236e-08, 2.0950306180542109e-08, 1.9950458768810593e-08, 
    1.8981908645899278e-08, 1.8043835540530416e-08, 1.7136241965426388e-08, 
    1.6259676714793512e-08, 1.5414912209739696e-08, 1.4602611605672759e-08, 
    1.382302280853975e-08, 1.3075732720692681e-08, 1.2359507833285648e-08, 
    1.1672236642568218e-08, 1.1010978038187119e-08, 1.0372108080336165e-08, 
    9.7515480191135186e-09, 9.1450488461546905e-09, 8.5485037460312395e-09, 
    7.9582584769452328e-09, 7.371391697745613e-09, 6.7859409828743088e-09, 
    6.2010561222793803e-09, 5.6170675213207217e-09, 5.0354647587705433e-09, 
    4.4587869748252233e-09, 3.8904336465478317e-09, 3.3344099237764835e-09, 
    2.7950258903976279e-09, 2.2765725657729212e-09, 1.7829997279605643e-09, 
    1.3176205486069584e-09, 8.8286636297621486e-10, 4.8011072561513941e-10, 
    1.0957636458401432e-10, -2.2966859519789574e-10, -5.396263198163941e-10, 
    -8.2320582862930282e-10, -1.0839958295315285e-09, 
    -1.3259945742392218e-09, -1.5533201802421004e-09, 
    -1.7699257746829723e-09, -1.9793419134721791e-09, 
    -2.1844653789509415e-09, -2.3874081012606662e-09, 
    -2.5894142795509299e-09, -2.790847420117457e-09, -2.9912435241998347e-09, 
    -3.1894216567804004e-09, -3.38363968859506e-09, -3.5717805319856834e-09, 
    -3.7515534462451478e-09, -3.9206949913179557e-09, 
    -4.0771556714253707e-09, -4.2192600241475327e-09, 
    -4.3458307207934366e-09, -4.4562698926510043e-09, 
    -4.5505942830357385e-09, -4.629423832310123e-09, -4.6939267863473513e-09, 
    -4.745727153881496e-09, -4.7867832957840628e-09, -4.8192482112602696e-09, 
    -4.8453235911818281e-09, -4.8671196719590305e-09, 
    -4.8865323196957213e-09, -4.9051465479184971e-09, 
    -4.9241730735877166e-09, -4.9444206998014175e-09, 
    -4.9663039107676769e-09, -4.9898813414458488e-09, 
    -5.0149182550882123e-09, -5.040964162326406e-09, -5.0674364015096006e-09, 
    -5.0937009208229275e-09, -5.1191432736933648e-09, 
    -5.1432249522674674e-09, -5.1655228264167282e-09, -5.185751570639284e-09, 
    -5.203770940845878e-09, -5.2195806406231634e-09, -5.2333060631346615e-09, 
    -5.2451776467634577e-09, -5.2555061621520299e-09, 
    -5.2646552257906838e-09, -5.2730119326850732e-09, 
    -5.2809559852253254e-09, -5.2888280544448857e-09, 
    -5.2968984251045446e-09, -5.3053378403116416e-09, 
    -5.3141929178213051e-09, -5.3233691602119294e-09, -5.332624268578172e-09, 
    -5.3415741335688842e-09, -5.3497125733868974e-09, 
    -5.3564445847209877e-09, -5.3611311117086676e-09, 
    -5.3631419403249642e-09, -5.3619120298238973e-09, 
    -5.3569961069583244e-09, -5.348116171606798e-09, -5.3351973962279625e-09, 
    -5.3183888250283007e-09, -5.2980669959563197e-09, 
    -5.2748219943190265e-09, -5.2494272357806711e-09, -5.22279534115532e-09, 
    -5.1959236867473402e-09, -5.1698335578124835e-09, 
    -5.1455073027136226e-09, -5.123827540584623e-09, -5.1055224270998177e-09, 
    -5.0911202080642046e-09, -5.0809159263632501e-09, 
    -5.0749521735244273e-09, -5.0730152054822223e-09, 
    -5.0746466037850368e-09, -5.0791699615163112e-09, 
    -5.0857308286212303e-09, -5.0933475102150441e-09, 
    -5.1009691965435478e-09, -5.1075376629239485e-09, 
    -5.1120481609597322e-09, -5.1136055152720871e-09, 
    -5.1114716311970813e-09, -5.1051016300562844e-09, 
    -5.0941666315706974e-09, -5.0785625770155458e-09, 
    -5.0584054128295679e-09, -5.0340141638406715e-09, 
    -5.0058839529055593e-09, -4.9746516993133141e-09, 
    -4.9410571384375786e-09, -4.9059018889352206e-09, 
    -4.8700086928808893e-09, -4.8341827798135125e-09, 
    -4.7991765990106983e-09, -4.7656590156769941e-09, 
    -4.7341895587984261e-09, -4.7051984042870192e-09, 
    -4.6789724566725976e-09, -4.6556481020228379e-09, 
    -4.6352108816623298e-09, -4.617502410428518e-09, -4.6022343284487098e-09, 
    -4.5890088695473161e-09, -4.5773449366629627e-09, 
    -4.5667082550977678e-09, -4.5565435137508701e-09, -4.546306370020177e-09, 
    -4.5354928950317925e-09, -4.5236644873305571e-09, 
    -4.5104664847019159e-09, -4.4956395833941104e-09, 
    -4.4790236770624223e-09, -4.4605546760178417e-09, 
    -4.4402552714631952e-09, -4.4182212805339029e-09, 
    -4.3946051583230753e-09, -4.3695985215828179e-09, 
    -4.3434150235411908e-09, -4.316274882398367e-09, -4.2883916996542543e-09, 
    -4.2599621202954406e-09, -4.2311583557535077e-09, 
    -4.2021236614157599e-09, -4.1729705225996944e-09, 
    -4.1437815156654438e-09, -4.1146125465583286e-09, -4.085498368136719e-09, 
    -4.0564599104664307e-09, -4.0275130395318209e-09, 
    -3.9986779401671178e-09, -3.9699883661002432e-09, 
    -3.9414996132052511e-09, -3.9132943258231464e-09, 
    -3.8854851358365467e-09, -3.8582136500728688e-09, 
    -3.8316454259770582e-09, -3.8059613062399267e-09, 
    -3.7813456963909318e-09, -3.7579729863651826e-09, 
    -3.7359933382362665e-09, -3.7155193826420299e-09, 
    -3.6966150517389227e-09, -3.6792877491644435e-09, 
    -3.6634844544768942e-09, -3.6490921983723461e-09, 
    -3.6359426649050987e-09, -3.6238205694079267e-09, 
    -3.6124749538096378e-09, -3.601632632829014e-09, -3.591012700884625e-09, 
    -3.5803412733543714e-09, -3.5693655078818329e-09, 
    -3.5578662323893577e-09, -3.545668411155764e-09, -3.5326490267377298e-09, 
    -3.5187417984291087e-09, -3.503938586951066e-09, -3.4882871954381375e-09, 
    -3.4718857585628248e-09, -3.4548739113828718e-09, 
    -3.4374214243516351e-09, -3.4197149718086887e-09, 
    -3.4019441962412094e-09, -3.3842880642194877e-09, 
    -3.3669027713066362e-09, -3.3499120810553905e-09, 
    -3.3334009959804626e-09, -3.3174130286269518e-09, 
    -3.3019512401886877e-09, -3.2869825432676384e-09, 
    -3.2724446758767905e-09, -3.2582547912033394e-09, -3.244318697695394e-09, 
    -3.2305396415658057e-09, -3.216825876654323e-09, -3.2030962806051151e-09, 
    -3.189283863292024e-09, -3.1753370300113697e-09, -3.1612190155280732e-09, 
    -3.1469058240438609e-09, -3.132383377511203e-09, -3.1176443256485279e-09, 
    -3.1026851641883473e-09, -3.0875039090540943e-09, 
    -3.0720986932729439e-09, -3.0564672402083589e-09, 
    -3.0406072808298294e-09, -3.0245176407910002e-09, 
    -3.0081999032184816e-09, -2.9916602851155806e-09, 
    -2.9749116052850485e-09, -2.9579749926585378e-09, -2.940881252560805e-09, 
    -2.9236715903218708e-09, -2.9063976433998579e-09, 
    -2.8891206084866636e-09, -2.8719095082158677e-09, 
    -2.8548384717064546e-09, -2.8379832522601936e-09, 
    -2.8214170358317401e-09, -2.8052059781853977e-09, 
    -2.7894046962334713e-09, -2.7740522956993042e-09, 
    -2.7591692426044733e-09, -2.7447555881026585e-09, 
    -2.7307907140799082e-09, -2.7172347968344745e-09, 
    -2.7040318327121051e-09, -2.6911140095529888e-09, 
    -2.6784068960093584e-09, -2.6658349792548132e-09, 
    -2.6533268287816073e-09, -2.6408194546412924e-09, 
    -2.6282613034172289e-09, -2.615613761438671e-09, -2.6028510156702541e-09, 
    -2.5899585545220223e-09, -2.5769305523500192e-09, 
    -2.5637667092339618e-09, -2.5504689380147302e-09, -2.537038467962656e-09, 
    -2.5234736291882339e-09, -2.5097686628703775e-09, 
    -2.4959135081935207e-09, -2.4818946012172643e-09, 
    -2.4676963970193206e-09, -2.453303457592719e-09, -2.4387026900843022e-09, 
    -2.4238855821774869e-09, -2.4088500639971996e-09, 
    -2.3936019443212189e-09, -2.3781556903959792e-09, 
    -2.3625346046420589e-09, -2.346770304766954e-09, -2.3309016575471839e-09, 
    -2.3149731513479397e-09, -2.2990329278080902e-09, 
    -2.2831305135881682e-09, -2.2673145242279029e-09, 
    -2.2516304023021588e-09, -2.2361184742821407e-09, 
    -2.2208123830933513e-09, -2.2057381148341319e-09, 
    -2.1909136029288473e-09, -2.1763490069088932e-09, 
    -2.1620475276307938e-09, -2.1480067066198587e-09, 
    -2.1342199509889015e-09, -2.1206781893808034e-09, 
    -2.1073713225147354e-09, -2.0942894078207797e-09, 
    -2.0814233542477167e-09, -2.0687651539588676e-09, 
    -2.0563075922946786e-09, -2.0440436239439284e-09, 
    -2.0319654684142669e-09, -2.0200637297158068e-09, -2.008326608131271e-09, 
    -1.9967394954806736e-09, -1.9852849606838486e-09, 
    -1.9739432710240552e-09, -1.9626933525024677e-09, 
    -1.9515141574397597e-09, -1.9403862529904662e-09, 
    -1.9292935105621765e-09, -1.9182246493086911e-09, 
    -1.9071745797370888e-09, -1.896145299721411e-09, -1.8851463643345457e-09, 
    -1.8741948270634943e-09, -1.8633147104645164e-09, 
    -1.8525359858894447e-09, -1.8418931901992681e-09, -1.831423680004336e-09, 
    -1.821165681694556e-09, -1.8111561448621235e-09, -1.8014285701701555e-09, 
    -1.7920108488503291e-09, -1.7829233012134739e-09, 
    -1.7741769822217268e-09, -1.7657724456017413e-09, 
    -1.7576990393814293e-09, -1.7499348938533239e-09, -1.742447586872509e-09, 
    -1.7351955649640064e-09, -1.7281301716367982e-09, 
    -1.7211982210046441e-09, -1.7143448506987354e-09, 
    -1.7075164840534956e-09, -1.7006636012650279e-09, 
    -1.6937431564959599e-09, -1.6867204001970504e-09, 
    -1.6795700656507242e-09, -1.6722768309868563e-09, 
    -1.6648351742075785e-09, -1.6572486672483197e-09, -1.649528931044403e-09, 
    -1.6416943586634405e-09, -1.6337688074595674e-09, 
    -1.6257803135560049e-09, -1.6177599396436772e-09, 
    -1.6097406907715269e-09, -1.6017565229060835e-09, -1.593841303697508e-09, 
    -1.5860277221346679e-09, -1.578346058178075e-09, -1.5708228570750489e-09, 
    -1.5634795362874084e-09, -1.5563310753915739e-09, 
    -1.5493848902810987e-09, -1.5426401263743864e-09, 
    -1.5360874346206408e-09, -1.529709423836132e-09, -1.5234817421402828e-09, 
    -1.5173748386027908e-09, -1.5113561981351332e-09, 
    -1.5053929349645512e-09, -1.4994544554632647e-09, 
    -1.4935149913812697e-09, -1.4875556992252701e-09, 
    -1.4815661795271559e-09, -1.4755452185415453e-09, 
    -1.4695007318846252e-09, -1.463448857210691e-09, -1.4574123314422244e-09, 
    -1.4514182340779945e-09, -1.4454953476220011e-09, 
    -1.4396712879782047e-09, -1.4339696929574733e-09, 
    -1.4284076349635554e-09, -1.4229935271947852e-09, 
    -1.4177256338408566e-09, -1.4125913700610286e-09, 
    -1.4075674215258083e-09, -1.4026207643259552e-09, 
    -1.3977104782026598e-09, -1.3927903321137545e-09, 
    -1.3878119037494314e-09, -1.3827280815747167e-09, 
    -1.3774966429401758e-09, -1.372083686783502e-09, -1.3664665670885074e-09, 
    -1.3606361406050393e-09, -1.354598045136981e-09, -1.3483729330231565e-09, 
    -1.3419955242053145e-09, -1.3355126010559975e-09, 
    -1.3289799952393523e-09, -1.3224588765022175e-09, 
    -1.3160115621340726e-09, -1.3096972379373762e-09, -1.303567896206326e-09, 
    -1.2976648597555354e-09, -1.2920161057542369e-09, 
    -1.2866346316217675e-09, -1.2815179163801672e-09, 
    -1.2766485255144948e-09, -1.2719956985089181e-09, 
    -1.2675178100711627e-09, -1.263165399737704e-09, -1.2588845676244636e-09, 
    -1.2546203966172503e-09, -1.2503201879638731e-09, 
    -1.2459362504469577e-09, -1.2414281429152205e-09, -1.236764176558636e-09, 
    -1.2319222338432034e-09, -1.2268898531971617e-09, 
    -1.2216637260740364e-09, -1.2162486545063747e-09, 
    -1.2106561795214919e-09, -1.2049029671612872e-09, 
    -1.1990091796146588e-09, -1.1929968718763263e-09, -1.186888643442219e-09, 
    -1.1807065113419187e-09, -1.1744711417912692e-09, 
    -1.1682013889407819e-09, -1.1619141927736853e-09, 
    -1.1556247006616581e-09, -1.1493466382339949e-09, 
    -1.1430927603657763e-09, -1.1368753742281928e-09, 
    -1.1307067683277524e-09, -1.1245995549174521e-09, 
    -1.1185667933570186e-09, -1.11262194141667e-09, -1.1067785575113433e-09, 
    -1.1010498372626891e-09, -1.095447973758005e-09, -1.0899834711782896e-09, 
    -1.0846643967476001e-09, -1.0794957395418595e-09, 
    -1.0744788505687392e-09, -1.0696111099834175e-09, 
    -1.0648857623048258e-09, -1.0602920441613919e-09, 
    -1.0558154917186889e-09, -1.0514385186649444e-09, 
    -1.0471411299572191e-09, -1.042901800959198e-09, -1.0386983975015271e-09, 
    -1.0345091589256059e-09, -1.0303135833729443e-09, -1.026093253474246e-09, 
    -1.0218324798711319e-09, -1.0175187957935122e-09, 
    -1.0131432102985075e-09, -1.0087002990945804e-09, 
    -1.0041880668036317e-09, -9.9960768082437195e-10, -9.949630546060814e-10, 
    -9.9026040307238079e-10, -9.8550772631551035e-10, 
    -9.8071435969749488e-10, -9.7589053065296843e-10, 
    -9.7104703584632095e-10, -9.6619494467904622e-10, 
    -9.6134541905025713e-10, -9.565095303375199e-10, -9.5169816306729656e-10, 
    -9.4692186397920475e-10, -9.4219071967412737e-10, 
    -9.3751416719289535e-10, -9.3290081577204547e-10, 
    -9.2835820320775992e-10, -9.2389258602526849e-10, 
    -9.1950870371307321e-10, -9.1520963687572222e-10, 
    -9.1099665441218493e-10, -9.0686923124604386e-10, 
    -9.0282507324886025e-10, -8.9886030091869474e-10, 
    -8.9496967372127469e-10, -8.9114693834832565e-10, 
    -8.8738517810487422e-10, -8.8367724998836875e-10, 
    -8.8001616272713547e-10, -8.7639548015136228e-10, 
    -8.7280961716083973e-10, -8.6925409937572383e-10, -8.65725674406098e-10, 
    -8.6222235914026509e-10, -8.5874332437941012e-10, 
    -8.5528871950155082e-10, -8.5185936364417731e-10, 
    -8.4845642466497022e-10, -8.4508102184421245e-10, 
    -8.4173388175044866e-10, -8.3841498720586671e-10, 
    -8.3512334913850891e-10, -8.3185682260326587e-10, 
    -8.2861205543909451e-10, -8.2538450032638922e-10, 
    -8.2216856690700295e-10, -8.1895777840265951e-10, -8.15745048641611e-10, 
    -8.1252292630345012e-10, -8.0928391040108165e-10, -8.060207218400921e-10, 
    -8.0272663192383884e-10, -7.9939574356522857e-10, 
    -7.9602332607544061e-10, -7.9260611745253683e-10, 
    -7.8914266350209369e-10, -7.8563360075665521e-10, 
    -7.8208194377408362e-10, -7.7849324940464251e-10, 
    -7.7487570674416999e-10, -7.7124003020894752e-10, 
    -7.6759921906327137e-10, -7.6396806765082959e-10, 
    -7.6036252655742127e-10, -7.5679885915086446e-10, 
    -7.5329273320708331e-10, -7.4985823432680116e-10, 
    -7.4650697480649062e-10, -7.4324731073921192e-10, 
    -7.4008382331967127e-10, -7.3701706291935606e-10, 
    -7.3404366486116639e-10, -7.3115676173130518e-10, 
    -7.2834674571335637e-10, -7.2560221759543096e-10, 
    -7.2291114261352983e-10, -7.2026197497005282e-10, 
    -7.1764475567789064e-10, -7.150519741650857e-10, -7.1247916498577136e-10, 
    -7.0992514412264792e-10, -7.0739188567042471e-10, 
    -7.0488400472932045e-10, -7.0240795624611714e-10, 
    -6.9997095445687076e-10, -6.97579805226613e-10, -6.9523967341263158e-10, 
    -6.9295300826645623e-10, -6.9071865118787122e-10, 
    -6.8853128684625362e-10, -6.8638125795355857e-10, 
    -6.8425479842826447e-10, -6.8213465631092137e-10, 
    -6.8000107924490402e-10, -6.7783305146253801e-10, 
    -6.7560973314565593e-10, -6.7331191702967465e-10, 
    -6.7092345845246864e-10, -6.684325035262447e-10, -6.658324893074484e-10, 
    -6.6312278093421423e-10, -6.6030897888800856e-10, 
    -6.5740280482725389e-10, -6.5442164222719162e-10, 
    -6.5138770522127833e-10, -6.4832693716267691e-10, 
    -6.4526763933222766e-10, -6.4223897356182132e-10, 
    -6.3926934351942475e-10, -6.3638482278194757e-10, 
    -6.3360765444949181e-10, -6.3095496412764992e-10, 
    -6.2843774256844473e-10, -6.2606019273845558e-10, 
    -6.2381947924051666e-10, -6.2170593202580097e-10, 
    -6.1970367841500283e-10, -6.1779170067374804e-10, 
    -6.1594521875260598e-10, -6.1413734890217602e-10, 
    -6.1234087171340747e-10, -6.1053003128176867e-10, 
    -6.0868219477659275e-10, -6.0677927840109198e-10, 
    -6.0480881147262466e-10, -6.0276459605436483e-10, 
    -6.0064687950977952e-10, -5.984620800030318e-10, -5.9622205228344642e-10, 
    -5.9394302045376474e-10, -5.9164419362154322e-10, 
    -5.8934627562038493e-10, -5.870698969336033e-10, -5.8483416578125842e-10, 
    -5.8265538832777278e-10, -5.8054609308520137e-10, 
    -5.7851436972137075e-10, -5.7656357367973167e-10, 
    -5.7469238000741915e-10, -5.7289514845735051e-10, 
    -5.7116253745476449e-10, -5.6948230461081153e-10, -5.678402040928712e-10, 
    -5.6622093094363476e-10, -5.6460901225938823e-10, 
    -5.6298965826691411e-10, -5.6134947400469541e-10, 
    -5.5967707258365599e-10, -5.5796354803564643e-10, 
    -5.5620283554968852e-10, -5.543919358338596e-10, -5.5253104133531056e-10, 
    -5.5062353184652853e-10, -5.4867586284736606e-10, 
    -5.4669733173540123e-10, -5.4469972509355413e-10, 
    -5.4269683278178332e-10, -5.4070388525665661e-10, 
    -5.3873686052971397e-10, -5.3681175312533896e-10, 
    -5.3494379500936851e-10, -5.331466963949267e-10, -5.3143193830222798e-10, 
    -5.2980815453305014e-10, -5.2828065267750357e-10, 
    -5.2685109071600257e-10, -5.255173226962127e-10, -5.2427344115952453e-10, 
    -5.2310996990820243e-10, -5.220142323889685e-10, -5.2097083751249536e-10, 
    -5.1996227474603015e-10, -5.1896958428034411e-10, 
    -5.1797306573675232e-10, -5.1695300864661643e-10, 
    -5.1589041878301825e-10, -5.1476771408755447e-10, 
    -5.1356936755011064e-10, -5.1228248694078628e-10, -5.108973015142107e-10, 
    -5.0940753920019648e-10, -5.0781068729629399e-10, -5.06108102539727e-10, 
    -5.0430498271276111e-10, -5.0241017602642855e-10, -5.004358642296449e-10, 
    -4.9839709705561459e-10, -4.9631121885763852e-10, 
    -4.9419720498433616e-10, -4.9207493576852637e-10, 
    -4.8996443658920321e-10, -4.8788510955716544e-10, 
    -4.8585497908962362e-10, -4.8388999342966207e-10, 
    -4.8200337808492722e-10, -4.802050934375583e-10, -4.7850139481893043e-10, 
    -4.7689452818970242e-10, -4.7538258559478753e-10, 
    -4.7395951932774082e-10, -4.7261535069315454e-10, 
    -4.7133656063396707e-10, -4.7010666315549495e-10, 
    -4.6890693828026452e-10, -4.6771730533166562e-10, 
    -4.6651729436031745e-10, -4.6528705027143202e-10, 
    -4.6400834932023453e-10, -4.6266552749276909e-10, 
    -4.6124629781090838e-10, -4.5974238854938427e-10, 
    -4.5814997758280726e-10, -4.5646986882399501e-10, -4.547074410618504e-10, 
    -4.5287232006620904e-10, -4.5097782168971026e-10, 
    -4.4904018160950881e-10, -4.4707761570476444e-10, 
    -4.4510925220804004e-10, -4.4315399698089313e-10, -4.412293878576717e-10, 
    -4.3935052053320076e-10, -4.3752908209625582e-10, 
    -4.3577259340175198e-10, -4.3408387946820195e-10, 
    -4.3246084555011958e-10, -4.3089656074691887e-10, 
    -4.2937968297078225e-10, -4.2789518078599878e-10, 
    -4.2642534086155211e-10, -4.2495096230106152e-10, 
    -4.2345269579711351e-10, -4.2191239098592065e-10, 
    -4.2031438162958002e-10, -4.1864658763550055e-10, 
    -4.1690139200790382e-10, -4.1507618118198311e-10, 
    -4.1317355414328092e-10, -4.1120118073127928e-10, -4.091713338004328e-10, 
    -4.0710012984559772e-10, -4.0500657588143459e-10, 
    -4.0291146152223975e-10, -4.0083620139004865e-10, 
    -3.9880170771979457e-10, -3.9682734773183607e-10, -3.949300523111033e-10, 
    -3.9312362247123504e-10, -3.9141822295503037e-10, 
    -3.8982012360089874e-10, -3.883316075139802e-10, -3.8695109341600564e-10, 
    -3.856733897306086e-10, -3.8449009474400284e-10, -3.8339007069768565e-10, 
    -3.8236000699697306e-10, -3.8138500495388374e-10, 
    -3.8044921153075135e-10, -3.7953645141594882e-10, -3.786308641540416e-10, 
    -3.7771751967270152e-10, -3.7678302671855809e-10, 
    -3.7581606979831276e-10, -3.7480790648550088e-10, 
    -3.7375274957551404e-10, -3.7264805520781431e-10, 
    -3.7149464067097481e-10, -3.7029667403686127e-10, 
    -3.6906145059181719e-10, -3.6779902266111028e-10, 
    -3.6652162294389059e-10, -3.6524297810978628e-10, 
    -3.6397747774476797e-10, -3.627392981600115e-10, -3.6154149670945044e-10, 
    -3.603951723036565e-10, -3.5930870852746917e-10, -3.5828718858827313e-10, 
    -3.5733197688254365e-10, -3.5644055674997457e-10, 
    -3.5560656188792085e-10, -3.5482005922377747e-10, 
    -3.5406801991202822e-10, -3.5333497496227482e-10, 
    -3.5260378945383196e-10, -3.5185653034912508e-10, 
    -3.5107534616227477e-10, -3.5024334951676399e-10, 
    -3.4934541408615431e-10, -3.4836889760095792e-10, 
    -3.4730419793357588e-10, -3.4614519489267041e-10, 
    -3.4488948613564403e-10, -3.4353847816071349e-10, 
    -3.4209727184440522e-10, -3.4057441188331918e-10, 
    -3.3898144572638057e-10, -3.373323819884734e-10, -3.3564300162672814e-10, 
    -3.3393013331298188e-10, -3.3221084402572002e-10, 
    -3.3050166898169108e-10, -3.2881785023568738e-10, 
    -3.2717267946826903e-10, -3.2557692407895179e-10, 
    -3.2403844288372453e-10, -3.2256191140999258e-10, 
    -3.2114877922075152e-10, -3.197973586163585e-10, -3.1850312160729096e-10, 
    -3.1725912695877147e-10, -3.1605659118082819e-10, 
    -3.1488555354939759e-10, -3.137356082313803e-10, -3.1259663377826575e-10, 
    -3.1145953973392076e-10, -3.1031688649067593e-10, 
    -3.0916344573983715e-10, -3.0799656128480821e-10, 
    -3.0681636060711769e-10, -3.0562572888856871e-10, 
    -3.0443011433289781e-10, -3.032370893842879e-10, -3.0205578425555211e-10, 
    -3.0089614724562719e-10, -2.9976816313050547e-10, 
    -2.9868102560135458e-10, -2.9764238237928843e-10, 
    -2.9665766318997044e-10, -2.9572960642140459e-10, 
    -2.9485795669769855e-10, -2.9403942829158665e-10, -2.932678792189975e-10, 
    -2.9253473931076426e-10, -2.9182960184610318e-10, 
    -2.9114100239137388e-10, -2.9045723686598534e-10, 
    -2.8976724795127352e-10, -2.8906141495746108e-10, 
    -2.8833226042765249e-10, -2.8757495174507703e-10, 
    -2.8678762759199327e-10, -2.8597143473695148e-10, 
    -2.8513039686466934e-10, -2.8427100284328622e-10, 
    -2.8340167359670204e-10, -2.8253206060795276e-10, 
    -2.8167233628887791e-10, -2.8083243548358648e-10, 
    -2.8002140880451542e-10, -2.7924684397791852e-10, 
    -2.7851447134117877e-10, -2.778278922579416e-10, -2.7718851492443711e-10, 
    -2.7659560117416318e-10, -2.7604648129687695e-10, 
    -2.7553683217063748e-10, -2.7506106839197323e-10, 
    -2.7461272836218177e-10, -2.7418491865924319e-10, 
    -2.7377070505035443e-10, -2.7336350454178157e-10, 
    -2.7295739850871216e-10, -2.7254742627118688e-10, 
    -2.7212976052890382e-10, -2.7170184345045745e-10, 
    -2.7126240504446712e-10, -2.7081142080633844e-10, 
    -2.7034995214696081e-10, -2.6987994886680448e-10, 
    -2.6940394741713519e-10, -2.6892476030628745e-10, 
    -2.6844511138234363e-10, -2.6796731631789273e-10, 
    -2.6749295858621813e-10, -2.6702265825794055e-10, 
    -2.6655589226588525e-10, -2.660909393033198e-10, -2.6562489688936634e-10, 
    -2.6515383320598089e-10, -2.6467299850835136e-10, 
    -2.6417715783386226e-10, -2.6366094760130453e-10, 
    -2.6311929581998298e-10, -2.6254782130514547e-10, 
    -2.6194324275671379e-10, -2.6130369580885922e-10, 
    -2.6062899641712782e-10, -2.5992076031220241e-10, 
    -2.5918242942533302e-10, -2.5841911928069096e-10, 
    -2.5763736443302461e-10, -2.5684471541416006e-10, 
    -2.5604926019231889e-10, -2.552590593552168e-10, -2.5448161297938444e-10, 
    -2.5372331644137877e-10, -2.5298903837183557e-10, 
    -2.5228178142228935e-10, -2.5160254268594921e-10, 
    -2.5095029389067192e-10, -2.5032216465598918e-10, 
    -2.4971374636963314e-10, -2.4911954747745169e-10, 
    -2.4853350350815109e-10, -2.4794955040511736e-10, 
    -2.4736215780699755e-10, -2.467668353483063e-10, -2.4616050913339002e-10, 
    -2.4554180197832519e-10, -2.4491112815452816e-10, 
    -2.4427067357170691e-10, -2.436241914666686e-10, -2.429767049058874e-10, 
    -2.4233409277629974e-10, -2.4170263772106145e-10, -2.410885466161698e-10, 
    -2.4049752644926131e-10, -2.3993440036651042e-10, 
    -2.3940284041603184e-10, -2.3890517912620046e-10, 
    -2.3844236399864125e-10, -2.3801398562324482e-10, 
    -2.3761838970487604e-10, -2.3725282357813226e-10, 
    -2.3691364641272979e-10, -2.3659649052769033e-10, 
    -2.3629642604792017e-10, -2.3600806880664621e-10, 
    -2.3572568563081836e-10, -2.3544322758449895e-10, 
    -2.3515438381563081e-10, -2.3485261408962341e-10, -2.345312198560387e-10, 
    -2.3418344678942607e-10, -2.3380266624698267e-10, 
    -2.3338259102382919e-10, -2.3291757815849845e-10, 
    -2.3240294942444497e-10, -2.3183535104985747e-10, 
    -2.3121307266616651e-10, -2.305363381392176e-10, -2.2980746694360122e-10, 
    -2.2903093645822175e-10, -2.2821326670531984e-10, 
    -2.2736276640507036e-10, -2.2648909910133832e-10, 
    -2.2560276478406723e-10, -2.2471446788950895e-10, 
    -2.2383449144001749e-10, -2.229720816168745e-10, -2.2213496582140858e-10, 
    -2.2132897598414773e-10, -2.2055786920923755e-10, 
    -2.1982330499015747e-10, -2.1912501182555217e-10, 
    -2.1846105448249568e-10, -2.1782822068233226e-10, 
    -2.1722240626020924e-10, -2.1663901787880501e-10, 
    -2.1607329792069826e-10, -2.155206071409944e-10, -2.1497660322494598e-10, 
    -2.1443738776245511e-10, -2.1389959187336111e-10, -2.133604848327161e-10, 
    -2.1281807726317722e-10, -2.1227128773411828e-10, -2.117201205808825e-10, 
    -2.1116590044255405e-10, -2.1061146958896203e-10, 
    -2.1006135170938521e-10, -2.0952180464017519e-10, 
    -2.0900075947351466e-10, -2.0850756304781097e-10, 
    -2.0805257185356009e-10, -2.0764656398278498e-10, 
    -2.0730003128267641e-10, -2.0702237648954901e-10, 
    -2.0682113686925689e-10, -2.0670123007246921e-10, 
    -2.0666435167588897e-10, -2.0670854698331876e-10, 
    -2.0682802998540831e-10, -2.0701321754724024e-10, 
    -2.0725102959006022e-10, -2.0752537609044974e-10, 
    -2.0781783374843521e-10, -2.0810840804184689e-10, 
    -2.0837637637217375e-10, -2.0860109006858191e-10, -2.087627625871134e-10, 
    -2.0884314657372983e-10, -2.088261306618446e-10, -2.0869821188190646e-10, 
    -2.0844891411908311e-10, -2.0807109643290825e-10, 
    -2.0756121914809179e-10, -2.0691954764839816e-10, 
    -2.0615030906900754e-10, -2.052617577262212e-10, -2.0426616702274237e-10, 
    -2.0317966083098877e-10, -2.020218873804839e-10, -2.0081547749539571e-10, 
    -1.9958532443193001e-10, -1.9835762451283037e-10, 
    -1.9715877232192627e-10, -1.9601412016434301e-10, 
    -1.9494674020985858e-10, -1.9397620582303722e-10, -1.931175522588158e-10, 
    -1.9238045694112204e-10, -1.9176876023821112e-10, 
    -1.9128031976803019e-10, -1.9090726991609491e-10, 
    -1.9063661686406626e-10, -1.9045119350729719e-10, 
    -1.9033082834655493e-10, -1.9025370397228457e-10, 
    -1.9019775628578702e-10, -1.9014203504056245e-10, 
    -1.9006790344534291e-10, -1.89960023220148e-10, -1.8980700439176426e-10, 
    -1.8960173642585568e-10, -1.8934133955150964e-10, 
    -1.8902678801146103e-10, -1.8866223711871336e-10, 
    -1.8825413872127897e-10, -1.8781021766049117e-10, 
    -1.8733845686728914e-10, -1.8684612608651276e-10, 
    -1.8633901126651848e-10, -1.8582085038820917e-10, 
    -1.8529308197513185e-10, -1.8475484188014905e-10, 
    -1.8420323747402076e-10, -1.8363381877924191e-10, 
    -1.8304119833922716e-10, -1.8241970660854944e-10, 
    -1.8176405074295455e-10, -1.8106986285973861e-10, 
    -1.8033414111820881e-10, -1.7955550986411724e-10, 
    -1.7873434461317491e-10, -1.7787273636658396e-10, 
    -1.7697437442647195e-10, -1.7604433848692879e-10, 
    -1.7508887885216284e-10, -1.7411518621855021e-10, -1.731312075579559e-10, 
    -1.72145467512114e-10, -1.7116696280453247e-10, -1.7020504552884229e-10, 
    -1.6926934109626932e-10, -1.6836962556930328e-10, 
    -1.6751570906481501e-10, -1.6671724116693748e-10, 
    -1.6598348070561075e-10, -1.6532299159429898e-10, -1.647433173183042e-10, 
    -1.6425058537389233e-10, -1.6384911983556137e-10, 
    -1.6354105157628102e-10, -1.6332598611774752e-10, 
    -1.6320072533744398e-10, -1.6315914347278538e-10, 
    -1.6319217555223467e-10, -1.6328798506368337e-10, 
    -1.6343231081872432e-10, -1.6360899991816905e-10, 
    -1.6380067166199145e-10, -1.6398952564863494e-10, 
    -1.6415818802385306e-10, -1.6429057708670176e-10, -1.643726758427863e-10, 
    -1.6439320169385336e-10, -1.6434405136432045e-10, -1.642205399414063e-10, 
    -1.64021377487063e-10, -1.6374841222870594e-10, -1.6340614420746998e-10, 
    -1.6300109407985323e-10, -1.6254104057701017e-10, 
    -1.6203424831251957e-10, -1.6148871101108542e-10, 
    -1.6091150889099701e-10, -1.6030830195437145e-10, -1.596830247150364e-10, 
    -1.5903776371786904e-10, -1.5837283983006877e-10, 
    -1.5768705770197147e-10, -1.5697810216847621e-10, 
    -1.5624302234358719e-10, -1.5547876082684374e-10, 
    -1.5468267715017817e-10, -1.5385302571453756e-10, -1.529893302818309e-10, 
    -1.5209265055085765e-10, -1.5116569033645694e-10, 
    -1.5021278158863802e-10, -1.4923970973628858e-10, 
    -1.4825341592980001e-10, -1.4726159266613504e-10, 
    -1.4627222959504513e-10, -1.4529310584525797e-10, 
    -1.4433131167292655e-10, -1.4339281050630124e-10, 
    -1.4248210157717807e-10, -1.4160200182979566e-10, 
    -1.4075357851621989e-10, -1.3993623391799455e-10, 
    -1.3914795696739524e-10, -1.383857065039665e-10, -1.3764590404322013e-10, 
    -1.3692499468505607e-10, -1.3622002331344276e-10, 
    -1.3552915731710757e-10, -1.3485214181580243e-10, 
    -1.3419058588022465e-10, -1.335481008636497e-10, -1.3293022825510545e-10, 
    -1.3234420723772461e-10, -1.3179854582146276e-10, 
    -1.3130247925774169e-10, -1.3086533384013984e-10, 
    -1.3049584689376631e-10, -1.3020151823648038e-10, 
    -1.2998802320690939e-10, -1.2985873183684268e-10, 
    -1.2981438819975705e-10, -1.2985293472332415e-10, -1.299695229405128e-10, 
    -1.3015668516603455e-10, -1.3040467135553042e-10, 
    -1.3070190968264593e-10, -1.3103557396212783e-10, -1.313922197977725e-10, 
    -1.3175844121616167e-10, -1.3212151225976705e-10, 
    -1.3246998945630893e-10, -1.3279420471496044e-10, 
    -1.3308665153818101e-10, -1.3334221681639812e-10, 
    -1.3355827874549457e-10, -1.3373463579749029e-10, 
    -1.3387330315936966e-10, -1.3397819238977436e-10, 
    -1.3405469889696475e-10, -1.3410924771246082e-10, 
    -1.3414880881019827e-10, -1.341804412440886e-10, -1.3421087823874526e-10, 
    -1.342461770735253e-10, -1.3429144228941044e-10, -1.3435062509308788e-10, 
    -1.3442639691137541e-10, -1.3452007718547825e-10, 
    -1.3463161550217811e-10, -1.3475960172743659e-10, 
    -1.3490132589754778e-10, -1.3505285084710004e-10, 
    -1.3520913108260503e-10, -1.3536417594606306e-10, 
    -1.3551125472903519e-10, -1.356431673529807e-10, -1.3575258479007305e-10, 
    -1.358324242723375e-10, -1.3587628191340216e-10, -1.3587887155516542e-10, 
    -1.3583644865661151e-10, -1.3574718137804818e-10, 
    -1.3561143293889222e-10, -1.3543191745336521e-10, 
    -1.3521371038815148e-10, -1.3496409605924764e-10, 
    -1.3469225367114248e-10, -1.3440879926900114e-10, -1.341252094278797e-10, 
    -1.3385316444668712e-10, -1.3360386465857951e-10, 
    -1.3338734640007523e-10, -1.3321188062791259e-10, 
    -1.3308345639704375e-10, -1.3300539940010912e-10, 
    -1.3297814220406498e-10, -1.3299917406726473e-10, 
    -1.3306314093057008e-10, -1.3316210353994203e-10, 
    -1.3328594269659794e-10, -1.3342287070676122e-10, 
    -1.3356002687251864e-10, -1.3368414148220662e-10, 
    -1.3378219740712827e-10, -1.3384208429731093e-10, 
    -1.3385319357584846e-10, -1.3380692517604632e-10, 
    -1.3369708007239969e-10, -1.3352011833229895e-10, 
    -1.3327527363287282e-10, -1.3296450723662447e-10, 
    -1.3259232685287485e-10, -1.3216550108773703e-10, 
    -1.3169265303641723e-10, -1.3118380625570442e-10, 
    -1.3064989025059138e-10, -1.3010225118462212e-10, 
    -1.2955218863049402e-10, -1.2901054178873341e-10, 
    -1.2848733673244812e-10, -1.27991527647119e-10, -1.2753079910275013e-10, 
    -1.2711146407924603e-10, -1.2673842528785563e-10, 
    -1.2641521720040708e-10, -1.2614409458278252e-10, 
    -1.2592617203902218e-10, -1.257615892931511e-10, -1.2564969830617307e-10, 
    -1.2558923867937309e-10, -1.2557850059132167e-10, 
    -1.2561544913459178e-10, -1.2569781041700057e-10, 
    -1.2582310625671466e-10, -1.2598863326971268e-10, 
    -1.2619140755314919e-10, -1.264280817847885e-10, -1.2669483807104051e-10, 
    -1.2698730513342003e-10, -1.2730048413747006e-10, 
    -1.2762872324101628e-10, -1.2796574128502761e-10, 
    -1.2830469016302912e-10, -1.2863827823189012e-10, 
    -1.2895892901704825e-10, -1.2925896254864172e-10, 
    -1.2953078682326049e-10, -1.2976708792529846e-10, 
    -1.2996101399694291e-10, -1.3010631873177415e-10, -1.301975023184133e-10, 
    -1.3022991628345213e-10, -1.3019983457399362e-10, 
    -1.3010451850881609e-10, -1.2994225777428153e-10, 
    -1.2971238620411277e-10, -1.2941529602930621e-10, 
    -1.2905241645804941e-10, -1.2862618141137223e-10, 
    -1.2813996581514535e-10, -1.275980007998854e-10, -1.2700524982368766e-10, 
    -1.2636727068559427e-10, -1.2569003569522523e-10, 
    -1.2497975151208163e-10, -1.2424264388967688e-10, 
    -1.2348476789160409e-10, -1.2271180862421225e-10, 
    -1.2192891671030682e-10, -1.2114057752622123e-10, 
    -1.2035053363348484e-10, -1.1956176282461056e-10, 
    -1.1877651713981299e-10, -1.1799642470356691e-10, 
    -1.1722264869430608e-10, -1.1645608265596537e-10, 
    -1.1569757390717628e-10, -1.1494814271530886e-10, 
    -1.1420918699006364e-10, -1.1348262384335057e-10, 
    -1.1277099031161572e-10, -1.1207744514019457e-10, 
    -1.1140570151179558e-10, -1.1075987121544582e-10, 
    -1.1014426221480282e-10, -1.0956312092683019e-10, 
    -1.0902035199708324e-10, -1.0851925722442701e-10, 
    -1.0806231206902125e-10, -1.0765098359384356e-10, 
    -1.0728563864263498e-10, -1.0696551475841043e-10, 
    -1.0668878609700222e-10, -1.0645268916879325e-10, 
    -1.0625371259464442e-10, -1.0608782699833751e-10, 
    -1.0595073157005915e-10, -1.058381004867868e-10, -1.0574581185394442e-10, 
    -1.0567013012546477e-10, -1.0560784418867379e-10, 
    -1.0555634073720328e-10, -1.0551361587421227e-10, 
    -1.0547822320032843e-10, -1.0544918585077048e-10, 
    -1.0542585663488874e-10, -1.0540778294328999e-10, -1.053945639753728e-10, 
    -1.0538574692667981e-10, -1.0538076020616617e-10, 
    -1.0537889979505818e-10, -1.0537936087450587e-10, 
    -1.0538132748058312e-10, -1.0538405557046931e-10, 
    -1.0538698604695897e-10, -1.0538980793077869e-10, 
    -1.0539248502406963e-10, -1.05395217205635e-10, -1.0539834191929546e-10, 
    -1.0540217475590477e-10, -1.0540683157930262e-10, 
    -1.0541202942699343e-10, -1.0541694149471697e-10, 
    -1.0542009311369249e-10, -1.0541936887171246e-10, 
    -1.0541210611397324e-10, -1.0539528957980547e-10, 
    -1.0536583583706007e-10, -1.0532092217786501e-10, 
    -1.0525833010438373e-10, -1.0517677081515204e-10, 
    -1.0507613005175672e-10, -1.0495762944098204e-10, 
    -1.0482385524444387e-10, -1.0467869273792122e-10, 
    -1.0452713345248659e-10, -1.0437499957271388e-10, 
    -1.0422861019438497e-10, -1.0409444571069991e-10, 
    -1.0397879984559918e-10, -1.0388749097991062e-10, 
    -1.0382563109142484e-10, -1.0379746355681367e-10, 
    -1.0380627875382652e-10, -1.0385439177663074e-10, 
    -1.0394316948802475e-10, -1.0407308874564264e-10, 
    -1.0424380027489405e-10, -1.0445420441365994e-10, -1.047024903328403e-10, 
    -1.0498617450280562e-10, -1.0530211490409919e-10, 
    -1.0564651264965317e-10, -1.0601492131967841e-10, 
    -1.0640228692436925e-10, -1.0680300479586959e-10, -1.072110309118443e-10, 
    -1.0762003477168159e-10, -1.0802360718426384e-10, 
    -1.0841548015089668e-10, -1.08789777407814e-10, -1.0914124180817585e-10, 
    -1.0946541771977547e-10, -1.0975876835605673e-10, 
    -1.1001872849812024e-10, -1.102436413668568e-10, -1.1043262962158351e-10, 
    -1.1058538190132427e-10, -1.107019192546185e-10, -1.1078233571036765e-10, 
    -1.1082658793273179e-10, -1.1083434843685396e-10, 
    -1.1080495230110414e-10, -1.1073744417996746e-10, 
    -1.1063074516070899e-10, -1.1048388097948467e-10, 
    -1.1029627961575233e-10, -1.1006806780596408e-10, 
    -1.0980033198959293e-10, -1.0949529645415125e-10, 
    -1.0915642058058477e-10, -1.0878834617676116e-10, 
    -1.0839674403075727e-10, -1.0798804597350134e-10, -1.075691249712976e-10, 
    -1.0714692365475537e-10, -1.0672810876410342e-10, 
    -1.0631875982847875e-10, -1.0592412993563771e-10, 
    -1.0554848890770812e-10, -1.0519505677359571e-10, 
    -1.0486598831545883e-10, -1.0456243347578916e-10, 
    -1.0428460785909132e-10, -1.0403187010367006e-10, 
    -1.0380279749095257e-10, -1.0359524082616051e-10, 
    -1.0340636041493082e-10, -1.0323265945516844e-10, 
    -1.0307002112263458e-10, -1.0291377396074527e-10, 
    -1.0275877573969529e-10, -1.0259956987142355e-10, 
    -1.0243056828501231e-10, -1.0224627727273623e-10, 
    -1.0204155282828911e-10, -1.0181187953068243e-10, 
    -1.0155361776259329e-10, -1.0126423776293402e-10, 
    -1.0094249408119783e-10, -1.0058853555237095e-10, 
    -1.0020393150971903e-10, -9.9791629059022466e-11, 
    -9.9355814404611268e-11, -9.8901713236936777e-11, -9.84353239389405e-11, 
    -9.796312336618561e-11, -9.749174304215754e-11, -9.7027669475913381e-11, 
    -9.6576959823127402e-11, -9.6145024773741303e-11, -9.573646616875994e-11, 
    -9.5354993426741204e-11, -9.5003404214562995e-11, 
    -9.4683635499624471e-11, -9.4396843416113697e-11, 
    -9.4143520456020924e-11, -9.3923601042008899e-11, 
    -9.3736555028528166e-11, -9.3581452654311781e-11, 
    -9.3456992179752979e-11, -9.3361492869355007e-11, 
    -9.3292890939254431e-11, -9.3248715708096204e-11, 
    -9.3226106028944909e-11, -9.3221854036805052e-11, 
    -9.3232514923181645e-11, -9.3254566318927731e-11, 
    -9.3284602893296274e-11, -9.3319571325152509e-11, 
    -9.3356999291305851e-11, -9.3395178358200396e-11, 
    -9.3433301116478294e-11, -9.347148111101928e-11, -9.3510682579869108e-11, 
    -9.3552520429353483e-11, -9.3598962152424882e-11, 
    -9.3651955133128663e-11, -9.3713015510049357e-11, 
    -9.3782823903726995e-11, -9.386089224066176e-11, -9.3945341249162906e-11, 
    -9.4032819682884528e-11, -9.4118617053778014e-11, 
    -9.4196950108658373e-11, -9.4261426837346703e-11, 
    -9.4305632772487179e-11, -9.4323793450141094e-11, 
    -9.4311462475627908e-11, -9.4266128554906555e-11, 
    -9.4187691341467619e-11, -9.4078748214102842e-11, 
    -9.3944644341492294e-11, -9.3793280592726336e-11, 
    -9.3634685298645754e-11, -9.3480381433231532e-11, -9.334262914743822e-11, 
    -9.3233596524378346e-11, -9.3164529090160246e-11, 
    -9.3145013701086279e-11, -9.318239455173144e-11, -9.3281367335121854e-11, 
    -9.3443780823434661e-11, -9.3668664108596487e-11, 
    -9.3952443921309634e-11, -9.4289329443095036e-11, 
    -9.4671801388175887e-11, -9.5091186689444808e-11, -9.553825062280098e-11, 
    -9.6003756417707625e-11, -9.6478969266327101e-11, 
    -9.6956057790019833e-11, -9.7428377314750928e-11, 
    -9.7890613512930015e-11, -9.8338799518177515e-11, 
    -9.8770194694280509e-11, -9.9183042382436654e-11, -9.957624337231556e-11, 
    -9.9948969459687538e-11, -1.0030024963377561e-10, 
    -1.0062857950179827e-10, -1.0093159195980151e-10, 
    -1.0120582338569124e-10, -1.0144660778922387e-10, 
    -1.0164811313167535e-10, -1.0180353910274087e-10, 
    -1.0190543165684371e-10, -1.019461342255508e-10, -1.0191830643399935e-10, 
    -1.0181547261587496e-10, -1.0163256474989071e-10, 
    -1.0136638916397364e-10, -1.0101599331769694e-10, 
    -1.0058289432173381e-10, -1.0007115677910779e-10, 
    -9.9487318408161817e-11, -9.8840171330817425e-11, 
    -9.8140433186245164e-11, -9.7400326079160308e-11, 
    -9.6633115751075823e-11, -9.5852617781203409e-11, 
    -9.5072715672451617e-11, -9.4306908606072075e-11, -9.356788084279663e-11, 
    -9.2867120606125114e-11, -9.2214579265484998e-11, 
    -9.1618368203069536e-11, -9.1084520640829237e-11, 
    -9.0616802121824287e-11, -9.0216617213848282e-11, 
    -8.9883009822399395e-11, -8.961279785907028e-11, -8.940083323218561e-11, 
    -8.9240418624754513e-11, -8.9123854657617492e-11, 
    -8.9043090717919227e-11, -8.899044600437618e-11, -8.8959332610167114e-11, 
    -8.8944912254382773e-11, -8.8944623418256101e-11, -8.895850608547336e-11, 
    -8.8989287429791831e-11, -8.9042171112145325e-11, 
    -8.9124360141414728e-11, -8.9244330858708781e-11, 
    -8.9410899421678659e-11, -8.9632183009813508e-11, -8.991453661574089e-11, 
    -9.0261588463273042e-11, -9.0673457584053032e-11, 
    -9.1146248454835027e-11, -9.1671884565006293e-11, 
    -9.2238302259427116e-11, -9.2829997800126581e-11, 
    -9.3428884345360168e-11, -9.4015383799636098e-11, 
    -9.4569636884414583e-11, -9.5072756916676917e-11, 
    -9.5507975038351159e-11, -9.5861618147616192e-11, 
    -9.6123822676217446e-11, -9.6288957207732643e-11, 
    -9.6355732219031399e-11, -9.6327024755100875e-11, 
    -9.6209447427697103e-11, -9.6012748076735564e-11, 
    -9.5749073046277841e-11, -9.5432193728520331e-11, 
    -9.5076726989006318e-11, -9.4697410776597844e-11, 
    -9.4308458504060611e-11, -9.3923012383453368e-11, 
    -9.3552699416045912e-11, -9.3207293186978983e-11, 
    -9.2894473612047161e-11, -9.2619694150418856e-11, 
    -9.2386131906284256e-11, -9.2194748381305997e-11, 
    -9.2044441779336574e-11, -9.193228745555201e-11, -9.1853871555237067e-11, 
    -9.1803692764507097e-11, -9.177561891304246e-11, -9.1763371989069205e-11, 
    -9.1761007556274976e-11, -9.1763367809476246e-11, 
    -9.1766466004800748e-11, -9.1767785875656464e-11,
  // Sqw-F(7, 0-1999)
    0.022461199858423913, 0.022458902354948074, 0.022452032896436217, 
    0.022440657643187669, 0.022424877181850319, 0.022404813043979292, 
    0.022380590818404749, 0.022352321630514937, 0.022320083971389352, 
    0.022283907866738974, 0.022243763165561661, 0.022199553312190843, 
    0.022151115382781344, 0.022098226485634136, 0.022040615931654878, 
    0.021977981971535318, 0.021910011455810327, 0.021836400563436616, 
    0.021756874786882867, 0.021671206636534001, 0.021579229973816789, 
    0.021480850411451455, 0.021376051730237228, 0.021264898663805834, 
    0.021147536632803568, 0.021024189045531268, 0.020895152645255967, 
    0.020760791136014572, 0.020621527044142843, 0.020477831562313198, 
    0.020330212051128359, 0.020179196981764101, 0.020025318390019441, 
    0.019869092331706625, 0.019710998300876633, 0.019551458996877439, 
    0.019390822107132499, 0.019229345836262107, 0.019067189724012418, 
    0.018904411866170957, 0.018740973040581078, 0.018576747534449718, 
    0.018411539775321391, 0.018245105288140096, 0.018077174113824063, 
    0.01790747467410574, 0.017735756155610804, 0.017561807778311806, 
    0.017385473747468322, 0.017206663189180006, 0.017025354865417088, 
    0.016841596897449528, 0.016655502061824465, 0.016467239448921554, 
    0.016277023398819729, 0.016085100673124113, 0.015891736808576876, 
    0.015697202549145389, 0.015501761180218166, 0.015305657495064221, 
    0.015109109006726717, 0.014912299872634741, 0.014715377821409069, 
    0.014518454164679917, 0.014321606752087251, 0.014124885503019382, 
    0.01392831994656904, 0.013731928044692417, 0.0135357254819406, 
    0.013339734590332292, 0.013143992142225639, 0.012948555379525209, 
    0.012753505837337028, 0.012558950741124874, 0.012365021982725332, 
    0.012171872887790612, 0.01197967315566678, 0.011788602470046899, 
    0.011598843340929777, 0.011410573749200542, 0.011223960133930452, 
    0.011039151201391404, 0.010856272955356773, 0.010675425258886, 
    0.010496680142247633, 0.010320081969361478, 0.010145649463089428, 
    0.009973379465279977, 0.0098032521716835182, 0.0096352374417489235, 
    0.0094693016527368414, 0.0093054144659197348, 0.0091435548214730579, 
    0.0089837154971103977, 0.0088259056652099932, 0.0086701510641764897, 
    0.0085164916484596221, 0.008364976871316045, 0.0082156590486031893, 
    0.0080685855099898868, 0.0079237904277825247, 0.0077812872939203928, 
    0.0076410629774782074, 0.0075030741398686091, 0.0073672465310891042, 
    0.0072334773697504667, 0.0071016406629268594, 0.0069715949924032423, 
    0.0068431930214601115, 0.0067162917920178464, 0.0065907628045419825, 
    0.0064665009075086767, 0.0063434311608964664, 0.0062215130592049306, 
    0.0061007417759037187, 0.0059811463907985902, 0.0058627853521179786, 
    0.0057457396770211402, 0.0056301045846442431, 0.0055159803696293898, 
    0.0054034633550173834, 0.0052926377137852126, 0.0051835688281852898, 
    0.005076298681393485, 0.0049708435666760593, 0.0048671941768507225, 
    0.0047653179222136811, 0.0046651631369237952, 0.0045666646868824995, 
    0.00446975039658273, 0.0043743476733328866, 0.0042803897248284749, 
    0.0041878208357391863, 0.0040966002823040592, 0.0040067046091271418, 
    0.0039181281554100398, 0.0038308818834924489, 0.0037449907155847366, 
    0.0036604897111052882, 0.0035774195059320164, 0.0034958214788704863, 
    0.0034157331072133816, 0.0033371839249791021, 0.0032601924116500559, 
    0.0031847640272368929, 0.0031108904849506671, 0.0030385502299437564, 
    0.0029677099845107952, 0.0028983271369726346, 0.0028303526993758393, 
    0.0027637345398657427, 0.0026984206067025545, 0.0026343618966181517, 
    0.0025715149727305606, 0.0025098438980411392, 0.0024493215117839012, 
    0.0023899300313418139, 0.0023316610080546508, 0.0022745146992609469, 
    0.0022184989415977526, 0.0021636276236148932, 0.0021099188616053601, 
    0.0020573929837685752, 0.0020060704265502443, 0.0019559696446173375, 
    0.0019071051329216677, 0.001859485655338037, 0.0018131127684761572, 
    0.0017679797201755681, 0.0017240707886533528, 0.0016813611094014572, 
    0.0016398170125130288, 0.0015993968638034946, 0.0015600523704857531, 
    0.0015217302787303973, 0.0014843743593197204, 0.0014479275521921383, 
    0.0014123341242047002, 0.0013775416894734689, 0.0013435029496457016, 
    0.0013101770324584273, 0.0012775303394752925, 0.0012455368550809071, 
    0.001214177914678341, 0.0011834414759945024, 0.0011533209788268609, 
    0.0011238139113512982, 0.0010949202221415986, 0.0010666407245239124, 
    0.0010389756334731636, 0.0010119233560417571, 0.00098547962662888641, 
    0.00095963704150700524, 0.00093438500674030507, 0.00090971007392650781, 
    0.00088559660281495789, 0.00086202766197313843, 0.00083898606062623603, 
    0.00081645539787897304, 0.00079442101992837895, 0.00077287079065963416, 
    0.00075179560427357495, 0.0007311895976392529, 0.00071105005174518406, 
    0.0006913770026451807, 0.00067217260958352273, 0.00065344034898525793, 
    0.00063518411593658033, 0.00061740731880761772, 0.00060011204791958071, 
    0.00058329838667795907, 0.0005669639152002438, 0.00055110343450276889, 
    0.00053570891637288987, 0.00052076966267492755, 0.00050627264021784444, 
    0.00049220294505167251, 0.00047854434400876051, 0.00046527984148300912, 
    0.00045239222508222849, 0.00043986455349054044, 0.00042768056184133626, 
    0.00041582497221819768, 0.00040428370786296694, 0.0003930440180137346, 
    0.00038209452538227862, 0.00037142521013421449, 0.00036102734347702182, 
    0.00035089338161475284, 0.00034101682807625229, 0.00033139207032861984, 
    0.00032201419587112051, 0.00031287879389682138, 0.00030398175082620827, 
    0.000295319050843224, 0.00028688659504128846, 0.00027868005394276742, 
    0.00027069476724803792, 0.00026292570136542668, 0.00025536746974859814, 
    0.00024801441399151106, 0.00024086073605064794, 0.00023390066510294892, 
    0.00022712863757614598, 0.00022053946669338108, 0.00021412847890009924, 
    0.00020789159870051116, 0.00020182537013190769, 0.00019592691135610473, 
    0.00019019380744350416, 0.00018462395414717818, 0.00017921537128316145, 
    0.0001739660075506027, 0.0001688735589635461, 0.00016393532066213745, 
    0.00015914808722275345, 0.00015450811043244328, 0.00015001111668958226, 
    0.00014565237957853928, 0.00014142683746928329, 0.00013732924175509351, 
    0.00013335431889752226, 0.0001294969289165392, 0.00012575220427768483, 
    0.00012211565605313877, 0.00011858323841040807, 0.00011515136744939916, 
    0.00011181689564266369, 0.00010857704808079348, 0.00010542933085342465, 
    0.00010237142474198408, 9.9401078631273333e-05, 9.6516016505938525e-05, 
    9.3713869644850356e-05, 9.0992141938355152e-05, 8.8348211607993852e-05, 
    8.5779367617641115e-05, 8.3282874400021864e-05, 8.0856054807143957e-05, 
    7.8496378918787245e-05, 7.6201545785749058e-05, 7.3969546373309575e-05, 
    7.1798698680554024e-05, 6.9687649813145172e-05, 6.7635344113758456e-05, 
    6.5640960700991756e-05, 6.3703827378407631e-05, 6.1823320430730676e-05, 
    5.9998761083636351e-05, 5.82293193304931e-05, 5.6513934565893267e-05, 
    5.4851260295801535e-05, 5.3239637474028157e-05, 5.1677098116922641e-05, 
    5.0161398097465532e-05, 4.8690075663217279e-05, 4.7260530404738683e-05, 
    4.587011617731456e-05, 4.4516240828294121e-05, 4.3196465443833551e-05, 
    4.1908596123551319e-05, 4.0650761951958002e-05, 3.9421473808909758e-05, 
    3.8219659915805054e-05, 3.7044675519550765e-05, 3.5896285834149301e-05, 
    3.4774623220206008e-05, 3.3680121481159031e-05, 3.2613431945461022e-05, 
    3.1575327517348706e-05, 3.0566601938748119e-05, 2.9587971962840907e-05, 
    2.8639989897843784e-05, 2.7722973021092965e-05, 2.6836954758921949e-05, 
    2.5981660439941543e-05, 2.5156508088650842e-05, 2.4360632407135046e-05, 
    2.3592928066537449e-05, 2.2852106931621263e-05, 2.2136763026208453e-05, 
    2.1445438973857619e-05, 2.0776688266874648e-05, 2.0129128886639581e-05, 
    1.9501485307758087e-05, 1.8892617529688624e-05, 1.8301537262645414e-05, 
    1.772741257066246e-05, 1.7169563034988699e-05, 1.6627447822649289e-05, 
    1.6100648979255049e-05, 1.5588851923240053e-05, 1.5091824637118624e-05, 
    1.4609396566981739e-05, 1.4141437858788595e-05, 1.3687839339598e-05, 
    1.3248493598935533e-05, 1.2823277602010216e-05, 1.2412037401039396e-05, 
    1.201457562510992e-05, 1.1630642452130549e-05, 1.1259930657939609e-05, 
    1.0902075089296612e-05, 1.0556656550240927e-05, 1.0223209680394746e-05, 
    9.9012340120594798e-06, 9.5902070885162585e-06, 9.2895983640039535e-06, 
    8.9988826116152831e-06, 8.7175517365950995e-06, 8.4451241940829348e-06, 
    8.1811515893203065e-06, 7.9252224280464771e-06, 7.6769633245074226e-06, 
    7.436038213857216e-06, 7.2021462295691976e-06, 6.975018891241596e-06, 
    6.7544171270640324e-06, 6.5401284650075874e-06, 6.3319645163547807e-06, 
    6.129758688422042e-06, 5.9333639373383615e-06, 5.742650324873024e-06, 
    5.5575021781706134e-06, 5.377814750795579e-06, 5.2034904217748743e-06, 
    5.0344346109817785e-06, 4.8705517042713882e-06, 4.7117413445660528e-06, 
    4.5578954448112712e-06, 4.4088962152592071e-06, 4.2646153855621927e-06, 
    4.1249146620487765e-06, 3.9896473192002455e-06, 3.8586607039209462e-06, 
    3.7317993509847325e-06, 3.6089083750199687e-06, 3.4898368190853897e-06, 
    3.3744406912064509e-06, 3.2625854943916278e-06, 3.1541481343861017e-06, 
    3.0490181593111731e-06, 2.9470983352986796e-06, 2.84830459059823e-06, 
    2.7525653694662236e-06, 2.6598204360759242e-06, 2.5700191662068711e-06, 
    2.4831183713387046e-06, 2.3990797194107299e-06, 2.3178668505780082e-06, 
    2.2394423278809554e-06, 2.1637646042665158e-06, 2.090785216471047e-06, 
    2.0204464251475331e-06, 1.9526795021150647e-06, 1.8874038207256838e-06, 
    1.8245268379945614e-06, 1.7639449781728852e-06, 1.7055453474748912e-06, 
    1.6492081417731287e-06, 1.5948095608111691e-06, 1.5422250197417849e-06, 
    1.4913324496507814e-06, 1.4420154995526665e-06, 1.3941664836051089e-06, 
    1.3476889519162104e-06, 1.3024997924075375e-06, 1.258530792279735e-06, 
    1.2157295991022646e-06, 1.1740600285400669e-06, 1.1335016727614394e-06, 
    1.0940487788902572e-06, 1.055708393933292e-06, 1.0184978149367185e-06, 
    9.8244143703434229e-07, 9.4756715280680608e-07, 9.1390251334286979e-07, 
    8.8147090603058474e-07, 8.5028802564389582e-07, 8.2035890925591516e-07, 
    7.9167576857922416e-07, 7.6421679021824031e-07, 7.3794599072520158e-07, 
    7.1281412129084079e-07, 6.8876052620322198e-07, 6.6571578193575923e-07, 
    6.4360488659080337e-07, 6.223507384037681e-07, 6.018776364015727e-07, 
    5.8211455484619403e-07, 5.6299797921611794e-07, 5.4447414020011136e-07, 
    5.2650053566744692e-07, 5.0904668488204596e-07, 4.9209410908296702e-07, 
    4.756355771854713e-07, 4.5967369259962382e-07, 4.4421892864440183e-07, 
    4.2928724461373033e-07, 4.1489743391196215e-07, 4.0106836806537219e-07, 
    3.878163062053132e-07, 3.7515243624761596e-07, 3.6308080165395691e-07, 
    3.5159674443077707e-07, 3.4068596262318769e-07, 3.3032423931587043e-07, 
    3.2047785425512147e-07, 3.1110464105450718e-07, 3.0215560813199066e-07, 
    2.935770027963008e-07, 2.8531267002112426e-07, 2.773065412752958e-07, 
    2.6950508650282485e-07, 2.6185957200241534e-07, 2.5432798813160487e-07, 
    2.4687653938986432e-07, 2.3948062385860692e-07, 2.3212526480052261e-07, 
    2.2480499322712448e-07, 2.1752321288189442e-07, 2.1029110833176513e-07, 
    2.0312618039669343e-07, 1.9605051169123446e-07, 1.8908887690096359e-07, 
    1.8226681864211781e-07, 1.7560880852264367e-07, 1.6913660570756729e-07, 
    1.6286791024079568e-07, 1.5681538754305566e-07, 1.5098611329886667e-07, 
    1.4538145741041064e-07, 1.3999739265672619e-07, 1.3482518223955896e-07, 
    1.2985237204981897e-07, 1.2506399232610891e-07, 1.204438602128667e-07, 
    1.1597587207014458e-07, 1.116451810353334e-07, 1.0743917172438439e-07, 
    1.0334816641955648e-07, 9.9365824667102584e-08, 9.5489226214823306e-08, 
    9.1718654423935296e-08, 8.805711982561617e-08, 8.4509681205740929e-08, 
    8.1082632272594248e-08, 7.7782626892205144e-08, 7.4615814354318817e-08, 
    7.1587050386866814e-08, 6.8699239406379904e-08, 6.5952851295867573e-08, 
    6.3345641392826973e-08, 6.0872587559483449e-08, 5.8526042540962897e-08, 
    5.629608531950728e-08, 5.4171041191923226e-08, 5.2138128895326161e-08, 
    5.0184183778375213e-08, 4.8296400796618704e-08, 4.6463039405292672e-08, 
    4.4674035942387961e-08, 4.2921476456778462e-08, 4.1199895132682392e-08, 
    3.9506378199351366e-08, 3.7840470505139187e-08, 3.6203898766037961e-08, 
    3.4600141527823705e-08, 3.3033888107271879e-08, 3.1510437353467192e-08, 
    3.0035089792630095e-08, 2.8612584870298774e-08, 2.7246627722833379e-08, 
    2.5939539525942912e-08, 2.4692051987057076e-08, 2.3503252940684093e-08, 
    2.2370676290562041e-08, 2.1290518403600069e-08, 2.0257953977836927e-08, 
    1.9267519094146663e-08, 1.831352649893706e-08, 1.7390478949556858e-08, 
    1.6493449089654178e-08, 1.5618399315102314e-08, 1.4762420707739876e-08, 
    1.3923877072476192e-08, 1.3102446768509681e-08, 1.2299062382789093e-08, 
    1.15157548889986e-08, 1.0755415722557746e-08, 1.0021495768889291e-08, 
    9.3176653032956053e-09, 8.6474619417100543e-09, 8.0139552894006272e-09, 
    7.4194556836697935e-09, 6.865291260269171e-09, 6.3516713668363149e-09, 
    5.8776467668914215e-09, 5.4411676767531363e-09, 5.0392316136446584e-09, 
    4.6681042315482096e-09, 4.3235900122835225e-09, 4.0013254412309062e-09, 
    3.6970668732545403e-09, 3.4069472936829516e-09, 3.1276815107547018e-09, 
    2.8567058781257866e-09, 2.5922466537185398e-09, 2.3333182928404026e-09, 
    2.0796595612879594e-09, 1.8316197121566287e-09, 1.5900097823476168e-09, 
    1.3559344137409329e-09, 1.1306189012900509e-09, 9.1524391534605298e-10, 
    7.1079808355878121e-10, 5.179558573787638e-10, 3.369861364736984e-10, 
    1.6769499808116047e-10, 9.4046085535232973e-12, -1.3903128424465674e-10, 
    -2.7917614606072059e-10, -4.1292660553904922e-10, 
    -5.4240022798919259e-10, -6.6980220090175734e-10, 
    -7.9727981761450436e-10, -9.2677552369057516e-10, 
    -1.0598899520733302e-09, -1.1977664044995922e-09, 
    -1.3410067084738192e-09, -1.4896262225768095e-09, 
    -1.6430522288088041e-09, -1.8001663670299108e-09, 
    -1.9593876215314326e-09, -2.1187890327856241e-09, 
    -2.2762382995117176e-09, -2.4295508273027563e-09, 
    -2.5766429826834731e-09, -2.7156740399815607e-09, 
    -2.8451665999249079e-09, -2.9640977358506544e-09, 
    -3.0719555668169277e-09, -3.1687589839927617e-09, 
    -3.2550406431557485e-09, -3.3317959339169271e-09, 
    -3.4004022763182623e-09, -3.4625148420413481e-09, 
    -3.5199456415563598e-09, -3.5745339047884444e-09, 
    -3.6280159087274515e-09, -3.6819027497276213e-09, 
    -3.7373740929953882e-09, -3.7951954637466082e-09, 
    -3.8556651589725595e-09, -3.9185952972577013e-09, 
    -3.9833289231279879e-09, -4.0487925752440415e-09, 
    -4.1135805911990687e-09, -4.1760649001089584e-09, 
    -4.2345215322439478e-09, -4.287263811802885e-09, -4.3327714241146803e-09, 
    -4.3698053099991673e-09, -4.3974995938596655e-09, 
    -4.4154242809321135e-09, -4.4236149658016967e-09, 
    -4.4225689419265196e-09, -4.4132095903815382e-09, 
    -4.3968234247650865e-09, -4.3749756009200597e-09, 
    -4.3494109110639626e-09, -4.3219474181186042e-09, 
    -4.2943699331018994e-09, -4.2683296984392109e-09, 
    -4.2452560655495561e-09, -4.2262846975594986e-09, 
    -4.2122060051725236e-09, -4.2034360759102925e-09, 
    -4.2000114389702032e-09, -4.2016074281837656e-09, 
    -4.2075787833974405e-09, -4.2170195324484287e-09, 
    -4.2288380780650767e-09, -4.2418420282820795e-09, 
    -4.2548267097408401e-09, -4.2666606844905956e-09, 
    -4.2763619688133778e-09, -4.2831591593612821e-09, 
    -4.2865331968937621e-09, -4.2862370148635006e-09, 
    -4.2822925175708056e-09, -4.2749661578603799e-09, 
    -4.2647264333753134e-09, -4.2521878404379949e-09, 
    -4.2380469292776315e-09, -4.2230161767487696e-09, 
    -4.2077612784543914e-09, -4.1928464534453774e-09, 
    -4.1786914531723359e-09, -4.1655424195659776e-09, 
    -4.1534577215360595e-09, -4.142308534859152e-09, -4.1317932287747428e-09, 
    -4.1214637716620925e-09, -4.1107620778116161e-09, 
    -4.0990637141924188e-09, -4.0857263628045522e-09, 
    -4.0701400306155528e-09, -4.0517761017038203e-09, 
    -4.0302320140455308e-09, -4.0052686413635071e-09, 
    -3.9768375112295783e-09, -3.9450957072000603e-09, 
    -3.9104068228034171e-09, -3.8733275606203716e-09, 
    -3.8345804693771363e-09, -3.7950146999552478e-09, 
    -3.7555574606572248e-09, -3.7171599109493227e-09, 
    -3.6807414967434155e-09, -3.6471370064542618e-09, 
    -3.6170501336270559e-09, -3.59101682612713e-09, -3.5693806547635071e-09, 
    -3.552281452937309e-09, -3.5396572679536691e-09, -3.5312587760682621e-09, 
    -3.5266742754066196e-09, -3.5253629406221599e-09, 
    -3.5266934546837992e-09, -3.5299852041121967e-09, -3.534549117236094e-09, 
    -3.5397257175181415e-09, -3.5449182059174665e-09, 
    -3.5496190304408046e-09, -3.5534288024096055e-09, 
    -3.5560671052507109e-09, -3.5573750910818127e-09, 
    -3.5573104134651361e-09, -3.5559352730150848e-09, 
    -3.5533988702855732e-09, -3.5499156775299653e-09, 
    -3.5457412917606791e-09, -3.5411475191760835e-09, 
    -3.5363985019750338e-09, -3.5317293874460188e-09, 
    -3.5273289161038095e-09, -3.5233267937918291e-09, 
    -3.5197864605603432e-09, -3.5167032094081685e-09, 
    -3.5140073742112758e-09, -3.5115717522579159e-09, 
    -3.5092223418159817e-09, -3.5067511725994219e-09, 
    -3.5039301633650814e-09, -3.5005249154980495e-09, -3.496307690615121e-09, 
    -3.4910688795693313e-09, -3.484626682059412e-09, -3.4768347145895049e-09, 
    -3.4675875671077743e-09, -3.4568242182156071e-09, -3.444529426744828e-09, 
    -3.4307330360281117e-09, -3.4155073344395857e-09, -3.398962473390448e-09, 
    -3.381240191995342e-09, -3.3625060811134981e-09, -3.3429408619638407e-09, 
    -3.3227311361820369e-09, -3.3020603071249047e-09, 
    -3.2811001768002252e-09, -3.2600038891386106e-09, 
    -3.2389005504143226e-09, -3.217891908609284e-09, -3.1970510869857542e-09, 
    -3.1764233618003947e-09, -3.1560286931865752e-09, 
    -3.1358657454576396e-09, -3.1159169331834152e-09, 
    -3.0961541651040665e-09, -3.0765448331663498e-09, 
    -3.0570577746787039e-09, -3.0376687725495948e-09, -3.018365399603651e-09, 
    -2.9991508049345854e-09, -2.9800462771839701e-09, 
    -2.9610922314480839e-09, -2.9423475286876832e-09, 
    -2.9238869364319121e-09, -2.9057968431738126e-09, 
    -2.8881693372510401e-09, -2.871095093688618e-09, -2.8546555171742601e-09, 
    -2.8389149114390352e-09, -2.8239133090925598e-09, 
    -2.8096608152296981e-09, -2.796133997221351e-09, -2.7832748762210666e-09, 
    -2.7709926453519036e-09, -2.7591681263210078e-09, 
    -2.7476605238873124e-09, -2.7363159548079653e-09, 
    -2.7249769155063067e-09, -2.7134919203249573e-09, 
    -2.7017244096533986e-09, -2.689560312671974e-09, -2.6769136780142225e-09, 
    -2.6637301536027019e-09, -2.6499881786517349e-09, 
    -2.6356981084512854e-09, -2.6208994837641194e-09, -2.605656916178085e-09, 
    -2.5900549235884528e-09, -2.5741922149941599e-09, 
    -2.5581757050281768e-09, -2.5421146337470659e-09, 
    -2.5261149686491786e-09, -2.5102743595072909e-09, 
    -2.4946777190014277e-09, -2.4793936807010119e-09, 
    -2.4644719611260314e-09, -2.4499418533500675e-09, 
    -2.4358118498041264e-09, -2.4220705344364345e-09, 
    -2.4086886522139823e-09, -2.3956223414420464e-09, 
    -2.3828172575616441e-09, -2.3702133915164481e-09, -2.357750143138587e-09, 
    -2.3453713498015235e-09, -2.3330297328763754e-09, 
    -2.3206904968051401e-09, -2.3083336677463899e-09, 
    -2.2959550625870031e-09, -2.283565741951682e-09, -2.271190106959453e-09, 
    -2.2588627703997664e-09, -2.2466246229530635e-09, 
    -2.2345183984878863e-09, -2.2225842581566391e-09, 
    -2.2108557285821646e-09, -2.1993564259173448e-09, 
    -2.1880977691771713e-09, -2.1770778926248823e-09, 
    -2.1662817751803496e-09, -2.1556825447312046e-09, 
    -2.1452437627096143e-09, -2.1349225298970741e-09, 
    -2.1246730293866877e-09, -2.1144502904143916e-09, 
    -2.1042137804040657e-09, -2.0939306046112827e-09, -2.083577975209118e-09, 
    -2.0731448417553912e-09, -2.062632473891522e-09, -2.0520540544655902e-09, 
    -2.0414332403232163e-09, -2.0308019179437993e-09, 
    -2.0201972863088263e-09, -2.0096585956267638e-09, -1.999223756405082e-09, 
    -1.9889261597685019e-09, -1.9787918858063567e-09, -1.968837555946546e-09, 
    -1.9590688708394693e-09, -1.9494799727970701e-09, 
    -1.9400535211138087e-09, -1.9307615070956559e-09, 
    -1.9215666230892754e-09, -1.9124241441987462e-09, 
    -1.9032841362814388e-09, -1.8940939421823864e-09, 
    -1.8848007787669857e-09, -1.8753544262281915e-09, 
    -1.8657098415112899e-09, -1.8558296930355854e-09, 
    -1.8456866281179901e-09, -1.8352652490417948e-09, 
    -1.8245636085905613e-09, -1.813594174206387e-09, -1.8023840920386046e-09, 
    -1.7909747313997317e-09, -1.7794204028398591e-09, 
    -1.7677863356770672e-09, -1.7561458859452964e-09, 
    -1.7445772011882577e-09, -1.7331594416203168e-09, 
    -1.7219688521059554e-09, -1.7110748902814925e-09, 
    -1.7005367381692842e-09, -1.6904003783076072e-09, -1.680696538865763e-09, 
    -1.671439574328683e-09, -1.6626274608194553e-09, -1.6542428212738567e-09, 
    -1.6462549853986872e-09, -1.6386228461565698e-09, 
    -1.6312983417435083e-09, -1.6242302350689339e-09, 
    -1.6173679377032192e-09, -1.6106650071474944e-09, 
    -1.6040821016128642e-09, -1.5975890930620325e-09, 
    -1.5911662610202329e-09, -1.5848044068482305e-09, 
    -1.5785039902062764e-09, -1.5722733307681976e-09, 
    -1.5661261479678714e-09, -1.5600786191783004e-09, 
    -1.5541463227286554e-09, -1.5483413157632795e-09, 
    -1.5426697012988976e-09, -1.5371298472211293e-09, 
    -1.5317115141651646e-09, -1.5263958927776104e-09, 
    -1.5211566221189596e-09, -1.5159616199963699e-09, 
    -1.5107756207918997e-09, -1.5055631118372104e-09, 
    -1.5002914547971838e-09, -1.4949338424338574e-09, 
    -1.4894718825363408e-09, -1.4838974887181672e-09, 
    -1.4782139784048903e-09, -1.4724361916152111e-09, 
    -1.4665896843063796e-09, -1.4607089666974338e-09, 
    -1.4548350171154227e-09, -1.4490121756823076e-09, 
    -1.4432847603804174e-09, -1.4376936005034944e-09, 
    -1.4322728273367529e-09, -1.4270471248748375e-09, 
    -1.4220297025092958e-09, -1.4172210826473519e-09, 
    -1.4126088396219943e-09, -1.4081682421582723e-09, -1.403863780564375e-09, 
    -1.3996513863706084e-09, -1.3954812204149635e-09, 
    -1.3913007368065583e-09, -1.3870578515094918e-09, -1.382703906393713e-09, 
    -1.3781962739447104e-09, -1.3735003654927436e-09, 
    -1.3685909894392824e-09, -1.3634529218413233e-09, 
    -1.3580807701261668e-09, -1.3524781448612663e-09, 
    -1.3466563366532361e-09, -1.3406325950916556e-09, 
    -1.3344282845381867e-09, -1.3280670373210761e-09, 
    -1.3215731366064745e-09, -1.3149701973639211e-09, 
    -1.3082803090227931e-09, -1.3015235584175611e-09, 
    -1.2947179966538253e-09, -1.2878798873338573e-09, 
    -1.2810242167809855e-09, -1.2741652520904282e-09, 
    -1.2673171178683408e-09, -1.2604942187480678e-09, 
    -1.2537115148596475e-09, -1.2469845397714551e-09, -1.240329241023242e-09, 
    -1.2337616028587825e-09, -1.2272971772876185e-09, 
    -1.2209505235586665e-09, -1.2147346823288347e-09, 
    -1.2086606893008161e-09, -1.2027372370316672e-09, 
    -1.1969704369147699e-09, -1.1913637607070458e-09, -1.185918069659619e-09, 
    -1.180631770513536e-09, -1.1755009871280647e-09, -1.170519769208517e-09, 
    -1.1656802330403049e-09, -1.1609726700854096e-09, 
    -1.1563855447311908e-09, -1.1519054539268977e-09, 
    -1.1475169993381032e-09, -1.1432027015908143e-09, 
    -1.1389429081231555e-09, -1.1347158434186366e-09, 
    -1.1304977777200597e-09, -1.126263424859009e-09, -1.1219865243951977e-09, 
    -1.1176406947385898e-09, -1.1132004476009649e-09, 
    -1.1086423962814751e-09, -1.1039465216926784e-09, 
    -1.0990974624985519e-09, -1.0940856729838221e-09, 
    -1.0889083867378162e-09, -1.083570236429721e-09, -1.0780834985050509e-09, 
    -1.0724678416728551e-09, -1.0667496154256046e-09, 
    -1.0609606321802919e-09, -1.055136570712366e-09, -1.0493150282397616e-09, 
    -1.0435334242153126e-09, -1.0378268563626265e-09, 
    -1.0322261347131717e-09, -1.026756101977851e-09, -1.0214344389374606e-09, 
    -1.0162709963715774e-09, -1.0112677881017088e-09, 
    -1.0064195456674178e-09, -1.0017148888847199e-09, 
    -9.9713788644442229e-10, -9.9266994226771729e-10, 
    -9.8829176924958313e-10, -9.8398530549486628e-10, 
    -9.7973534867981823e-10, -9.7553082877575906e-10, 
    -9.7136553714031349e-10, -9.6723835098504343e-10, 
    -9.6315287647405448e-10, -9.5911664290323502e-10, 
    -9.5513987917137757e-10, -9.5123407619757502e-10, 
    -9.4741040478780562e-10, -9.4367820735618712e-10, 
    -9.4004363152848008e-10, -9.365085844589876e-10, -9.3307002314358644e-10, 
    -9.2971969236897852e-10, -9.2644426283231472e-10, 
    -9.2322591708769315e-10, -9.2004327230232411e-10, -9.168725927025884e-10, 
    -9.1368918945542604e-10, -9.1046891764031749e-10, 
    -9.0718960300525462e-10, -9.0383238506501324e-10, 
    -9.0038277668655168e-10, -8.9683147229859857e-10, 
    -8.9317477535508599e-10, -8.8941471665217017e-10, 
    -8.8555879616126997e-10, -8.8161945346170757e-10, 
    -8.7761327258797446e-10, -8.7356002598240327e-10, 
    -8.6948157095146041e-10, -8.6540073061551665e-10, 
    -8.6134013064681978e-10, -8.5732111828432858e-10, 
    -8.5336273523944482e-10, -8.4948085602380623e-10, 
    -8.4568745561266263e-10, -8.4199011592521123e-10, 
    -8.3839174340996815e-10, -8.3489059034206673e-10, 
    -8.3148053699888486e-10, -8.2815169187399997e-10, -8.2489123200537938e-10, 
    -8.2168447953740007e-10, -8.1851608568702077e-10, 
    -8.1537128473106971e-10, -8.1223704074095513e-10, 
    -8.0910305326807962e-10, -8.0596244596163325e-10, 
    -8.0281217275065511e-10, -7.9965299766634704e-10, 
    -7.9648916313884715e-10, -7.9332770789766373e-10, 
    -7.9017756139916116e-10, -7.8704848408488839e-10, 
    -7.8394999344676527e-10, -7.8089032993193968e-10, 
    -7.7787560958358445e-10, -7.7490916849136028e-10, 
    -7.7199120430327221e-10, -7.6911865664836668e-10, 
    -7.6628538625946134e-10, -7.6348254877662492e-10, 
    -7.6069918567415867e-10, -7.5792291910158144e-10, 
    -7.5514075006260968e-10, -7.5233986049057818e-10, 
    -7.4950841738749254e-10, -7.4663628693686782e-10, -7.437156904572727e-10, 
    -7.4074169884216747e-10, -7.3771261669466911e-10, 
    -7.3463017191229042e-10, -7.3149956524775117e-10, 
    -7.2832930930663822e-10, -7.251309265802738e-10, -7.2191844231183468e-10, 
    -7.1870776799148676e-10, -7.1551592099473116e-10, 
    -7.1236019489190492e-10, -7.0925725518836594e-10, 
    -7.0622227718278381e-10, -7.0326811735430654e-10, 
    -7.0040464551289933e-10, -6.9763822321253325e-10, 
    -6.9497143291119546e-10, -6.9240303312102841e-10, 
    -6.8992819050792097e-10, -6.87538930472104e-10, -6.852248170511767e-10, 
    -6.8297374381130424e-10, -6.8077282550019797e-10, 
    -6.7860925464660692e-10, -6.7647109199387434e-10, 
    -6.7434788550628059e-10, -6.7223111688885335e-10, 
    -6.7011439829056967e-10, -6.6799347358299211e-10, 
    -6.6586599958517633e-10, -6.6373119394820768e-10, 
    -6.6158935707788918e-10, -6.5944136825225324e-10, 
    -6.5728817203864714e-10, -6.5513034912406484e-10, 
    -6.5296775492106319e-10, -6.5079931764141539e-10, 
    -6.4862294394278218e-10, -6.4643559185893787e-10, 
    -6.4423345457343841e-10, -6.4201228754488742e-10, 
    -6.3976780547932035e-10, -6.3749615481199514e-10, 
    -6.3519440183662521e-10, -6.328610167270005e-10, -6.3049628970514419e-10, 
    -6.2810266015912524e-10, -6.2568490555817712e-10, 
    -6.2325019022940687e-10, -6.208079235694751e-10, -6.1836947083258667e-10, 
    -6.1594769065674292e-10, -6.1355636859814771e-10, 
    -6.1120955505106815e-10, -6.0892088762684616e-10, 
    -6.0670292715446137e-10, -6.0456658153230088e-10, 
    -6.0252063641788873e-10, -6.0057144314997639e-10, 
    -5.9872275442191174e-10, -5.9697572893519681e-10, 
    -5.9532904172861207e-10, -5.9377912575637015e-10, 
    -5.9232043016912321e-10, -5.9094571358408791e-10, 
    -5.8964628724306538e-10, -5.8841221953791747e-10, 
    -5.8723246172166875e-10, -5.860949202118519e-10, -5.8498648819435844e-10, 
    -5.8389308404298422e-10, -5.8279971315409938e-10, 
    -5.8169062924544646e-10, -5.805495804768898e-10, -5.79360186474401e-10, 
    -5.7810641347403534e-10, -5.7677314640270219e-10, 
    -5.7534678473923259e-10, -5.7381583813316199e-10, 
    -5.7217143171740196e-10, -5.7040771115016055e-10, 
    -5.6852206662148929e-10, -5.6651518987553434e-10, 
    -5.6439095046169359e-10, -5.6215612234223122e-10, 
    -5.5981998499171731e-10, -5.5739387870711421e-10, 
    -5.5489071813176672e-10, -5.5232454717519208e-10, 
    -5.4971012953612861e-10, -5.4706263241110131e-10, 
    -5.4439734855741054e-10, -5.4172948315933199e-10, 
    -5.3907394830949026e-10, -5.3644516893546026e-10, -5.338568483504848e-10, 
    -5.3132170311727874e-10, -5.2885115696059452e-10, 
    -5.2645503344979795e-10, -5.2414124448745188e-10, 
    -5.2191556413917649e-10, -5.1978147360057945e-10, 
    -5.1774015796940364e-10, -5.1579063996736989e-10, 
    -5.1393007309711125e-10, -5.1215414730557053e-10, 
    -5.1045759902274863e-10, -5.0883472847258408e-10, 
    -5.0727989176875943e-10, -5.0578788234668817e-10, 
    -5.0435417725999475e-10, -5.0297497551747396e-10, 
    -5.0164708658994532e-10, -5.0036762367929186e-10, 
    -4.9913361011719181e-10, -4.9794152516714643e-10, 
    -4.9678689627426338e-10, -4.9566398516166169e-10, 
    -4.9456566712595178e-10, -4.9348349764212354e-10, -4.924080113350301e-10, 
    -4.9132920010048285e-10, -4.9023713997212684e-10, 
    -4.8912267205610741e-10, -4.8797805490328886e-10, 
    -4.8679749151138792e-10, -4.8557748498344714e-10, 
    -4.8431692607252547e-10, -4.8301694892341162e-10, 
    -4.8168053344535916e-10, -4.8031192917253741e-10, 
    -4.7891595711673049e-10, -4.774973027451515e-10, -4.760598584410642e-10, 
    -4.7460622585012041e-10, -4.7313739976286932e-10, 
    -4.7165269854861727e-10, -4.7014990708798271e-10, 
    -4.6862562475000008e-10, -4.6707574697803769e-10, 
    -4.6549604893364361e-10, -4.6388275978159423e-10, 
    -4.6223310194333571e-10, -4.6054571688041926e-10, 
    -4.5882096225861817e-10, -4.5706103193403658e-10, 
    -4.5526993884853622e-10, -4.5345331597040063e-10, 
    -4.5161810194981908e-10, -4.4977210326793075e-10, 
    -4.4792348692495724e-10, -4.460802160642588e-10, -4.4424949074784602e-10, 
    -4.4243719323559288e-10, -4.4064742933968519e-10, 
    -4.3888214856996065e-10, -4.3714092737875347e-10, 
    -4.3542091110240496e-10, -4.3371696559533016e-10, 
    -4.3202200776946931e-10, -4.3032753905633985e-10, 
    -4.2862431148748502e-10, -4.269031146547841e-10, -4.2515558455548677e-10, 
    -4.2337499203053547e-10, -4.2155691738422176e-10, -4.196997795775811e-10, 
    -4.1780512953115056e-10, -4.1587773907201154e-10, 
    -4.1392542467774033e-10, -4.119586779740205e-10, -4.0999009444074464e-10, 
    -4.0803370266321425e-10, -4.0610420524987729e-10, 
    -4.0421623003024812e-10, -4.0238360987015261e-10, 
    -4.0061877477621754e-10, -3.9893222945107219e-10, 
    -3.9733218843410238e-10, -3.9582430813750127e-10, 
    -3.9441156902339965e-10, -3.9309422235220715e-10, 
    -3.9186985719217606e-10, -3.907334966996456e-10, -3.8967778383014462e-10, 
    -3.8869319098015818e-10, -3.8776829385044487e-10, 
    -3.8689008271260858e-10, -3.8604434637615326e-10, 
    -3.8521609068626941e-10, -3.8439002493210161e-10, 
    -3.8355106649869578e-10, -3.8268487985104208e-10, 
    -3.8177837966825003e-10, -3.8082022086156597e-10, 
    -3.7980118027949555e-10, -3.7871446853036137e-10, 
    -3.7755589049389164e-10, -3.7632390354352718e-10, 
    -3.7501951143249588e-10, -3.7364608069896029e-10, 
    -3.7220901790461691e-10, -3.707154124705784e-10, -3.6917360113690344e-10, 
    -3.6759274507162939e-10, -3.6598237790623874e-10, 
    -3.6435201205776134e-10, -3.6271074891301815e-10, 
    -3.6106696874189683e-10, -3.5942804630611208e-10, 
    -3.5780017277000332e-10, -3.5618821651103502e-10, 
    -3.5459569939251594e-10, -3.5302483654309035e-10, 
    -3.5147668379866867e-10, -3.4995134493449361e-10, 
    -3.4844827636499219e-10, -3.4696660211316496e-10, 
    -3.4550548034682355e-10, -3.4406441802341046e-10, 
    -3.4264357564109327e-10, -3.4124393809486514e-10, 
    -3.3986743437873456e-10, -3.385168866423298e-10, -3.3719586611089888e-10, 
    -3.3590840632933131e-10, -3.3465865776126011e-10, 
    -3.3345043874647744e-10, -3.3228681907644736e-10, 
    -3.3116967411594369e-10, -3.3009936530564007e-10, 
    -3.2907448286360993e-10, -3.2809177351941748e-10, 
    -3.2714619526145722e-10, -3.2623117521001638e-10, 
    -3.2533898591474255e-10, -3.2446128459949302e-10, 
    -3.2358969939469252e-10, -3.2271647413072495e-10, 
    -3.2183504264572946e-10, -3.2094054968408318e-10, 
    -3.2003017371437975e-10, -3.191033164177566e-10, -3.1816154729304291e-10, 
    -3.1720838247488319e-10, -3.1624887310890239e-10, 
    -3.1528910575256789e-10, -3.1433560720197189e-10, 
    -3.1339481422821504e-10, -3.1247256387105786e-10, 
    -3.1157375749441031e-10, -3.1070213932462419e-10, 
    -3.0986028496636237e-10, -3.0904969653715177e-10, 
    -3.0827105276811353e-10, -3.075244895308964e-10, -3.0680992915362719e-10, 
    -3.0612732705788721e-10, -3.054768818170411e-10, -3.048590954339808e-10, 
    -3.0427475524514491e-10, -3.0372478776549038e-10, 
    -3.0321007887512145e-10, -3.0273122485628205e-10, 
    -3.0228834347043021e-10, -3.0188089202178129e-10, 
    -3.0150760248318362e-10, -3.0116645896369236e-10, 
    -3.0085480787825373e-10, -3.0056946779702043e-10, 
    -3.0030691452561686e-10, -3.0006341438078031e-10, 
    -2.9983515902978701e-10, -2.9961830024644049e-10, 
    -2.9940897055033672e-10, -2.9920321475935539e-10, 
    -2.9899693956746056e-10, -2.9878583758439246e-10, 
    -2.9856540775981831e-10, -2.9833100701167096e-10, 
    -2.9807803222747035e-10, -2.9780214414467915e-10, -2.974995901184094e-10, 
    -2.9716749009931193e-10, -2.96804128326213e-10, -2.9640910408138967e-10, 
    -2.959833872777545e-10, -2.9552917097760469e-10, -2.9504959833413704e-10, 
    -2.9454830316161392e-10, -2.9402891294889684e-10, 
    -2.9349446832637048e-10, -2.9294691373038009e-10, 
    -2.9238665734240975e-10, -2.9181231215077925e-10, 
    -2.9122057105315142e-10, -2.9060631781458876e-10, 
    -2.8996286090646662e-10, -2.8928234408026973e-10, -2.885562186269309e-10, 
    -2.8777581305145766e-10, -2.8693286095528011e-10, 
    -2.8602004322234554e-10, -2.8503143205173058e-10, 
    -2.8396291233908444e-10, -2.828124694004546e-10, -2.8158043117177648e-10, 
    -2.8026958850032831e-10, -2.7888525954761987e-10, 
    -2.7743522671860757e-10, -2.7592962015829126e-10, 
    -2.7438066737738197e-10, -2.7280238398004107e-10, 
    -2.7121014311220537e-10, -2.6962019433609412e-10, -2.680490752737629e-10, 
    -2.6651302668179097e-10, -2.650273373123321e-10, -2.6360574345803784e-10, 
    -2.6225983682197802e-10, -2.609985892238143e-10, -2.5982795548815445e-10, 
    -2.5875067485481793e-10, -2.5776619779868323e-10, 
    -2.5687084803618102e-10, -2.56058135175933e-10, -2.553193036864557e-10, 
    -2.5464399170718917e-10, -2.5402102686622781e-10, 
    -2.5343924952880667e-10, -2.5288836164894022e-10, 
    -2.5235964796874622e-10, -2.5184656993695306e-10, 
    -2.5134512901229215e-10, -2.5085402694765487e-10, 
    -2.5037452519405665e-10, -2.4991011595536084e-10, -2.494659712901762e-10, 
    -2.4904829316736614e-10, -2.4866359711435009e-10, 
    -2.4831806600406387e-10, -2.4801698440507898e-10, 
    -2.4776437577356869e-10, -2.475628012449584e-10, -2.474133855427052e-10, 
    -2.4731596240631103e-10, -2.4726934996189392e-10, 
    -2.4727161141638829e-10, -2.4732028974423522e-10, 
    -2.4741249151069836e-10, -2.4754483776455407e-10, 
    -2.4771321403702623e-10, -2.4791242122436426e-10, 
    -2.4813571365299037e-10, -2.4837437628841124e-10, -2.486173744223939e-10, 
    -2.4885123841590727e-10, -2.4906016747406177e-10, 
    -2.4922646261087073e-10, -2.4933121275094626e-10, 
    -2.4935526510851488e-10, -2.4928030758261696e-10, 
    -2.4909005030092234e-10, -2.4877130629141028e-10, 
    -2.4831493406143156e-10, -2.477164946637395e-10, -2.4697662366047547e-10, 
    -2.4610103698365735e-10, -2.4510024626084888e-10, 
    -2.4398896896107957e-10, -2.4278535843605681e-10, 
    -2.4151007881208398e-10, -2.4018535399153936e-10, 
    -2.3883400427572034e-10, -2.3747859540419921e-10, -2.361406631321878e-10, 
    -2.3484008779780603e-10, -2.3359458655751525e-10, 
    -2.3241935677956836e-10, -2.3132680591385575e-10, 
    -2.3032640661206485e-10, -2.2942463331925855e-10, -2.28624994761392e-10, 
    -2.2792812659717229e-10, -2.2733200641546686e-10, 
    -2.2683220216559923e-10, -2.2642221913550092e-10, 
    -2.2609388264375039e-10, -2.2583777975598924e-10, 
    -2.2564368572545318e-10, -2.2550099621136205e-10, 
    -2.2539908176116002e-10, -2.2532759488797938e-10, 
    -2.2527665451986763e-10, -2.2523695332061475e-10, 
    -2.2519973534822589e-10, -2.2515673066970273e-10, 
    -2.2510001129645989e-10, -2.2502185532030879e-10, 
    -2.2491462922755783e-10, -2.2477076644622385e-10, 
    -2.2458282294016886e-10, -2.2434367224889262e-10, 
    -2.2404680261289099e-10, -2.2368672899857371e-10, 
    -2.2325944070689327e-10, -2.2276288704063301e-10, 
    -2.2219738795231222e-10, -2.2156594304116488e-10, 
    -2.2087437140276309e-10, -2.2013128071860161e-10, 
    -2.1934779019436772e-10, -2.1853707207918811e-10, 
    -2.1771369327827547e-10, -2.1689285527080923e-10, 
    -2.1608953767442867e-10, -2.1531765981696608e-10, 
    -2.1458929362541201e-10, -2.1391403050441127e-10, 
    -2.1329850262247771e-10, -2.1274613512595325e-10, 
    -2.1225710352437516e-10, -2.1182852868073021e-10, 
    -2.1145484230834809e-10, -2.1112832767602328e-10, 
    -2.1083973360855961e-10, -2.1057895326999844e-10, 
    -2.1033565790564421e-10, -2.1009987905563828e-10, 
    -2.0986244031448621e-10, -2.0961525096348432e-10, 
    -2.0935141404258161e-10, -2.0906518093804056e-10, 
    -2.0875175868332571e-10, -2.0840704138292181e-10, 
    -2.0802728939257768e-10, -2.0760887476186046e-10, 
    -2.0714808561530293e-10, -2.0664109983908818e-10, 
    -2.0608409373713588e-10, -2.054735498660667e-10, -2.0480665694716623e-10, 
    -2.0408181574822178e-10, -2.0329912175413045e-10, 
    -2.0246079698329812e-10, -2.0157144957054151e-10, 
    -2.0063814531851825e-10, -1.9967023377574253e-10, 
    -1.9867895664372425e-10, -1.9767685062592332e-10, 
    -1.9667702985577505e-10, -1.9569239267781853e-10, 
    -1.9473488402541144e-10, -1.9381483445256883e-10, -1.929404823904373e-10, 
    -1.9211767661608012e-10, -1.9134980298873999e-10, 
    -1.9063787972580035e-10, -1.8998082421486552e-10, 
    -1.8937580607777397e-10, -1.8881866605532703e-10, 
    -1.8830431550603772e-10, -1.8782713706882531e-10, 
    -1.8738128776350076e-10, -1.8696095523688308e-10, 
    -1.8656051956341355e-10, -1.8617467422625723e-10, 
    -1.8579846843015769e-10, -1.8542731940971862e-10, 
    -1.8505699322537166e-10, -1.8468356930754804e-10, -1.843033849396988e-10, 
    -1.8391301309173871e-10, -1.8350922378566301e-10, 
    -1.8308898612683463e-10, -1.8264949651873236e-10, 
    -1.8218826194316911e-10, -1.8170320022604643e-10, 
    -1.8119280495438511e-10, -1.8065630230059994e-10, 
    -1.8009383683995211e-10, -1.7950660412867884e-10, 
    -1.7889695819288018e-10, -1.7826841734622565e-10, 
    -1.7762559077576794e-10, -1.7697399126620988e-10, 
    -1.7631975905832741e-10, -1.7566929581870068e-10, 
    -1.7502886714871548e-10, -1.7440417101359949e-10, 
    -1.7379995137486806e-10, -1.732196632239943e-10, -1.7266523647221128e-10, 
    -1.7213694323545444e-10, -1.7163339638378717e-10, 
    -1.7115164785205277e-10, -1.7068738794971292e-10, 
    -1.7023520801698246e-10, -1.6978892012895744e-10, 
    -1.6934187363650338e-10, -1.6888727454692281e-10, 
    -1.6841846124837862e-10, -1.6792915179805526e-10, -1.674136200000429e-10, 
    -1.6686685034552135e-10, -1.6628462616878831e-10, 
    -1.6566360946519072e-10, -1.6500139479883801e-10, 
    -1.6429654926362157e-10, -1.6354865962532003e-10, -1.627583946280486e-10, 
    -1.6192754501765498e-10, -1.610590802346579e-10, -1.6015716260726772e-10, 
    -1.5922714637528882e-10, -1.5827550748403049e-10, -1.573097198198195e-10, 
    -1.5633804946962138e-10, -1.5536929255739845e-10, 
    -1.5441243860315553e-10, -1.5347630734487692e-10, -1.525691679436681e-10, 
    -1.5169838080783803e-10, -1.5087008189217042e-10, 
    -1.5008895990458398e-10, -1.4935811011368742e-10, 
    -1.4867900212228803e-10, -1.4805153691655895e-10, 
    -1.4747420411573405e-10, -1.4694429150206636e-10, 
    -1.4645815138507848e-10, -1.4601148861407244e-10, 
    -1.4559964800515026e-10, -1.4521790147647993e-10, 
    -1.4486172455602447e-10, -1.4452704353752657e-10, 
    -1.4421048624423815e-10, -1.4390959289945114e-10, 
    -1.4362301603896801e-10, -1.4335066935538731e-10, 
    -1.4309384418481682e-10, -1.4285523016928661e-10, 
    -1.4263885978617743e-10, -1.424499414957223e-10, -1.4229456889388141e-10, 
    -1.4217933030130466e-10, -1.4211082981547406e-10, 
    -1.4209514450310241e-10, -1.4213727579614205e-10, 
    -1.4224063336650539e-10, -1.4240662990905147e-10, -1.426343919380266e-10, 
    -1.4292065348906562e-10, -1.4325983338832031e-10, 
    -1.4364429569088176e-10, -1.440647702248519e-10, -1.4451088401988175e-10, 
    -1.4497176479411014e-10, -1.4543665041016367e-10, 
    -1.4589544576064798e-10, -1.4633918909956383e-10, 
    -1.4676037639354868e-10, -1.4715315255641598e-10, 
    -1.4751333754010856e-10, -1.4783833260536357e-10, 
    -1.4812690955329587e-10, -1.4837895252846116e-10, 
    -1.4859515776617087e-10, -1.487767499603257e-10, -1.4892524399765325e-10, 
    -1.4904225170975697e-10, -1.4912935711028452e-10, 
    -1.4918804935357286e-10, -1.4921968810776248e-10, -1.492254901960749e-10, 
    -1.4920651622867641e-10, -1.4916364460175098e-10, 
    -1.4909751764625397e-10, -1.490084910308521e-10, -1.4889656504556641e-10, 
    -1.4876135863716059e-10, -1.4860212260661322e-10, 
    -1.4841782391606999e-10, -1.4820731181663716e-10, 
    -1.4796956044035129e-10, -1.4770397335779747e-10, 
    -1.4741070886317574e-10, -1.4709098771885489e-10, 
    -1.4674734516522123e-10, -1.4638376660117768e-10, 
    -1.4600567719796324e-10, -1.4561977482573775e-10, 
    -1.4523371776756929e-10, -1.4485567207658639e-10, 
    -1.4449377102626252e-10, -1.4415555102304217e-10, 
    -1.4384741248409332e-10, -1.4357415948695601e-10, -1.433386916296279e-10, 
    -1.4314183517006015e-10, -1.4298235743657336e-10, 
    -1.4285714032697526e-10, -1.427614864466652e-10, -1.4268951858229663e-10, 
    -1.4263464085741946e-10, -1.4259000408773457e-10, 
    -1.4254893863097914e-10, -1.425053376078766e-10, -1.4245398733462241e-10, 
    -1.4239080705422608e-10, -1.4231303796403536e-10, 
    -1.4221936567416093e-10, -1.4211000210820937e-10, 
    -1.4198670996784609e-10, -1.4185278214591768e-10, 
    -1.4171295276271514e-10, -1.4157324283696578e-10, 
    -1.4144070632696486e-10, -1.4132308250718224e-10, 
    -1.4122834919945691e-10, -1.41164200473248e-10, -1.4113747175029969e-10, 
    -1.4115355916189914e-10, -1.4121588151911092e-10, 
    -1.4132546661485669e-10, -1.4148066729498924e-10, 
    -1.4167709932046831e-10, -1.4190777237723495e-10, 
    -1.4216345270612354e-10, -1.4243320352136534e-10, 
    -1.4270506729567397e-10, -1.42966825670852e-10, -1.4320678117321243e-10, 
    -1.4341445922472915e-10, -1.4358122221965006e-10, 
    -1.4370069425918105e-10, -1.4376901180888019e-10, 
    -1.4378488427458263e-10, -1.4374945130239006e-10, 
    -1.4366600014741669e-10, -1.4353955946900728e-10, 
    -1.4337640773573107e-10, -1.4318354447224038e-10, 
    -1.4296816108086969e-10, -1.4273714737404322e-10, 
    -1.4249664337269864e-10, -1.4225167812849685e-10, -1.420058930379966e-10, 
    -1.417613483111692e-10, -1.4151843527986881e-10, -1.4127589448086193e-10, 
    -1.4103090366304253e-10, -1.4077928115270552e-10, 
    -1.4051574342287882e-10, -1.4023424067645673e-10, 
    -1.3992833102602675e-10, -1.3959158203539837e-10, 
    -1.3921797179701911e-10, -1.3880227438936413e-10, 
    -1.3834038561862508e-10, -1.3782960433130776e-10, 
    -1.3726880786029885e-10, -1.3665856633019185e-10, -1.360011467651585e-10, 
    -1.353004413793365e-10, -1.345618185650174e-10, -1.3379191972773028e-10, 
    -1.3299840891593463e-10, -1.3218970250079433e-10, 
    -1.3137468521224704e-10, -1.3056243631416058e-10, 
    -1.2976196066100654e-10, -1.2898194781801695e-10, 
    -1.2823053995954242e-10, -1.2751513269067864e-10, 
    -1.2684218020700256e-10, -1.2621704004519451e-10, 
    -1.2564382310961734e-10, -1.2512528184700637e-10, 
    -1.2466272079272358e-10, -1.2425596445815227e-10, 
    -1.2390336686259741e-10, -1.2360187884854431e-10, 
    -1.2334718509393276e-10, -1.2313391183943543e-10, 
    -1.2295588851056365e-10, -1.2280646230246226e-10, 
    -1.2267884472776001e-10, -1.2256647097912903e-10, 
    -1.2246333694417977e-10, -1.2236429469892904e-10, 
    -1.2226527770622857e-10, -1.221634421507759e-10, -1.2205720278078117e-10, 
    -1.2194617251558441e-10, -1.2183100329018979e-10, 
    -1.2171315808605562e-10, -1.2159461945132704e-10, 
    -1.2147758896683699e-10, -1.2136417796851813e-10, 
    -1.2125615223976422e-10, -1.2115471958476865e-10, 
    -1.2106040959162368e-10, -1.2097302736287412e-10, 
    -1.2089170185095784e-10, -1.2081500963102459e-10, 
    -1.2074115812202178e-10, -1.2066821315906686e-10, 
    -1.2059435607623444e-10, -1.2051811732598969e-10, 
    -1.2043860338369287e-10, -1.203556578046483e-10, -1.2026996547889494e-10, 
    -1.2018307648926791e-10, -1.2009735464347335e-10, 
    -1.2001583466101104e-10, -1.1994202247057464e-10, 
    -1.1987961790472637e-10, -1.198322173630431e-10, -1.1980297688322665e-10, 
    -1.1979430258699122e-10, -1.1980756159582112e-10, 
    -1.1984285083672349e-10, -1.1989884625332927e-10, 
    -1.1997274421564007e-10, -1.2006030600661122e-10, 
    -1.2015601401794073e-10, -1.202533242165234e-10, -1.2034500779292512e-10, 
    -1.204235610419375e-10, -1.2048166206982045e-10, -1.2051263327923254e-10, 
    -1.2051088123363258e-10, -1.2047227484208476e-10, 
    -1.2039445309613903e-10, -1.2027699880425534e-10, 
    -1.2012149960124089e-10, -1.1993145926304939e-10, 
    -1.1971208056750825e-10, -1.1946992238556731e-10, 
    -1.1921247080649759e-10, -1.1894764297088485e-10, 
    -1.1868328066892194e-10, -1.1842665812535374e-10, -1.181840719188117e-10, 
    -1.1796052017585507e-10, -1.1775951725968877e-10, 
    -1.1758305551337412e-10, -1.1743169568164424e-10, 
    -1.1730478459346597e-10, -1.1720078949106764e-10, 
    -1.1711765783903534e-10, -1.1705321424469417e-10, 
    -1.1700551005696718e-10, -1.1697311405419373e-10, 
    -1.1695528161394835e-10, -1.1695202039968946e-10, 
    -1.1696401495267304e-10, -1.1699243822544547e-10, 
    -1.1703866797700634e-10, -1.1710395664270033e-10, 
    -1.1718906733871828e-10, -1.1729394016949201e-10, 
    -1.1741740290827704e-10, -1.1755698173646797e-10, 
    -1.1770879821153127e-10, -1.1786758153982326e-10, 
    -1.1802678769119614e-10, -1.1817880819377555e-10, 
    -1.1831526037555258e-10, -1.1842734858930719e-10, 
    -1.1850626406884242e-10, -1.1854362626975582e-10, 
    -1.1853194995309845e-10, -1.1846511504077244e-10, 
    -1.1833883399026324e-10, -1.181511173739805e-10, -1.1790267077575475e-10, 
    -1.1759722348500246e-10, -1.1724174629495393e-10, 
    -1.1684651335141717e-10, -1.1642497764953514e-10, 
    -1.1599342871813929e-10, -1.155704263729094e-10, -1.1517600466828935e-10, 
    -1.1483067636148781e-10, -1.1455430158828917e-10, 
    -1.1436485273873086e-10, -1.1427720098257402e-10, 
    -1.1430197677644863e-10, -1.1444461886880875e-10, 
    -1.1470468488417299e-10, -1.1507549047927447e-10, 
    -1.1554412954172722e-10, -1.1609188411280949e-10, 
    -1.1669502038009059e-10, -1.1732593271389707e-10, 
    -1.1795455499099427e-10, -1.1854997880902973e-10, -1.190821449896305e-10, 
    -1.1952349957212826e-10, -1.1985051513448077e-10, 
    -1.2004496437214915e-10, -1.2009484582684666e-10, 
    -1.1999492164118746e-10, -1.1974681323705093e-10, 
    -1.1935866678668535e-10, -1.1884441038455304e-10, 
    -1.1822267113101463e-10, -1.1751542940671027e-10, 
    -1.1674651549661264e-10, -1.1594005351104228e-10, 
    -1.1511897543171026e-10, -1.1430369561477299e-10, 
    -1.1351103553445292e-10, -1.127534802266037e-10, -1.1203878596314769e-10, 
    -1.1136997522078928e-10, -1.1074568465130302e-10, 
    -1.1016083777302124e-10, -1.0960757134002043e-10, 
    -1.0907632787381629e-10, -1.0855701879099128e-10, 
    -1.0804016145970518e-10, -1.0751788835925292e-10, 
    -1.0698475495796092e-10, -1.0643827397942455e-10, 
    -1.0587914977070168e-10, -1.0531120894491385e-10, 
    -1.0474103605841098e-10, -1.0417738389961695e-10, 
    -1.0363039761874383e-10, -1.0311077439634522e-10, 
    -1.0262890975010641e-10, -1.0219412008346415e-10, -1.018140207376988e-10, 
    -1.0149409764110999e-10, -1.0123748893471841e-10, 
    -1.0104499685909214e-10, -1.0091527596512347e-10, 
    -1.0084517948187569e-10, -1.0083018857375116e-10, 
    -1.0086486974818383e-10, -1.0094330277022204e-10, 
    -1.0105943656788651e-10, -1.0120733267175428e-10, 
    -1.0138130208532942e-10, -1.0157594241553924e-10, 
    -1.0178608664596822e-10, -1.0200672984522154e-10, 
    -1.0223294757842721e-10, -1.0245986005597854e-10, 
    -1.0268264376629859e-10, -1.0289661329698097e-10, 
    -1.0309737648235799e-10, -1.0328100684573439e-10, 
    -1.0344423381209665e-10, -1.0358460631338393e-10, 
    -1.0370060355424407e-10, -1.0379167833321139e-10, 
    -1.0385822797623889e-10, -1.0390150071117383e-10, 
    -1.0392346804750466e-10, -1.0392668072442098e-10, 
    -1.0391413498720389e-10, -1.0388917546899546e-10, 
    -1.0385545403707231e-10, -1.0381692743326067e-10, 
    -1.0377787821181476e-10, -1.0374295388858898e-10, 
    -1.0371718457010868e-10, -1.0370595040935444e-10, 
    -1.0371487649770498e-10, -1.0374964980080441e-10, 
    -1.0381576277141158e-10, -1.0391818623887038e-10, 
    -1.0406100793971189e-10, -1.0424706982936771e-10, 
    -1.0447763044137437e-10, -1.0475210036662223e-10, 
    -1.0506787806889087e-10, -1.0542030021543025e-10, 
    -1.0580271756363849e-10, -1.0620670339987201e-10, -1.066223749738588e-10, 
    -1.0703880363562487e-10, -1.0744449200449538e-10, -1.078278785038706e-10, 
    -1.081778403952921e-10, -1.0848415584318895e-10, -1.0873790194172985e-10, 
    -1.0893177343583273e-10, -1.0906027609373939e-10, 
    -1.0911983321301508e-10, -1.0910876902972505e-10, 
    -1.0902719478344025e-10, -1.0887680804563463e-10, 
    -1.0866063084315969e-10, -1.0838269546515384e-10, 
    -1.0804771798019918e-10, -1.076607767034087e-10, -1.0722701945455946e-10, 
    -1.0675141782006141e-10, -1.0623859144019027e-10, 
    -1.0569270445696612e-10, -1.0511744716853412e-10, 
    -1.0451609092104143e-10, -1.0389161367328384e-10, 
    -1.0324688154187972e-10, -1.0258485177963753e-10, 
    -1.0190878494150979e-10, -1.0122243210237201e-10, 
    -1.0053016945030482e-10, -9.9837076339225289e-11, 
    -9.9148916922875958e-11, -9.8472057569530177e-11, 
    -9.7813306222002033e-11, -9.7179703388288322e-11, 
    -9.6578279326605001e-11, -9.6015826377759533e-11, 
    -9.5498692911697211e-11, -9.50326415704013e-11, -9.46227733666207e-11, 
    -9.4273530713053983e-11, -9.3988769513364441e-11, 
    -9.3771875615790257e-11, -9.3625914250390904e-11, 
    -9.3553760758119499e-11, -9.3558190743108134e-11, 
    -9.3641893716469247e-11, -9.3807401804581046e-11, 
    -9.4056907388567137e-11, -9.4391981432879108e-11, 
    -9.4813214744070456e-11, -9.5319813886913369e-11, 
    -9.5909190455185955e-11, -9.6576591552618747e-11, 
    -9.7314827584402042e-11, -9.8114138326668845e-11, 
    -9.8962225102714311e-11, -9.9844477630928879e-11, -1.007443950835993e-10, 
    -1.0164417759999785e-10, -1.0252546822093809e-10, 
    -1.0337018105430258e-10, -1.0416136592930529e-10, -1.048840449091764e-10, 
    -1.0552595466906234e-10, -1.0607813711295191e-10, 
    -1.0653533948415012e-10, -1.0689618591933401e-10, 
    -1.0716311646401284e-10, -1.0734209613525889e-10, 
    -1.0744212013315721e-10, -1.0747455203776407e-10, 
    -1.0745235360368869e-10, -1.0738924671760789e-10, 
    -1.0729889509756622e-10, -1.0719413333571873e-10, 
    -1.0708632519082813e-10, -1.0698486087209116e-10, 
    -1.0689684424019685e-10, -1.068269600777606e-10, -1.0677752508840515e-10, 
    -1.067487003609829e-10, -1.0673882393868125e-10, -1.0674483361816563e-10, 
    -1.0676272322447928e-10, -1.0678800949363666e-10, 
    -1.0681616019008204e-10, -1.068429686877157e-10, -1.0686485939759933e-10, 
    -1.0687912249890758e-10, -1.0688406786470634e-10,
  // Sqw-F(8, 0-1999)
    0.019794563054794996, 0.019792074128530197, 0.019784629834060999, 
    0.019772296272408774, 0.019755179227821437, 0.019733418010918206, 
    0.019707177644694093, 0.019676640120572859, 0.019641995545845364, 
    0.019603434014026182, 0.019561138945140926, 0.019515282463667367, 
    0.019466023121808274, 0.019413505964081583, 0.019357864607813198, 
    0.019299224732043749, 0.019237708172214592, 0.019173436746418675, 
    0.019106535007980433, 0.019037131320811335, 0.018965356955121516, 
    0.018891343248183149, 0.018815217204171172, 0.018737096157506541, 
    0.018657082250155606, 0.018575257455429928, 0.018491679730093476, 
    0.018406380632715092, 0.018319364468842303, 0.018230608778703663, 
    0.018140065827741289, 0.018047664728654114, 0.017953313918869247, 
    0.01785690390990257, 0.017758310459148597, 0.017657398520964301, 
    0.017554027446041263, 0.017448057868429526, 0.017339360531615822, 
    0.017227826978515541, 0.017113381618347082, 0.016995994262637051, 
    0.016875691877346086, 0.016752568103219383, 0.016626789102239154, 
    0.0164985945101929, 0.016368292692155357, 0.016236250054602823, 
    0.016102874788433041, 0.015968596017144954, 0.015833839826662657, 
    0.015699003999703601, 0.015564433436478474, 0.01543039821105196, 
    0.015297076009088693, 0.015164540354563291, 0.015032755604116732, 
    0.014901579210641882, 0.014770771267797512, 0.014640010870491308, 
    0.014508918380733963, 0.014377082286904409, 0.014244089000705135, 
    0.014109553667040678, 0.013973149890086398, 0.013834636229980133, 
    0.013693877424136065, 0.013550858553224524, 0.013405690808443444, 
    0.013258608108358074, 0.013109954522720742, 0.012960163228805338, 
    0.012809728478840229, 0.012659172714144394, 0.012509011445538936, 
    0.012359718768489871, 0.012211696357732796, 0.01206524848321415, 
    0.011920565033447197, 0.011777713780771963, 0.011636642256304392, 
    0.011497188715210912, 0.011359100862001802, 0.011222060357435566, 
    0.011085710709248112, 0.010949685995549118, 0.010813637986857224, 
    0.010677259592287981, 0.010540303101088052, 0.010402592346176699, 
    0.010264028595891699, 0.010124590600461888, 0.009984329711274333, 
    0.0098433613069385788, 0.0097018538817867771, 0.0095600170902221497, 
    0.009418089830165512, 0.0092763291446414341, 0.0091350003840645327, 
    0.0089943687618888445, 0.0088546921993412388, 0.0087162152181991977, 
    0.0085791636093798616, 0.0084437396645499225, 0.0083101178779144518, 
    0.0081784411679171713, 0.0080488177962514968, 0.0079213192442589009, 
    0.0077959793266735274, 0.0076727947761007784, 0.0075517274279972551, 
    0.0074327079943603772, 0.0073156412589582536, 0.0072004123820740389, 
    0.0070868938889286394, 0.0069749528473318344, 0.0068644577234594764, 
    0.0067552844397683835, 0.0066473212400628059, 0.0065404720837416129, 
    0.0064346584319577432, 0.0063298194392613456, 0.0062259107113231847, 
    0.0061229019188569489, 0.006020773657117705, 0.0059195139984944307, 
    0.0058191151950174914, 0.0057195709449296061, 0.0056208745454994404, 
    0.0055230181221756804, 0.0054259929673700948, 0.0053297908607447611, 
    0.0052344060991121374, 0.0051398378589532067, 0.0050460924643236293, 
    0.0049531851459289978, 0.0048611409521088188, 0.0047699945982429487, 
    0.0046797891983132358, 0.0045905739865916189, 0.0045024012833049746, 
    0.004415323063652497, 0.004329387539759655, 0.0042446361544765379, 
    0.0041611013187843075, 0.0040788051141943862, 0.0039977590472548598, 
    0.0039179648069688393, 0.0038394158580683682, 0.0037620996194546496, 
    0.0036859999364631398, 0.0036110995587905707, 0.0035373823764538021, 
    0.0034648352321148212, 0.0033934492048390435, 0.0033232203334755059, 
    0.0032541498059628247, 0.0031862436774974297, 0.0031195121948495979, 
    0.0030539688006116015, 0.0029896288779041229, 0.002926508282544074, 
    0.0028646217042810687, 0.0028039809066006953, 0.0027445929163627853, 
    0.0026864582660092672, 0.0026295694241969475, 0.0025739095754580515, 
    0.0025194519162077371, 0.0024661596161780997, 0.0024139865487531691, 
    0.0023628788237001264, 0.0023127770695489172, 0.0022636193223023629, 
    0.0022153442959053091, 0.002167894750894715, 0.0021212206507878186, 
    0.0020752818061809059, 0.0020300497537316547, 0.0019855086951934518, 
    0.0019416554200094129, 0.0018984982405058129, 0.0018560550676871735, 
    0.0018143508357788343, 0.0017734145359778271, 0.0017332761397537552, 
    0.0016939636796451231, 0.0016555007153698979, 0.0016179043530842149, 
    0.0015811839154959983, 0.0015453402901576072, 0.0015103659211561852, 
    0.0014762453616019747, 0.0014429562736761991, 0.0014104707493201535, 
    0.0013787568251746459, 0.0013477800757979335, 0.0013175051847790365, 
    0.0012878974100490337, 0.0012589238748349409, 0.0012305546284116654, 
    0.0012027634318230477, 0.001175528234870818, 0.0011488313240166173, 
    0.0011226591379831859, 0.0010970017691821715, 0.0010718521935350147, 
    0.001047205296257985, 0.0010230567832235488, 0.00099940208278196632, 
    0.00097623534814597916, 0.0009535486635964119, 0.00093133153859695987, 
    0.0009095707440831284, 0.00088825050809644744, 0.00086735304816504223, 
    0.00084685938045784106, 0.00082675031553535849, 0.00080700753123407246, 
    0.00078761460706669689, 0.00076855791190040882, 0.00074982725621561849, 
    0.00073141624906476787, 0.00071332233402955538, 0.00069554651364108725, 
    0.00067809280365380912, 0.00066096748369871849, 0.00064417822672601819, 
    0.00062773319514458973, 0.00061164018691843688, 0.000595905901564469, 
    0.00058053537644124512, 0.00056553162089814733, 0.00055089545285039382, 
    0.00053662552191164866, 0.00052271848744241145, 0.00050916930995860573, 
    0.00049597161054680766, 0.00048311805464356435, 0.00047060072251261723, 
    0.00045841143739778421, 0.00044654203200979707, 0.00043498454331896704, 
    0.00042373133358936403, 0.00041277514170771375, 0.00040210907309346552, 
    0.00039172653911620487, 0.00038162115845004433, 0.00037178663360685137, 
    0.00036221661631841097, 0.00035290457557535899, 0.00034384368187280234, 
    0.00033502672031699901, 0.00032644604345324207, 0.00031809357180992448, 
    0.00030996084623367408, 0.00030203913135366805, 0.00029431956441377394, 
    0.00028679333884112977, 0.00027945190791410257, 0.00027228719130351477, 
    0.00026529176646733694, 0.00025845902800939862, 0.00025178330103677873, 
    0.00024525989889644231, 0.00023888512090143211, 0.00023265619114425009, 
    0.00022657114462770709, 0.00022062867119422404, 0.00021482793072923422, 
    0.00020916835465305527, 0.00020364944878451706, 0.00019827061140149113, 
    0.00019303097800877603, 0.00018792930129412339, 0.00018296387138077216, 
    0.0001781324781154038, 0.0001734324140549355, 0.00016886051423487927, 
    0.00016441322682603351, 0.00016008670743131268, 0.00015587692899216566, 
    0.00015177979897310973, 0.00014779127558125593, 0.0001439074751821535, 
    0.00014012476376540109, 0.00013643982630167438, 0.00013284970915569601, 
    0.00012935183240942149, 0.00012594397100717812, 0.0001226242059927052, 
    0.00011939084962371452, 0.00011624235059906245, 0.00011317718774415919, 
    0.00011019376198305607, 0.00010729029703450829, 0.00010446475884145157, 
    0.00010171480224606574, 9.9037750962596639e-05, 9.6430613725839799e-05, 
    9.3890135955468533e-05, 9.1412882787515911e-05, 8.8995346290121033e-05, 
    8.663406744795324e-05, 8.4325762301151242e-05, 8.206744155404078e-05, 
    7.9856513968848603e-05, 7.7690865744246498e-05, 7.556891056325829e-05, 
    7.3489607752371975e-05, 7.1452448697680417e-05, 6.9457414043429665e-05, 
    6.7504906061921288e-05, 6.5595661840965697e-05, 6.3730653585136168e-05, 
    6.1910982446349163e-05, 6.0137772003827466e-05, 5.8412066935633688e-05, 
    5.6734741676069751e-05, 5.5106423018695041e-05, 5.3527429744204182e-05, 
    5.1997731437573965e-05, 5.0516927699515178e-05, 4.9084247946337493e-05, 
    4.7698570935493323e-05, 4.6358462087103199e-05, 4.5062225655839293e-05, 
    4.3807967929815491e-05, 4.2593666985494854e-05, 4.141724419709542e-05, 
    4.0276632741895349e-05, 3.9169838778887178e-05, 3.8094991775612141e-05, 
    3.7050381541490865e-05, 3.603448077896374e-05, 3.5045953251102471e-05, 
    3.4083648844893191e-05, 3.3146587763380085e-05, 3.2233936718942709e-05, 
    3.134498028564483e-05, 3.0479090508465164e-05, 2.9635697516938919e-05, 
    2.8814263335026703e-05, 2.8014260421117467e-05, 2.7235155808885883e-05, 
    2.6476401131749719e-05, 2.5737428347608066e-05, 2.5017650652027141e-05, 
    2.4316467858576407e-05, 2.3633275399554268e-05, 2.2967476013763707e-05, 
    2.231849310689605e-05, 2.1685784676864134e-05, 2.1068856601135793e-05, 
    2.0467274015506651e-05, 1.9880669520283147e-05, 1.9308747074712587e-05, 
    1.8751280716916394e-05, 1.820810767738669e-05, 1.767911601255117e-05, 
    1.7164227507389921e-05, 1.666337719832376e-05, 1.6176491353162204e-05, 
    1.5703466029316705e-05, 1.5244148354886551e-05, 1.4798322422752381e-05, 
    1.4365701181593299e-05, 1.3945925021633186e-05, 1.3538566986115942e-05, 
    1.3143143806987232e-05, 1.2759131369027782e-05, 1.2385982831450908e-05, 
    1.2023147517733629e-05, 1.1670088819649582e-05, 1.132629970261638e-05, 
    1.0991314872393899e-05, 1.0664719177125807e-05, 1.0346152290309351e-05, 
    1.0035310082059635e-05, 9.731943303382687e-06, 9.4358542752934546e-06, 
    9.1468922181812235e-06, 8.8649477194680175e-06, 8.5899466728360203e-06, 
    8.321843875657858e-06, 8.0606163771891306e-06, 7.8062566403294471e-06, 
    7.5587656096640387e-06, 7.3181458451206857e-06, 7.0843949560009455e-06, 
    6.8574996243998913e-06, 6.637430520358283e-06, 6.4241383736360889e-06, 
    6.2175513848266044e-06, 6.0175740461031473e-06, 5.8240873226045319e-06, 
    5.6369500402597982e-06, 5.4560012533343122e-06, 5.2810633322437156e-06, 
    5.1119455189276166e-06, 4.9484477320547563e-06, 4.7903644533781829e-06, 
    4.6374885724482004e-06, 4.4896150981890396e-06, 4.3465446550407327e-06, 
    4.2080866710431394e-06, 4.0740621422331524e-06, 3.9443058354874096e-06, 
    3.8186677822394678e-06, 3.6970139300838514e-06, 3.5792258614941235e-06, 
    3.4651995584825049e-06, 3.3548432791775275e-06, 3.2480747052099917e-06, 
    3.144817601010749e-06, 3.0449982846861079e-06, 2.9485422333073845e-06, 
    2.8553711298374073e-06, 2.7654006050904108e-06, 2.6785388451010579e-06, 
    2.5946861333450883e-06, 2.5137352941185851e-06, 2.435572911276517e-06, 
    2.3600811283868016e-06, 2.2871397983805434e-06, 2.216628746381587e-06, 
    2.1484299343963945e-06, 2.0824293649027448e-06, 2.0185186207828003e-06, 
    1.9565960019663031e-06, 1.8965672733746443e-06, 1.8383460781228368e-06, 
    1.78185408942859e-06, 1.7270209752860906e-06, 1.673784233964148e-06, 
    1.6220889327486674e-06, 1.5718873529986406e-06, 1.5231385197520015e-06, 
    1.475807578264556e-06, 1.4298649776778273e-06, 1.3852854332414034e-06, 
    1.3420466625231024e-06, 1.3001279229934463e-06, 1.2595084140580552e-06, 
    1.2201656393416183e-06, 1.1820738504748972e-06, 1.145202706579096e-06, 
    1.1095162823923974e-06, 1.0749725408223938e-06, 1.0415233546200261e-06, 
    1.0091151186062384e-06, 9.7768994346055915e-07, 9.4718736831818468e-07, 
    9.1754647874866314e-07, 8.8870827319014196e-07, 8.6061809025030728e-07, 
    8.3322789420661186e-07, 8.0649821965639349e-07, 7.8039959829992399e-07, 
    7.5491333092695541e-07, 7.3003152170148939e-07, 7.0575635595929515e-07, 
    6.8209866987223476e-07, 6.5907592460867415e-07, 6.3670975136540576e-07, 
    6.1502327194774862e-07, 5.9403841714774962e-07, 5.7377346107588027e-07, 
    5.5424096334251044e-07, 5.3544626673794866e-07, 5.1738664015258699e-07, 
    5.000510927495254e-07, 4.8342082231400532e-07, 4.6747020620215018e-07, 
    4.5216820204979373e-07, 4.3748000186450451e-07, 4.2336877736868668e-07, 
    4.0979736607641275e-07, 3.9672977217007368e-07, 3.8413239002962087e-07, 
    3.7197489507114556e-07, 3.6023078257724562e-07, 3.4887756573939978e-07, 
    3.3789666794014697e-07, 3.2727305976083593e-07, 3.1699469993703568e-07, 
    3.0705184210343765e-07, 2.9743626844152594e-07, 2.8814050800451207e-07, 
    2.7915709349438688e-07, 2.7047790499354163e-07, 2.6209364326635392e-07, 
    2.5399346700698706e-07, 2.4616481827375849e-07, 2.3859344693758143e-07, 
    2.3126362975401603e-07, 2.2415856284163593e-07, 2.1726089058786554e-07, 
    2.1055332059607746e-07, 2.0401926602761188e-07, 1.9764345437633245e-07, 
    1.9141244665085694e-07, 1.8531502198375019e-07, 1.7934239914828962e-07, 
    1.7348828523037337e-07, 1.6774876098541654e-07, 1.621220286548827e-07, 
    1.5660806000870213e-07, 1.5120818800881246e-07, 1.4592468535389955e-07, 
    1.4076036719328329e-07, 1.357182458681528e-07, 1.3080125383635265e-07, 
    1.2601203975639376e-07, 1.2135283306053545e-07, 1.1682536598497977e-07, 
    1.1243083884756075e-07, 1.0816991466239507e-07, 1.0404273161214062e-07, 
    1.0004892602196487e-07, 9.6187662500665524e-08, 9.245767155816421e-08, 
    8.8857296827676287e-08, 8.5384554579476273e-08, 8.2037206689688903e-08, 
    7.8812845972939908e-08, 7.5708989471640273e-08, 7.272317255125698e-08, 
    6.9853034234600665e-08, 6.7096383537337367e-08, 6.4451237007374704e-08, 
    6.1915820161798492e-08, 5.948852887364293e-08, 5.7167851463158504e-08, 
    5.4952256680747976e-08, 5.284005732360417e-08, 5.0829262283864222e-08, 
    4.8917431954069525e-08, 4.7101551998487606e-08, 4.5377939448417914e-08, 
    4.3742192244587319e-08, 4.218918993535593e-08, 4.0713148836350846e-08, 
    3.9307730794488738e-08, 3.7966200218991701e-08, 3.6681620440756865e-08, 
    3.5447076966394412e-08, 3.4255912953884682e-08, 3.3101960449717216e-08, 
    3.1979750597332338e-08, 3.0884686619056578e-08, 2.981316561560693e-08, 
    2.8762638524973635e-08, 2.7731602413940113e-08, 2.6719524710081286e-08, 
    2.5726705187256559e-08, 2.4754087063327752e-08, 2.380303372347396e-08, 
    2.2875090652613518e-08, 2.1971753727713425e-08, 2.1094263815062252e-08, 
    2.0243444810528098e-08, 1.9419597051769544e-08, 1.8622452200016926e-08, 
    1.7851188976292791e-08, 1.7104503296597037e-08, 1.6380721188151634e-08, 
    1.567793977626625e-08, 1.4994180053498822e-08, 1.4327535868115051e-08, 
    1.3676305456855122e-08, 1.3039095312608142e-08, 1.2414889849946066e-08, 
    1.1803084472310849e-08, 1.1203482935268069e-08, 1.061626295081612e-08, 
    1.0041915731820739e-08, 9.4811664755707252e-09, 8.9348829452494275e-09, 
    8.4039793347079827e-09, 7.889321821566068e-09, 7.3916416744310805e-09, 
    6.911460727020678e-09, 6.4490333461020506e-09, 6.0043079121713987e-09, 
    5.5769099973996191e-09, 5.1661481331322692e-09, 4.7710419960659062e-09, 
    4.3903713161518314e-09, 4.0227426207303287e-09, 3.6666694377966796e-09, 
    3.3206607269021939e-09, 2.9833113236418754e-09, 2.6533881336208779e-09, 
    2.3299057419415702e-09, 2.0121860239803835e-09, 1.6998972350668075e-09, 
    1.3930696803600825e-09, 1.0920865255204124e-09, 7.976502230946576e-10, 
    5.1072652340158088e-10, 2.3246974619131875e-10, -3.5865825586051255e-11, 
    -2.930224225260298e-10, -5.3783658165805411e-10, -7.6933126309490195e-10, 
    -9.8679570035838739e-10, -1.1898468775347662e-09, 
    -1.3784679880984514e-09, -1.5530206732885677e-09, -1.714230137159218e-09, 
    -1.8631443050266272e-09, -2.0010706392862903e-09, 
    -2.1294960034974848e-09, -2.2499966414937982e-09, 
    -2.3641459355928322e-09, -2.4734277331188653e-09, 
    -2.5791620145540409e-09, -2.6824483029476687e-09, 
    -2.7841300010360209e-09, -2.8847807732179687e-09, 
    -2.9847116831767178e-09, -3.0839962018538413e-09, 
    -3.1825086033002045e-09, -3.2799708183675762e-09, 
    -3.3760025393666039e-09, -3.4701700353581391e-09, 
    -3.5620297993616948e-09, -3.6511644518526846e-09, 
    -3.7372092225630382e-09, -3.8198685878770005e-09, 
    -3.8989232935046538e-09, -3.9742288408439699e-09, 
    -4.0457068036733994e-09, -4.1133307894163462e-09, 
    -4.1771088807793831e-09, -4.2370646414045984e-09, 
    -4.2932185764756718e-09, -4.3455720661495018e-09, -4.39409532994337e-09, 
    -4.4387209309568329e-09, -4.4793436065872068e-09, 
    -4.5158268722825805e-09, -4.5480159940783659e-09, 
    -4.5757564643570613e-09, -4.5989163270147594e-09, -4.617410411162901e-09, 
    -4.6312240997274718e-09, -4.6404343679723699e-09, 
    -4.6452258790888133e-09, -4.6459004789738642e-09, 
    -4.6428788897439523e-09, -4.6366942431048389e-09, 
    -4.6279776191539408e-09, -4.6174366285188692e-09, 
    -4.6058284087053785e-09, -4.5939289921964511e-09, 
    -4.5825009632554321e-09, -4.5722615628236944e-09, 
    -4.5638530289007855e-09, -4.5578169080218856e-09, 
    -4.5545735398737416e-09, -4.5544077441932408e-09, 
    -4.5574612037765755e-09, -4.5637318679457389e-09, -4.573080183090485e-09, 
    -4.5852418437145684e-09, -4.599846220446202e-09, -4.6164395212951843e-09, 
    -4.6345112573337125e-09, -4.6535225028159253e-09, 
    -4.6729341012768281e-09, -4.6922330803695728e-09, 
    -4.7109554853477104e-09, -4.7287042556270944e-09, 
    -4.7451610316829842e-09, -4.7600914915155765e-09, -4.77334423313966e-09, 
    -4.7848440084124659e-09, -4.7945804136333033e-09, 
    -4.8025936612481347e-09, -4.8089590523737002e-09, 
    -4.8137718419399647e-09, -4.8171337553326091e-09, 
    -4.8191421859935251e-09, -4.8198824532799887e-09, 
    -4.8194231840949729e-09, -4.8178143613905592e-09, 
    -4.8150874919208477e-09, -4.8112571012110231e-09, 
    -4.8063230299986939e-09, -4.8002730116163117e-09, 
    -4.7930854474449402e-09, -4.7847323194617154e-09, 
    -4.7751825228177177e-09, -4.7644057524404144e-09, 
    -4.7523771471536173e-09, -4.7390825256826793e-09, 
    -4.7245239856825729e-09, -4.7087252161035541e-09, 
    -4.6917359170429656e-09, -4.673634484619318e-09, -4.6545284368370621e-09, 
    -4.6345521156573612e-09, -4.6138617245967314e-09, 
    -4.5926279437223252e-09, -4.5710268955403107e-09, 
    -4.5492303025380851e-09, -4.5273959311089338e-09, 
    -4.5056592379481221e-09, -4.4841270994907088e-09, 
    -4.4628740757597298e-09, -4.4419414968244087e-09, 
    -4.4213391998677472e-09, -4.4010496540599167e-09, 
    -4.3810338642546882e-09, -4.3612385321242862e-09, 
    -4.3416037992801034e-09, -4.3220710758209839e-09, 
    -4.3025903833965204e-09, -4.2831268519253457e-09, -4.263665920450222e-09, 
    -4.2442169809740662e-09, -4.224815089206396e-09, -4.2055205966383272e-09, 
    -4.1864165161379784e-09, -4.1676037280013631e-09, 
    -4.1491941809250293e-09, -4.1313026011497682e-09, 
    -4.1140372899834276e-09, -4.0974908404681492e-09, 
    -4.0817315690541635e-09, -4.0667965232776571e-09, 
    -4.0526866459029796e-09, -4.0393645731265366e-09, 
    -4.0267551281165737e-09, -4.01474839791604e-09, -4.0032048953423953e-09, 
    -3.9919622580739568e-09, -3.9808427358780315e-09, 
    -3.9696608801618775e-09, -3.9582308196526514e-09, 
    -3.9463728332204568e-09, -3.933918988575704e-09, -3.9207179186406899e-09, 
    -3.9066387802435865e-09, -3.8915746424651715e-09, 
    -3.8754453552007811e-09, -3.8582000160972339e-09, 
    -3.8398188857310891e-09, -3.8203146273601699e-09, 
    -3.7997325194418298e-09, -3.7781494400098598e-09, 
    -3.7556712954889367e-09, -3.7324288875180821e-09, 
    -3.7085722007769836e-09, -3.684263479505296e-09, -3.6596694653364632e-09, 
    -3.6349534734174343e-09, -3.6102678972948087e-09, 
    -3.5857478353808744e-09, -3.5615063038966143e-09, 
    -3.5376314402099183e-09, -3.5141857656337038e-09, 
    -3.4912074535335588e-09, -3.4687132504911219e-09, 
    -3.4467026490535376e-09, -3.4251627190512585e-09, 
    -3.4040731001547998e-09, -3.3834106189720861e-09, 
    -3.3631532049079406e-09, -3.3432827822328236e-09, 
    -3.3237870844199755e-09, -3.3046603444051713e-09, 
    -3.2859030150010785e-09, -3.2675206335226756e-09, 
    -3.2495221062242057e-09, -3.2319175641205564e-09, 
    -3.2147161199518237e-09, -3.1979236540642043e-09, 
    -3.1815409415202742e-09, -3.1655622460672499e-09, 
    -3.1499746135522044e-09, -3.134757920672683e-09, -3.1198857686709065e-09, 
    -3.1053271420291147e-09, -3.0910487073677101e-09, 
    -3.0770174716702988e-09, -3.06320354876317e-09, -3.0495825965328548e-09, 
    -3.0361376593976133e-09, -3.0228600907839938e-09, 
    -3.0097494432413811e-09, -2.9968122597902103e-09, -2.984059957040674e-09, 
    -2.9715060027927005e-09, -2.9591628300663923e-09, 
    -2.9470387902192566e-09, -2.9351355868062683e-09, -2.923446407218947e-09, 
    -2.9119549463736257e-09, -2.900635296595257e-09, -2.8894526165382664e-09, 
    -2.8783643347290193e-09, -2.8673216754443855e-09, 
    -2.8562712261073918e-09, -2.8451564285959661e-09, 
    -2.8339188520464317e-09, -2.8224993389350964e-09, 
    -2.8108390552251555e-09, -2.7988806501354413e-09, 
    -2.7865696236213109e-09, -2.7738560196970457e-09, 
    -2.7606964210580918e-09, -2.7470561882678751e-09, 
    -2.7329117024670132e-09, -2.7182524210637822e-09, 
    -2.7030824198341604e-09, -2.6874212410142156e-09, 
    -2.6713038338796474e-09, -2.6547795910634203e-09, 
    -2.6379104927082137e-09, -2.6207685698395248e-09, 
    -2.6034328920446348e-09, -2.5859864138593919e-09, 
    -2.5685128916596859e-09, -2.5510941574363299e-09, 
    -2.5338078527714539e-09, -2.5167257373352607e-09, 
    -2.4999125216225962e-09, -2.4834251862475798e-09, 
    -2.4673126404332115e-09, -2.4516156430828557e-09, 
    -2.4363668341597752e-09, -2.4215908564152042e-09, 
    -2.4073044743384217e-09, -2.3935167527459783e-09, 
    -2.3802292606035294e-09, -2.3674363941006992e-09, 
    -2.3551257954837326e-09, -2.3432789625269112e-09, 
    -2.3318719745653281e-09, -2.3208763888750056e-09, 
    -2.3102602227139357e-09, -2.2999890319224224e-09, 
    -2.2900269853976099e-09, -2.2803379400960273e-09, 
    -2.2708864253996675e-09, -2.2616385526696733e-09, 
    -2.2525627452700605e-09, -2.2436303055640971e-09, 
    -2.2348157549260812e-09, -2.2260969487612836e-09, 
    -2.2174549301877235e-09, -2.2088735789377904e-09, 
    -2.2003390612139205e-09, -2.1918391900838799e-09, 
    -2.1833627687036445e-09, -2.1748990655270657e-09, 
    -2.1664374920901473e-09, -2.1579676142496491e-09, 
    -2.1494795008798246e-09, -2.1409644494177672e-09, 
    -2.1324159512345728e-09, -2.1238308181036492e-09, 
    -2.1152102313802011e-09, -2.1065605654598882e-09, 
    -2.0978937219783705e-09, -2.0892269045082957e-09, -2.080581669319931e-09, 
    -2.0719823450833882e-09, -2.0634538616183869e-09, 
    -2.0550192545065085e-09, -2.0466970395034402e-09, 
    -2.0384988379172268e-09, -2.0304274559070779e-09, 
    -2.0224757311721439e-09, -2.0146262622794976e-09, 
    -2.0068521178211987e-09, -1.9991184284095081e-09, 
    -1.9913847726017363e-09, -1.98360805085681e-09, -1.9757456386801034e-09, 
    -1.9677584497993977e-09, -1.9596136952429695e-09, 
    -1.9512870481515724e-09, -1.9427641358569156e-09, 
    -1.9340412013999598e-09, -1.9251250180682261e-09, 
    -1.9160320791192621e-09, -1.9067872549302563e-09, 
    -1.8974220146688509e-09, -1.8879724626050447e-09, 
    -1.8784772875885138e-09, -1.8689758295002255e-09, 
    -1.8595063121136343e-09, -1.8501044057980474e-09, 
    -1.8408020595876732e-09, -1.8316267115495697e-09, -1.822600799157708e-09, 
    -1.8137416012082351e-09, -1.8050613141860271e-09, 
    -1.7965673729062813e-09, -1.7882629018492612e-09, 
    -1.7801473038072591e-09, -1.7722168622397551e-09, 
    -1.7644653660497267e-09, -1.7568846407040178e-09, 
    -1.7494650403253694e-09, -1.7421957851175858e-09, 
    -1.7350652427854418e-09, -1.728061086534514e-09, -1.7211704483687201e-09, 
    -1.7143800262865769e-09, -1.707676270302587e-09, -1.701045588453083e-09, 
    -1.6944746655845723e-09, -1.6879507960937239e-09, 
    -1.6814622804687619e-09, -1.6749987267671125e-09, 
    -1.6685512921071363e-09, -1.6621127091296038e-09, 
    -1.6556771274313571e-09, -1.6492396774257275e-09, 
    -1.6427958778345286e-09, -1.6363408258046387e-09, 
    -1.6298683825621989e-09, -1.6233703689801574e-09, 
    -1.6168359841010687e-09, -1.6102514746146146e-09, -1.603600229918887e-09, 
    -1.5968632547664763e-09, -1.5900201060962778e-09, 
    -1.5830501530053288e-09, -1.5759341470194086e-09, 
    -1.5686558840600557e-09, -1.561203877686043e-09, -1.5535728110356216e-09, 
    -1.545764698485353e-09, -1.5377895471099852e-09, -1.5296655245161068e-09, 
    -1.5214184995923381e-09, -1.5130810656071357e-09, 
    -1.5046910065486688e-09, -1.4962893998788836e-09, 
    -1.4879184103939451e-09, -1.4796190261772871e-09, 
    -1.4714288303166709e-09, -1.4633800583464674e-09, 
    -1.4554980290288491e-09, -1.4478001525178939e-09, 
    -1.4402954992703834e-09, -1.432985069567028e-09, -1.4258626188040961e-09, 
    -1.4189160490696595e-09, -1.4121291577335085e-09, 
    -1.4054836346053595e-09, -1.398961051427203e-09, -1.3925447343649184e-09, 
    -1.3862212511762986e-09, -1.3799814901331126e-09, 
    -1.3738211348865901e-09, -1.367740618175716e-09, -1.3617444898622583e-09, 
    -1.3558403813037057e-09, -1.3500376114398143e-09, 
    -1.3443456689475822e-09, -1.3387726687017769e-09, 
    -1.3333240161335264e-09, -1.3280013310634309e-09, 
    -1.3228018050741238e-09, -1.3177179590957188e-09, 
    -1.3127378930362811e-09, -1.3078458855670885e-09, 
    -1.3030233380610023e-09, -1.2982499038759741e-09, 
    -1.2935047445781992e-09, -1.2887677132666078e-09, 
    -1.2840204837271778e-09, -1.2792474250672712e-09, -1.274436294586426e-09, 
    -1.2695786265026495e-09, -1.2646699177404633e-09, 
    -1.2597095461020758e-09, -1.2547005362716775e-09, 
    -1.2496491364825363e-09, -1.2445643138036522e-09, 
    -1.2394571228233029e-09, -1.234340064408701e-09, -1.2292263542909878e-09, 
    -1.2241292230013426e-09, -1.2190611874263808e-09, 
    -1.2140334020061752e-09, -1.2090550419861225e-09, -1.204132842333544e-09, 
    -1.1992707403796558e-09, -1.1944697397328715e-09, 
    -1.1897279255930957e-09, -1.1850407177130768e-09, -1.1804012633227109e-09, 
    -1.1758010145735932e-09, -1.1712303629140453e-09, 
    -1.1666793559486962e-09, -1.162138349265094e-09, -1.1575986335374912e-09, 
    -1.1530528912244936e-09, -1.1484955783121041e-09, 
    -1.1439230919951913e-09, -1.139333858292246e-09, -1.1347282625108184e-09, 
    -1.1301085203806674e-09, -1.1254784739402903e-09, 
    -1.1208433949410377e-09, -1.1162097400272352e-09, 
    -1.1115849540915295e-09, -1.1069772245304683e-09, -1.102395273814226e-09, 
    -1.0978480696996509e-09, -1.0933445393284206e-09, 
    -1.0888931797411308e-09, -1.0845016557671756e-09, -1.080176318686225e-09, 
    -1.0759217491805087e-09, -1.0717403032304322e-09, 
    -1.0676317774395594e-09, -1.0635931756635463e-09, 
    -1.0596187165520161e-09, -1.0557000104853052e-09, -1.051826529987116e-09, 
    -1.0479862501629226e-09, -1.0441665206868839e-09, 
    -1.0403550004874033e-09, -1.036540661539324e-09, -1.0327146708685028e-09, 
    -1.0288711381407715e-09, -1.0250075613455909e-09, 
    -1.0211249985920563e-09, -1.0172278527544146e-09, 
    -1.0133233815978631e-09, -1.0094208907961897e-09, 
    -1.0055308058367109e-09, -1.0016636278365239e-09, 
    -9.9782899947456386e-10, -9.9403490428475653e-10, 
    -9.9028716373986435e-10, -9.8658922487120815e-10, 
    -9.8294230090607858e-10, -9.7934577586262265e-10, 
    -9.7579785442518138e-10, -9.7229627453616374e-10, 
    -9.6883903942902204e-10, -9.6542497104328338e-10, 
    -9.6205405886455739e-10, -9.587274742304845e-10, -9.5544730115812049e-10, 
    -9.5221594744804503e-10, -9.4903539560610659e-10, 
    -9.4590632001360758e-10, -9.4282727747575168e-10, 
    -9.3979403195395517e-10, -9.3679918507110889e-10, 
    -9.3383211288321781e-10, -9.3087931623850697e-10, -9.279250772474945e-10, 
    -9.2495244021925953e-10, -9.2194433393071003e-10, 
    -9.1888480382678248e-10, -9.1576013627689331e-10, 
    -9.1255986224716403e-10, -9.0927745905807821e-10, 
    -9.0591078499544297e-10, -9.0246215945722002e-10, 
    -8.9893816442361382e-10, -8.9534916854153287e-10, 
    -8.9170869331472796e-10, -8.8803263843137021e-10, 
    -8.8433851146678318e-10, -8.8064465643308785e-10, 
    -8.7696961213724698e-10, -8.733315518517321e-10, -8.6974789584398184e-10, 
    -8.6623501047250397e-10, -8.628080489702643e-10, -8.5948080999477729e-10, 
    -8.5626566370752513e-10, -8.5317340475948093e-10, 
    -8.5021309614158714e-10, -8.4739177020261017e-10, -8.447141073786703e-10, 
    -8.4218197705543111e-10, -8.3979399609534136e-10, -8.375450642947118e-10, 
    -8.3542602601654051e-10, -8.3342346267575858e-10, 
    -8.3151973584890661e-10, -8.296932846999571e-10, -8.2791923868323724e-10, 
    -8.2617029634899357e-10, -8.2441787590863668e-10, 
    -8.2263340557857443e-10, -8.2078971932508742e-10, 
    -8.1886239727633965e-10, -8.1683098947847082e-10, 
    -8.1467999320894098e-10, -8.1239954225783945e-10, 
    -8.0998573541654017e-10, -8.0744063120671772e-10, 
    -8.0477187534592505e-10, -8.0199205331888092e-10, 
    -7.9911778481785926e-10, -7.9616866906789713e-10, 
    -7.9316611028371458e-10, -7.9013215193501203e-10, 
    -7.8708832926423714e-10, -7.8405465378995476e-10, 
    -7.8104873134998589e-10, -7.7808510457146974e-10, -7.75174790945784e-10, 
    -7.7232507375059925e-10, -7.6953951091449149e-10, -7.668181621185628e-10, 
    -7.6415798534727172e-10, -7.6155337443906035e-10, 
    -7.5899675889046594e-10, -7.5647925195294078e-10, 
    -7.5399124866178264e-10, -7.515229821462162e-10, -7.4906496917004927e-10, 
    -7.466083688447168e-10, -7.441452270243621e-10, -7.4166864662854755e-10, 
    -7.3917288521668128e-10, -7.3665342494792328e-10, 
    -7.3410701629840659e-10, -7.3153172748489304e-10, 
    -7.2892698917969617e-10, -7.2629366987610912e-10, 
    -7.2363410048894013e-10, -7.2095213331774033e-10, 
    -7.1825311056465714e-10, -7.1554381530538446e-10, 
    -7.1283232690341727e-10, -7.1012782048025715e-10, 
    -7.0744026333260399e-10, -7.0478007411836892e-10, 
    -7.0215768846777378e-10, -6.9958311157161791e-10, 
    -6.9706543642630266e-10, -6.9461238483009392e-10, -6.92229870868373e-10, 
    -6.8992163088316187e-10, -6.8768892020322647e-10, -6.855303200005389e-10, 
    -6.83441626974252e-10, -6.8141587174034584e-10, -6.7944343228663178e-10, 
    -6.7751226621463535e-10, -6.7560823793329361e-10, -6.737155578061613e-10, 
    -6.7181730019528569e-10, -6.698960161535755e-10, -6.6793441405359951e-10, 
    -6.6591610248782615e-10, -6.6382635589726894e-10, 
    -6.6165289401263406e-10, -6.5938659849545751e-10, 
    -6.5702217198653909e-10, -6.5455862247679539e-10, -6.519995830217703e-10, 
    -6.4935337239135998e-10, -6.4663280350486851e-10, 
    -6.4385468223752621e-10, -6.4103905349826334e-10, 
    -6.3820816319043385e-10, -6.3538524275528641e-10, 
    -6.3259315041936977e-10, -6.2985298355987247e-10, 
    -6.2718274869979103e-10, -6.2459620720043572e-10, 
    -6.2210196437976583e-10, -6.1970293056483942e-10, 
    -6.1739615200197961e-10, -6.1517308729148928e-10, 
    -6.1302027858852446e-10, -6.1092040797114254e-10, 
    -6.0885361727157599e-10, -6.0679902076731403e-10, 
    -6.0473625419255301e-10, -6.0264694880832519e-10, 
    -6.0051600037286642e-10, -5.9833253264961123e-10, 
    -5.9609048058658688e-10, -5.9378878379934686e-10, -5.914311627601923e-10, 
    -5.8902556961823619e-10, -5.865833419747216e-10, -5.8411819926547477e-10, 
    -5.8164513660645888e-10, -5.7917936440826231e-10, 
    -5.7673532420917178e-10, -5.7432587860238123e-10, -5.71961689812886e-10, 
    -5.6965082556433647e-10, -5.6739856501047267e-10, -5.652074094508503e-10, 
    -5.6307725633427454e-10, -5.6100573334155574e-10, 
    -5.5898862329650417e-10, -5.5702039596439675e-10, -5.55094760551569e-10, 
    -5.5320526182287836e-10, -5.5134582649148551e-10, -5.495112656164138e-10, 
    -5.4769766302244816e-10, -5.4590264517924988e-10, 
    -5.4412548027924872e-10, -5.4236701832053593e-10, -5.406294540834214e-10, 
    -5.3891595747668599e-10, -5.3723017272932343e-10, 
    -5.3557568027663113e-10, -5.3395542626947468e-10, 
    -5.3237123424395042e-10, -5.3082339688680504e-10, 
    -5.2931044346573756e-10, -5.2782906516280041e-10, 
    -5.2637425981819642e-10, -5.2493962236141568e-10, 
    -5.2351782128726248e-10, -5.2210115105355352e-10, 
    -5.2068215930652611e-10, -5.1925423340170444e-10, 
    -5.1781213778385308e-10, -5.1635239292709779e-10, 
    -5.1487350201352995e-10, -5.1337595891078236e-10, 
    -5.1186208631200535e-10, -5.1033565937203448e-10, 
    -5.0880142399954457e-10, -5.0726450349115863e-10, 
    -5.0572980078664856e-10, -5.0420143294398164e-10, 
    -5.0268227783756706e-10, -5.0117365341427345e-10, 
    -4.9967518128569356e-10, -4.9818480913907182e-10, 
    -4.9669902034902165e-10, -4.9521313236964123e-10, 
    -4.9372172100469227e-10, -4.9221904180436789e-10, 
    -4.9069945189863883e-10, -4.8915776479024795e-10, 
    -4.8758953132497268e-10, -4.8599118900544138e-10, 
    -4.8436014460717885e-10, -4.8269472369992403e-10, -4.809940902780113e-10, 
    -4.7925809219519262e-10, -4.7748712349103488e-10, 
    -4.7568198386527302e-10, -4.7384380352808874e-10, 
    -4.7197399759148612e-10, -4.7007430876179642e-10, 
    -4.6814688310359711e-10, -4.6619441078452655e-10, 
    -4.6422026695619175e-10, -4.6222868051353304e-10, 
    -4.6022484455877117e-10, -4.5821501274448725e-10, 
    -4.5620649912135189e-10, -4.5420762138105684e-10, 
    -4.5222754212437032e-10, -4.5027605867666611e-10, 
    -4.4836328927656393e-10, -4.4649935419213988e-10, 
    -4.4469398267306598e-10, -4.4295615754756096e-10, -4.4129374085866e-10, 
    -4.3971317837224967e-10, -4.3821923332650135e-10, 
    -4.3681482788050671e-10, -4.3550094989000611e-10, 
    -4.3427669084424681e-10, -4.3313934822863559e-10, 
    -4.3208466587874914e-10, -4.3110712553061738e-10, 
    -4.3020033289006323e-10, -4.2935742153369603e-10, 
    -4.2857150366557418e-10, -4.278360598457436e-10, -4.2714531222150651e-10, 
    -4.2649447649723079e-10, -4.2587992511249538e-10, 
    -4.2529918589146491e-10, -4.2475084327476837e-10, 
    -4.2423426435948439e-10, -4.2374925305527341e-10, 
    -4.2329560750540744e-10, -4.2287267449546696e-10, 
    -4.2247891363523962e-10, -4.2211156942225334e-10, 
    -4.2176644739347364e-10, -4.2143788904004336e-10, 
    -4.2111889182270629e-10, -4.2080145127221426e-10, 
    -4.2047700475517344e-10, -4.2013701310202405e-10, 
    -4.1977354271592666e-10, -4.1937983330032509e-10, -4.189507160251554e-10, 
    -4.184828997410636e-10, -4.179749924749733e-10, -4.1742734645043684e-10, 
    -4.1684166285877366e-10, -4.1622046108029893e-10, 
    -4.1556644584468218e-10, -4.1488190626253303e-10, 
    -4.1416816777157904e-10, -4.1342523262048676e-10, 
    -4.1265161182038015e-10, -4.1184441250445422e-10, 
    -4.1099961540964467e-10, -4.1011256366953406e-10, 
    -4.0917852876717771e-10, -4.0819332925762842e-10, 
    -4.0715387367114772e-10, -4.0605861533369016e-10, 
    -4.0490779695544773e-10, -4.037035324197919e-10, -4.024496627490239e-10, 
    -4.0115148788448044e-10, -3.9981534020611453e-10, 
    -3.9844812155549981e-10, -3.9705681413834002e-10, 
    -3.9564806092060442e-10, -3.9422780064152914e-10, 
    -3.9280104855393438e-10, -3.9137176536114289e-10, 
    -3.8994288066605685e-10, -3.8851639530995144e-10, 
    -3.8709359906805403e-10, -3.8567532657790783e-10, 
    -3.8426228209130485e-10, -3.8285534143359229e-10, 
    -3.8145586377561918e-10, -3.8006592313488588e-10, 
    -3.7868848925491449e-10, -3.7732747521390679e-10, 
    -3.7598769602882313e-10, -3.7467465954642051e-10, 
    -3.7339425973795677e-10, -3.7215232595266755e-10, 
    -3.7095413700549558e-10, -3.6980387387140909e-10, 
    -3.6870412667744685e-10, -3.6765547474191712e-10, 
    -3.6665625955617799e-10, -3.6570251884502316e-10, 
    -3.6478817307633289e-10, -3.6390541589940587e-10, 
    -3.6304532802420888e-10, -3.6219859822919916e-10, 
    -3.6135634076978954e-10, -3.6051086520195884e-10, 
    -3.5965636039469326e-10, -3.5878937051820585e-10, 
    -3.5790906649886764e-10, -3.5701721212333898e-10, 
    -3.5611790607333362e-10, -3.552170539991811e-10, -3.5432169778879464e-10, 
    -3.5343919751307955e-10, -3.5257641573239501e-10, -3.517389049452622e-10, 
    -3.5093023916388747e-10, -3.5015147216463898e-10, 
    -3.4940082462778088e-10, -3.4867356210792838e-10, 
    -3.4796213781966551e-10, -3.4725652569406252e-10, 
    -3.4654478190118062e-10, -3.458137510719682e-10, -3.4504993906139904e-10, 
    -3.4424042600630226e-10, -3.4337381504252164e-10, 
    -3.4244111748638184e-10, -3.4143652290080135e-10, -3.40357972790168e-10, 
    -3.3920750971270144e-10, -3.3799133332148421e-10, 
    -3.3671958851098844e-10, -3.3540586520179414e-10, 
    -3.3406648647702024e-10, -3.3271960751264808e-10, 
    -3.3138424352623405e-10, -3.3007926747369318e-10, 
    -3.2882250911556471e-10, -3.276299658968534e-10, -3.265152271714507e-10, 
    -3.2548907969248937e-10, -3.2455935601983365e-10, -3.237309347613477e-10, 
    -3.2300590764096794e-10, -3.2238381476652182e-10, 
    -3.2186196164157519e-10, -3.2143570263464149e-10, -3.210987227622085e-10, 
    -3.2084325874026917e-10, -3.2066028672871032e-10, 
    -3.2053964980891089e-10, -3.2047020458963292e-10, 
    -3.2043993242523419e-10, -3.2043608911531305e-10, -3.204453789507471e-10, 
    -3.2045418944085798e-10, -3.2044884395809632e-10, 
    -3.2041591579677564e-10, -3.2034254576672231e-10, -3.202167953186203e-10, 
    -3.2002797476781496e-10, -3.1976697466028162e-10, 
    -3.1942654410118567e-10, -3.1900154781772349e-10, 
    -3.1848914324131111e-10, -3.1788890500946058e-10, 
    -3.1720284964772764e-10, -3.1643540227513006e-10, 
    -3.1559323947416522e-10, -3.1468506428341138e-10, 
    -3.1372127594632566e-10, -3.1271359309642672e-10, 
    -3.1167459332013004e-10, -3.1061726528093259e-10, 
    -3.0955452698169761e-10, -3.0849879276961018e-10, 
    -3.0746156683332184e-10, -3.0645313268141984e-10, 
    -3.0548228396512918e-10, -3.0455614745855808e-10, 
    -3.0368005515834167e-10, -3.0285750381154751e-10, 
    -3.0209013517155345e-10, -3.0137777513849486e-10, 
    -3.0071849406269827e-10, -3.0010873317157956e-10, 
    -2.9954343638024177e-10, -2.9901625457792673e-10, 
    -2.9851977411198144e-10, -2.980458153241456e-10, -2.9758573932891178e-10, 
    -2.9713080864021193e-10, -2.9667252479423753e-10, 
    -2.9620296485221772e-10, -2.9571505294994394e-10, 
    -2.9520278925752169e-10, -2.94661368522997e-10, -2.9408723026780942e-10, 
    -2.9347800482821403e-10, -2.9283239353983424e-10, 
    -2.9214998965700809e-10, -2.9143108187417703e-10, 
    -2.9067643629938836e-10, -2.8988714320353919e-10, 
    -2.8906447474709357e-10, -2.8820982958075172e-10, 
    -2.8732471491906458e-10, -2.8641081062776607e-10, 
    -2.8547003922530795e-10, -2.8450466726864581e-10, 
    -2.8351737843644551e-10, -2.8251133189318618e-10, 
    -2.8149014569569902e-10, -2.8045784369950152e-10, 
    -2.7941873148052868e-10, -2.7837723764861951e-10, 
    -2.7733772582234253e-10, -2.7630430882469188e-10, -2.752806708988115e-10, 
    -2.742699520758142e-10, -2.7327465555879554e-10, -2.7229663282171393e-10, 
    -2.7133710888055876e-10, -2.7039676793267066e-10, 
    -2.6947585407883417e-10, -2.6857431794979981e-10, 
    -2.6769195172051162e-10, -2.6682853786209857e-10, -2.659839618077944e-10, 
    -2.6515833874860445e-10, -2.6435207296380715e-10, -2.635658998126444e-10, 
    -2.6280085707744182e-10, -2.6205822479745353e-10, 
    -2.6133937626869825e-10, -2.6064558924517683e-10, -2.599777938369407e-10, 
    -2.5933630810759921e-10, -2.5872054139623211e-10, 
    -2.5812877189287469e-10, -2.5755795772025962e-10, 
    -2.5700366036859779e-10, -2.5646008986670765e-10, 
    -2.5592029448292568e-10, -2.5537646277275915e-10, 
    -2.5482035850668645e-10, -2.5424381143716496e-10, 
    -2.5363926663319388e-10, -2.5300029218141947e-10, 
    -2.5232206436504831e-10, -2.5160173056821574e-10, 
    -2.5083866038780301e-10, -2.5003455570550197e-10, 
    -2.4919341887601776e-10, -2.4832137283521286e-10, 
    -2.4742637777342588e-10, -2.4651781287981132e-10, 
    -2.4560600151163241e-10, -2.447016526003258e-10, -2.4381528451113753e-10, 
    -2.4295661860031455e-10, -2.421340224122714e-10, -2.4135398641542728e-10, 
    -2.4062069789905979e-10, -2.3993573557352927e-10, 
    -2.3929792499833876e-10, -2.3870335603799221e-10, 
    -2.3814559127660717e-10, -2.3761603774694772e-10, 
    -2.3710448191518258e-10, -2.3659971208691608e-10, 
    -2.3609021980059018e-10, -2.3556486983288133e-10, 
    -2.3501353021455081e-10, -2.3442757023294742e-10, 
    -2.3380020998594916e-10, -2.3312668849385971e-10, 
    -2.3240428279615229e-10, -2.3163214604905193e-10, 
    -2.3081105144228282e-10, -2.2994304645900058e-10, 
    -2.2903109742334705e-10, -2.2807873729331133e-10, 
    -2.2708977628495047e-10, -2.2606807664324935e-10, 
    -2.2501741688708671e-10, -2.2394143341961978e-10, 
    -2.2284363189358524e-10, -2.2172744721968785e-10, -2.205963492559654e-10, 
    -2.1945394972919954e-10, -2.1830414536857467e-10, 
    -2.1715123767652849e-10, -2.1600006813776193e-10, 
    -2.1485613270659579e-10, -2.1372570741567318e-10, 
    -2.1261593928100675e-10, -2.1153492549669576e-10, 
    -2.1049174046331641e-10, -2.0949640624842698e-10, 
    -2.0855977619859425e-10, -2.0769332941396211e-10, 
    -2.0690883637296042e-10, -2.0621793902792313e-10, 
    -2.0563160613879809e-10, -2.0515953121179496e-10, -2.048094835727676e-10, 
    -2.0458669195174352e-10, -2.0449328182200974e-10, 
    -2.0452785440174509e-10, -2.0468524869422683e-10, 
    -2.0495650921625231e-10, -2.0532909787363608e-10, -2.057873507521604e-10, 
    -2.0631312758221949e-10, -2.0688663841471605e-10, 
    -2.0748735032587637e-10, -2.0809494760309469e-10, -2.086902221453167e-10, 
    -2.0925585479731438e-10, -2.0977702539675372e-10, 
    -2.1024182622474911e-10, -2.1064144839935413e-10, 
    -2.1097016972407398e-10, -2.1122515347620451e-10, 
    -2.1140612534965196e-10, -2.1151494688840785e-10, 
    -2.1155516586460856e-10, -2.1153155660449197e-10, 
    -2.1144972089714611e-10, -2.113157327267807e-10, -2.1113587030934217e-10, 
    -2.109164015169028e-10, -2.1066345406237256e-10, -2.1038291218613182e-10, 
    -2.1008035927740021e-10, -2.0976104276808983e-10, 
    -2.0942984586527921e-10, -2.0909127193344966e-10, 
    -2.0874943962129786e-10, -2.0840807265662676e-10, 
    -2.0807050469733046e-10, -2.0773967866650546e-10, 
    -2.0741816181729703e-10, -2.071081445532783e-10, -2.0681145912686622e-10, 
    -2.0652958232285931e-10, -2.0626365198475409e-10, 
    -2.0601448458562697e-10, -2.0578261001373738e-10, 
    -2.0556831489738862e-10, -2.0537171027422335e-10, 
    -2.0519280569912155e-10, -2.050315920373089e-10, -2.0488810762899577e-10, 
    -2.0476249649772124e-10, -2.0465501507628202e-10, 
    -2.0456599391319383e-10, -2.044957471452107e-10, -2.0444444721499725e-10, 
    -2.0441195458763394e-10, -2.0439765011316801e-10, 
    -2.0440028635107451e-10, -2.0441788882291089e-10, 
    -2.0444771753654351e-10, -2.0448633342365196e-10, -2.045297252753035e-10, 
    -2.0457351588771751e-10, -2.0461321805390606e-10, 
    -2.0464450008837741e-10, -2.0466343693346274e-10, 
    -2.0466672068459352e-10, -2.0465180478933769e-10, 
    -2.0461695849185276e-10, -2.045612515391146e-10, -2.0448448067481462e-10, 
    -2.0438702786413915e-10, -2.0426969863619459e-10, 
    -2.0413354164346943e-10, -2.0397967753975899e-10, -2.038091420793715e-10, 
    -2.0362275327880125e-10, -2.0342100093336653e-10, 
    -2.0320397702172393e-10, -2.0297132652599141e-10, -2.027222373242946e-10, 
    -2.0245546213423163e-10, -2.0216938687200365e-10, -2.01862134870881e-10, 
    -2.0153170722507694e-10, -2.0117615235445015e-10, 
    -2.0079376154345746e-10, -2.003832541113059e-10, -1.9994395015427916e-10, 
    -1.9947589862752684e-10, -1.9897995831009526e-10, -1.984578133361114e-10, 
    -1.9791191553051972e-10, -1.9734538240513937e-10, 
    -1.9676184981187532e-10, -1.9616529753550445e-10, 
    -1.9555990437838086e-10, -1.9494990882702465e-10, 
    -1.9433953264068712e-10, -1.9373296163194426e-10, 
    -1.9313437261070207e-10, -1.9254800694488779e-10, 
    -1.9197826698584984e-10, -1.9142978924591532e-10, 
    -1.9090747763861934e-10, -1.9041645667726749e-10, 
    -1.8996193267622252e-10, -1.8954893818335841e-10, 
    -1.8918199357689077e-10, -1.888646922624807e-10, -1.8859925090680121e-10, 
    -1.8838609235669215e-10, -1.8822352147117868e-10, 
    -1.8810753035369027e-10, -1.8803180927242878e-10, -1.879879665236587e-10, 
    -1.8796597579711002e-10, -1.8795482166259606e-10, 
    -1.8794329098781355e-10, -1.8792083507465885e-10, 
    -1.8787841882098224e-10, -1.8780924940813249e-10, 
    -1.8770931157028736e-10, -1.8757762184505196e-10, 
    -1.8741618771317053e-10, -1.8722964240989857e-10, 
    -1.8702459919541174e-10, -1.8680879806371849e-10, 
    -1.8659013831639704e-10, -1.8637570204954168e-10, 
    -1.8617088868532256e-10, -1.8597875679018906e-10, 
    -1.8579964347715407e-10, -1.856311018465997e-10, -1.8546814961498825e-10, 
    -1.8530379150581812e-10, -1.8512973513314712e-10, 
    -1.8493720743388612e-10, -1.8471778030129572e-10, 
    -1.8446409348911562e-10, -1.8417041462003943e-10, 
    -1.8383298063620771e-10, -1.8345012310224288e-10, 
    -1.8302217411105298e-10, -1.825512101474751e-10, -1.8204068749149685e-10, 
    -1.8149504182634588e-10, -1.8091929849457328e-10, 
    -1.8031874506636372e-10, -1.7969869342020501e-10, 
    -1.7906433520553629e-10, -1.7842067625609343e-10, 
    -1.7777253066317654e-10, -1.7712453658481296e-10, 
    -1.7648117449203098e-10, -1.7584675314966835e-10, 
    -1.7522537192752909e-10, -1.7462083620182323e-10, 
    -1.7403656316481032e-10, -1.7347548042098988e-10, 
    -1.7293994487534775e-10, -1.724317015635456e-10, -1.7195190342064396e-10, 
    -1.7150118278464737e-10, -1.7107978537556873e-10, 
    -1.7068774010356032e-10, -1.7032505721590001e-10, 
    -1.6999192690949003e-10, -1.6968888671709507e-10, 
    -1.6941694603304543e-10, -1.691776609812933e-10, -1.6897311346254065e-10, 
    -1.6880583666032105e-10, -1.686786481396406e-10, -1.6859441609306793e-10, 
    -1.6855576842641605e-10, -1.6856475414013642e-10, 
    -1.6862247143394776e-10, -1.6872870141468215e-10, 
    -1.6888154237075115e-10, -1.6907711460567902e-10, 
    -1.6930931865872873e-10, -1.6956973192822121e-10, 
    -1.6984762590944127e-10, -1.701301557429917e-10, -1.7040272835710173e-10, 
    -1.7064954370420615e-10, -1.7085429232978048e-10, 
    -1.7100098556104489e-10, -1.7107484737301839e-10, 
    -1.7106322569844794e-10, -1.7095642840071364e-10, 
    -1.7074844580314795e-10, -1.7043746272138936e-10, 
    -1.7002612810308226e-10, -1.6952153955760311e-10, 
    -1.6893495959000206e-10, -1.6828123099042661e-10, 
    -1.6757797775376145e-10, -1.6684460834767992e-10, 
    -1.6610121438792032e-10, -1.6536743435154181e-10, -1.646613679938315e-10, 
    -1.6399860623331646e-10, -1.6339147888734139e-10, 
    -1.6284851816181356e-10, -1.6237424681714827e-10, 
    -1.6196922377029712e-10, -1.6163040641791073e-10, 
    -1.6135175272099892e-10, -1.61125020972039e-10, -1.6094069231352511e-10, 
    -1.6078895170416783e-10, -1.6066060585454966e-10, 
    -1.6054789413688827e-10, -1.604450947103901e-10, -1.6034891217939672e-10, 
    -1.6025858675239268e-10, -1.6017576639398427e-10, 
    -1.6010414534227762e-10, -1.6004892082202286e-10, 
    -1.6001613805505281e-10, -1.6001200131026202e-10, 
    -1.6004218354845135e-10, -1.6011122638637136e-10, 
    -1.6022204818949052e-10, -1.6037560416901553e-10, 
    -1.6057069023360024e-10, -1.6080390368773475e-10, 
    -1.6106972590585351e-10, -1.6136072849041324e-10, 
    -1.6166785583654076e-10, -1.6198079956811689e-10, 
    -1.6228840203580649e-10, -1.6257912427453815e-10, 
    -1.6284153540557574e-10, -1.6306482547216528e-10, 
    -1.6323932301330732e-10, -1.6335702767808538e-10, 
    -1.6341208286654041e-10, -1.6340120749836769e-10, 
    -1.6332401669704194e-10, -1.6318322336453046e-10, 
    -1.6298466750270051e-10, -1.6273715391615785e-10, 
    -1.6245208842146761e-10, -1.6214291371720495e-10, 
    -1.6182435730995891e-10, -1.6151155407883618e-10, 
    -1.6121906134348955e-10, -1.609598844978556e-10, -1.6074454306517733e-10, 
    -1.6058029138411775e-10, -1.6047054088754121e-10, 
    -1.6041455675167418e-10, -1.6040745093278731e-10, 
    -1.6044049697628079e-10, -1.6050173007925778e-10, 
    -1.6057680823489771e-10, -1.6065003495563594e-10, 
    -1.6070550064571938e-10, -1.607281952969826e-10, -1.6070503256850398e-10, 
    -1.6062567023870001e-10, -1.6048309516101578e-10, 
    -1.6027388196712654e-10, -1.5999816016069145e-10, 
    -1.5965927316115844e-10, -1.5926319207696187e-10, 
    -1.5881774988071803e-10, -1.5833177409124013e-10, 
    -1.5781420820497881e-10, -1.5727330347080687e-10, 
    -1.5671594473939846e-10, -1.5614717947927264e-10, 
    -1.5556995875559979e-10, -1.5498511760242713e-10, -1.543915683974813e-10, 
    -1.5378669088498555e-10, -1.5316686224234764e-10, 
    -1.5252808912786521e-10, -1.5186667230725723e-10, 
    -1.5117987055675036e-10, -1.504664862725002e-10, -1.4972735550928703e-10, 
    -1.4896568617406722e-10, -1.4818723894766247e-10, 
    -1.4740032569245859e-10, -1.4661563089228904e-10, 
    -1.4584585897447172e-10, -1.4510525159590121e-10, 
    -1.4440897221709482e-10, -1.4377242733859097e-10, 
    -1.4321053980757167e-10, -1.4273704653562297e-10, 
    -1.4236384087474319e-10, -1.4210039648075626e-10, 
    -1.4195332560122306e-10, -1.4192607638934697e-10, 
    -1.4201878277574319e-10, -1.4222828542700826e-10, 
    -1.4254829136554232e-10, -1.4296968153225153e-10, 
    -1.4348092094383049e-10, -1.4406854591923892e-10, 
    -1.4471769692915128e-10, -1.4541266605012742e-10, 
    -1.4613740523694521e-10, -1.4687599891855883e-10, 
    -1.4761305460081614e-10, -1.4833400951888694e-10, 
    -1.4902535436077743e-10, -1.4967477901612318e-10, 
    -1.5027124865787107e-10, -1.5080503280552088e-10, 
    -1.5126770279379699e-10, -1.5165214111352971e-10, -1.519525429867564e-10, 
    -1.5216445856698335e-10, -1.5228486803357341e-10, 
    -1.5231229155416893e-10, -1.52246926866995e-10, -1.5209080972758536e-10, 
    -1.5184794893236868e-10, -1.5152444957599682e-10, 
    -1.5112855825253277e-10, -1.5067062178863244e-10, 
    -1.5016292955882767e-10, -1.4961944348253539e-10, 
    -1.4905539008451456e-10, -1.4848673360933739e-10, 
    -1.4792957079060974e-10, -1.4739947825432694e-10, 
    -1.4691085896526544e-10, -1.4647633641393309e-10, 
    -1.4610625386741408e-10, -1.4580831598823056e-10, 
    -1.4558738739525216e-10, -1.4544546357537489e-10, 
    -1.4538180280713349e-10, -1.4539318171724818e-10, 
    -1.4547424807591201e-10, -1.4561792872806357e-10, 
    -1.4581584454245786e-10, -1.4605870421504714e-10, 
    -1.4633665850988569e-10, -1.4663960813713859e-10, 
    -1.4695745921191857e-10, -1.4728035787242739e-10, 
    -1.4759889869770075e-10, -1.4790434067103099e-10, 
    -1.4818882867267602e-10, -1.4844562616290222e-10, 
    -1.4866934654785011e-10, -1.4885615961238869e-10, 
    -1.4900395890532935e-10, -1.4911244954142236e-10, 
    -1.4918313653168967e-10, -1.4921920061735475e-10, -1.492252419061419e-10, 
    -1.4920691295336236e-10, -1.491704426506856e-10, -1.4912210068027493e-10, 
    -1.4906763188149372e-10, -1.4901171200653823e-10, 
    -1.4895747059229745e-10, -1.4890613507086059e-10, 
    -1.4885682367126846e-10, -1.4880652019049448e-10, 
    -1.4875023919255231e-10, -1.486813837496368e-10, -1.4859226474345354e-10, 
    -1.484747563026244e-10, -1.4832102605405147e-10, -1.4812429721766857e-10, 
    -1.4787956469065532e-10, -1.4758421644092395e-10, 
    -1.4723849964266148e-10, -1.4684579908264033e-10, 
    -1.4641269413925023e-10, -1.4594878679114721e-10, -1.454663171689625e-10, 
    -1.4497959455705557e-10, -1.4450427056892804e-10, 
    -1.4405652594228553e-10, -1.4365220992205688e-10, 
    -1.4330600346600044e-10, -1.4303064214916899e-10, 
    -1.4283626992273603e-10, -1.4272993473597478e-10, 
    -1.4271526680202341e-10, -1.4279233718784791e-10, 
    -1.4295771191140491e-10, -1.4320466515709652e-10, 
    -1.4352353781023918e-10, -1.4390220800028682e-10, 
    -1.4432663399804097e-10, -1.4478143068702373e-10, 
    -1.4525044740833481e-10, -1.4571732219088375e-10, 
    -1.4616598830971127e-10, -1.4658113083679032e-10, 
    -1.4694858957119957e-10, -1.4725572102034985e-10, 
    -1.4749172625870187e-10, -1.476479543828592e-10, -1.4771819861819603e-10, 
    -1.4769895968444508e-10, -1.4758968620718586e-10, 
    -1.4739295247234396e-10, -1.4711455107243542e-10, 
    -1.4676345665560358e-10, -1.4635163929260851e-10, -1.458936954808611e-10, 
    -1.4540629310415255e-10, -1.4490744258954812e-10, 
    -1.4441562215854506e-10, -1.4394881690300368e-10, -1.435235343705249e-10, 
    -1.4315388003274186e-10, -1.4285077121433732e-10, 
    -1.4262135834368927e-10, -1.4246870000467e-10, -1.4239173076536356e-10, 
    -1.4238550505722688e-10, -1.4244169843658348e-10, 
    -1.4254930569566884e-10, -1.4269546354812385e-10, 
    -1.4286632277302365e-10, -1.4304788938316875e-10, -1.432267867260978e-10, 
    -1.4339087894029535e-10, -1.435297510158034e-10, -1.4363504594457239e-10, 
    -1.4370068297976953e-10, -1.4372297370065576e-10,
  // Sqw-F(9, 0-1999)
    0.017430167320618094, 0.017429969627323169, 0.017429310972700725, 
    0.017428000725615837, 0.017425740808424614, 0.017422152898051255, 
    0.017416812272557536, 0.017409284695805473, 0.017399162504062812, 
    0.017386096280343096, 0.017369819134626024, 0.017350161559430588, 
    0.017327055971704645, 0.017300531236022598, 0.01727069854468934, 
    0.017237730882629802, 0.017201838840593467, 0.017163245716969547, 
    0.017122164672705855, 0.017078780225669457, 0.017033235673958095, 
    0.016985627224972977, 0.016936004784813032, 0.016884378626150588, 
    0.016830730575702967, 0.016775027989941169, 0.016717238635475307, 
    0.016657344647934346, 0.016595353979291717, 0.016531308115160483, 
    0.01646528530202692, 0.016397399021705183, 0.016327791942520067, 
    0.016256626025585565, 0.016184069837611628, 0.016110284392242533, 
    0.016035408989327374, 0.015959548532404791, 0.01588276367512936, 
    0.015805064885241301, 0.015726411141179768, 0.015646713525984072, 
    0.015565843500798935, 0.015483645177024217, 0.015399950512010206, 
    0.015314596070358351, 0.015227439849384114, 0.0151383766732433, 
    0.01504735080713507, 0.014954364706471436, 0.014859483160893042, 
    0.01476283248041332, 0.01466459476397932, 0.014564997659483256, 
    0.014464300347892816, 0.014362776750216456, 0.014260697157633449, 
    0.014158309617482771, 0.014055822465068793, 0.0139533893651917, 
    0.01385109810843759, 0.013748964188075426, 0.013646929863086934, 
    0.013544869001948951, 0.013442597525241375, 0.013339888762642409, 
    0.0132364925625514, 0.013132156596762938, 0.013026648041135461, 
    0.012919773726358153, 0.012811396960732538, 0.012701449524413809, 
    0.012589937791391063, 0.01247694249963196, 0.012362612295339899, 
    0.0122471517542305, 0.012130805067575036, 0.012013836925188605, 
    0.011896512304362866, 0.011779076878784222, 0.011661739611543305, 
    0.011544658824014804, 0.011427932678956339, 0.011311594624306781, 
    0.011195613951728448, 0.011079901260056063, 0.010964318297461841, 
    0.010848691397160524, 0.01073282752315277, 0.010616531804847531, 
    0.01049962536200205, 0.010381962205208085, 0.010263444044685986, 
    0.010144031954480647, 0.010023754021723248, 0.009902708358814731, 
    0.009781061161455256, 0.0096590398413633552, 0.0095369216261681732, 
    0.0094150183716415238, 0.0092936586417119178, 0.0091731683489686099, 
    0.0090538513867334178, 0.0089359717056956521, 0.0088197381870257375, 
    0.0087052934457074443, 0.008592707380695631, 0.0084819759010532313, 
    0.0083730248354022558, 0.0082657186150574043, 0.0081598729471449166, 
    0.0080552703956121297, 0.0079516775895437531, 0.0078488626933390961, 
    0.0077466118046693091, 0.00764474308589183, 0.0075431176661414209, 
    0.0074416466514842343, 0.0073402939219856054, 0.0072390747480978518, 
    0.0071380505953694247, 0.0070373207790482692, 0.0069370118553504449, 
    0.0068372657760393434, 0.0067382278766133178, 0.0066400357134010352, 
    0.0065428096181517946, 0.0064466456166066225, 0.0063516110845913687, 
    0.0062577432217508959, 0.0061650501418005028, 0.0060735141399271041, 
    0.0059830965275626301, 0.0058937433376774137, 0.005805391204172403, 
    0.005717972799540171, 0.0056314213584566907, 0.0055456739972993881, 
    0.0054606737338758213, 0.0053763702922920353, 0.0052927199240447734, 
    0.0052096845743310827, 0.0051272307664237083, 0.005045328568414058, 
    0.0049639509532232711, 0.0048830737758470636, 0.0048026764842664799, 
    0.004722743565097668, 0.0046432666133390966, 0.0045642468171758965, 
    0.0044856975715985457, 0.0044076468848828904, 0.0043301392246016925, 
    0.0042532364680392797, 0.0041770176767862814, 0.0041015775051909641, 
    0.0040270231719370872, 0.0039534700640235345, 0.0038810361897566471, 
    0.0038098358361400215, 0.0037399728992909731, 0.0036715344284979287, 
    0.0036045849432423901, 0.0035391620418473184, 0.0034752737216402416, 
    0.0034128976826222797, 0.0033519827054301326, 0.0032924520005172654, 
    0.0032342082415834955, 0.0031771398437773126, 0.0031211279433174359, 
    0.003066053490684683, 0.00301180388742336, 0.0029582786720360492, 
    0.0029053938818202375, 0.0028530848682502379, 0.0028013075046377347, 
    0.0027500378773795222, 0.002699270679599249, 0.0026490166161667193, 
    0.0025992991751493575, 0.0025501511218789827, 0.0025016110328434449, 
    0.002453720117151299, 0.0024065194862653177, 0.0023600479423847871, 
    0.0023143402759601369, 0.002269426004416849, 0.0022253284540586027, 
    0.0021820640868741225, 0.0021396419997137262, 0.0020980635664832044, 
    0.00205732224297388, 0.0020174035961576403, 0.0019782856441559245, 
    0.0019399395922385357, 0.0019023310218766142, 0.0018654215375276133, 
    0.0018291708080714103, 0.0017935388688473343, 0.001758488489590112, 
    0.0017239873755691844, 0.0016900099627241789, 0.0016565385962070943, 
    0.0016235639432148846, 0.0015910845774680783, 0.0015591057720003364, 
    0.0015276376346314228, 0.0014966928022304659, 0.0014662839636517397, 
    0.001436421499295488, 0.0014071115052603782, 0.0013783544153097953, 
    0.0013501443526992088, 0.0013224692482640358, 0.0012953116647359904, 
    0.0012686501833364535, 0.0012424611482240193, 0.0012167205343784967, 
    0.0011914057072506957, 0.0011664968754059616, 0.0011419780936838615, 
    0.001117837744450537, 0.0010940684974948941, 0.0010706668146967485, 
    0.0010476321155026345, 0.0010249657482989867, 0.0010026699193506372, 
    0.0009807467168452082, 0.00095919733725823735, 0.00093802158094049898, 
    0.00091721764031251363, 0.00089678216360645666, 0.00087671054467226904, 
    0.00085699736807502138, 0.00083763692969324947, 0.0008186237555934463, 
    0.00079995305398049472, 0.00078162105344772566, 0.0007636252021344861, 
    0.00074596422342182759, 0.00072863804168382283, 0.00071164760442236062, 
    0.00069499463391154857, 0.00067868134233879435, 0.00066271014032795884, 
    0.00064708336128821106, 0.00063180301520387658, 0.00061687057717449304, 
    0.00060228680976352647, 0.00058805161490642452, 0.00057416391089255424, 
    0.00056062153216586278, 0.000547421153243272, 0.00053455824154064271, 
    0.0005220270460445822, 0.00050982062870732483, 0.00049793094293127207, 
    0.0004863489589777343, 0.0004750648305757194, 0.00046406809171978811, 
    0.00045334786891922482, 0.00044289309293759271, 0.00043269269571124321, 
    0.00042273578234167434, 0.0004130117738926466, 0.00040351052285321579, 
    0.00039422240812941244, 0.0003851384191150436, 0.00037625023810936085, 
    0.00036755032711914765, 0.00035903201962195035, 0.00035068961142441631, 
    0.00034251843884068091, 0.00033451492848203263, 0.00032667660205067692, 
    0.00031900202210675347, 0.00031149067056124964, 0.00030414275971274419, 
    0.00029695898461230076, 0.00028994023384861851, 0.00028308728207525959, 
    0.00027640049073672881, 0.00026987954305869995, 0.00026352323564217606, 
    0.00025732934268546772, 0.00025129456105229013, 0.00024541453633711714, 
    0.00023968396285699986, 0.00023409674492953488, 0.00022864620327864895, 
    0.0002233253089406893, 0.00021812692729634701, 0.00021304405632801703, 
    0.00020807004536940117, 0.00020319878305799142, 0.00019842484568368912, 
    0.00019374359960380833, 0.00018915125395378948, 0.00018464486265899524, 
    0.00018022227781937236, 0.00017588205983736839, 0.00017162335295990773, 
    0.00016744573783448151, 0.00016334907478448104, 0.00015933335236602682, 
    0.00015539855508026415, 0.00015154456180355193, 0.0001477710827385111, 
    0.00014407763790986487, 0.00014046357504339085, 0.00013692811978298662, 
    0.00013347044730000244, 0.00013008976197891801, 0.00012678537134316395, 
    0.00012355674176400686, 0.00012040352654104838, 0.00011732556118883, 
    0.00011432282557847315, 0.00011139537727537803, 0.00010854326433026158, 
    0.00010576642840718474, 0.00010306461015706147, 0.00010043726810398155, 
    9.7883520179850147e-05, 9.5402113806255156e-05, 9.299142660468172e-05, 
    9.0649496000609216e-05, 8.8374072718657665e-05, 8.6162690876734598e-05, 
    8.4012746326028249e-05, 8.1921575093615338e-05, 7.9886525097927475e-05, 
    7.7905016392478107e-05, 7.5974587612246446e-05, 7.4092928595214226e-05, 
    7.225790093426111e-05, 7.046754922402924e-05, 6.8720105918697755e-05, 
    6.7013992112784616e-05, 6.5347815452284591e-05, 6.3720365130226787e-05, 
    6.2130602883053433e-05, 6.0577648383211778e-05, 5.9060757583661169e-05, 
    5.7579293409420504e-05, 5.6132689535033845e-05, 5.4720409532953208e-05, 
    5.3341905058710373e-05, 5.1996577610780842e-05, 5.0683748518427608e-05, 
    4.9402641081554113e-05, 4.8152377300198628e-05, 4.6931989640523835e-05, 
    4.5740446147914706e-05, 4.457668533150698e-05, 4.3439655950956951e-05, 
    4.2328356361320172e-05, 4.124186847412422e-05, 4.0179382562117716e-05, 
    3.9140210815677355e-05, 3.8123789412561735e-05, 3.7129670536835376e-05, 
    3.6157506988472545e-05, 3.5207032586546488e-05, 3.4278041457760164e-05, 
    3.3370368626994131e-05, 3.2483873305975435e-05, 3.1618425177884878e-05, 
    3.0773893061711847e-05, 2.9950134804713236e-05, 2.9146987189470779e-05, 
    2.8364255029529943e-05, 2.7601699339532307e-05, 2.6859025303942682e-05, 
    2.6135871514175747e-05, 2.5431802401034696e-05, 2.4746305831303052e-05, 
    2.4078797426505449e-05, 2.3428632360390776e-05, 2.2795124340302507e-05, 
    2.2177570371212528e-05, 2.1575278942443131e-05, 2.0987598643168885e-05, 
    2.0413944016223335e-05, 1.9853815735731158e-05, 1.9306812891463368e-05, 
    1.8772636162962562e-05, 1.8251081802854552e-05, 1.7742027444351659e-05, 
    1.7245411641851904e-05, 1.6761209632439782e-05, 1.628940801459912e-05, 
    1.582998088991864e-05, 1.538286956781723e-05, 1.4947967296656964e-05, 
    1.4525109773520696e-05, 1.4114071511183347e-05, 1.3714567587590383e-05, 
    1.3326259920126701e-05, 1.2948767002218754e-05, 1.2581675991729597e-05, 
    1.2224556103405487e-05, 1.1876972381549537e-05, 1.1538499067202617e-05, 
    1.1208731898264205e-05, 1.0887298779284937e-05, 1.0573868339049851e-05, 
    1.0268155976142174e-05, 9.9699270984545745e-06, 9.6789974062470271e-06, 
    9.3952302541451307e-06, 9.1185313416000806e-06, 8.8488411993348668e-06, 
    8.5861261262527732e-06, 8.3303683551471521e-06, 8.0815562600957189e-06, 
    7.8396753553742269e-06, 7.6047006819921234e-06, 7.3765909606407932e-06, 
    7.1552846452730055e-06, 6.9406977835064279e-06, 6.7327234150042994e-06, 
    6.5312321441418111e-06, 6.3360735155352426e-06, 6.1470778912933363e-06, 
    5.9640586493358753e-06, 5.7868146577514744e-06, 5.6151330916862395e-06, 
    5.448792717008727e-06, 5.2875677505759427e-06, 5.1312323222603545e-06, 
    4.9795654257909788e-06, 4.8323560869890582e-06, 4.6894083361343387e-06, 
    4.5505454837061398e-06, 4.4156131908788207e-06, 4.2844809098801946e-06, 
    4.1570414357163364e-06, 4.033208536306195e-06, 3.9129128745199776e-06, 
    3.7960966624819121e-06, 3.6827076558011939e-06, 3.5726931768196064e-06, 
    3.4659948377890905e-06, 3.3625445240147644e-06, 3.2622620128598963e-06, 
    3.1650543807372216e-06, 3.0708171219731117e-06, 2.9794367063954964e-06, 
    2.8907941612496691e-06, 2.8047691928396518e-06, 2.7212443634183436e-06, 
    2.6401088996164313e-06, 2.5612618096376555e-06, 2.4846141064262363e-06, 
    2.410090050596842e-06, 2.3376274255775656e-06, 2.2671769283420978e-06, 
    2.1987008026090052e-06, 2.1321708614390478e-06, 2.0675660526343942e-06, 
    2.004869721096263e-06, 1.9440667251248048e-06, 1.885140570035433e-06, 
    1.8280707315577578e-06, 1.7728303464954278e-06, 1.7193844430095852e-06, 
    1.6676888597751159e-06, 1.6176899598355216e-06, 1.5693251809249492e-06, 
    1.5225243864264705e-06, 1.4772118988131044e-06, 1.433309023816797e-06, 
    1.3907368196526822e-06, 1.3494188417916313e-06, 1.309283603584688e-06, 
    1.2702665363199878e-06, 1.2323113011026416e-06, 1.195370389322517e-06, 
    1.1594050338264357e-06, 1.124384527629713e-06, 1.0902850996528769e-06, 
    1.0570885230760273e-06, 1.0247806298349657e-06, 9.9334988003637263e-07, 
    9.6278609439312776e-07, 9.3307941192373715e-07, 9.0421949206290547e-07, 
    8.7619494816119181e-07, 8.4899298040276882e-07, 8.2259917177059185e-07, 
    7.9699741627512276e-07, 7.721699604274165e-07, 7.4809754998584035e-07, 
    7.247596808155213e-07, 7.0213495150484684e-07, 6.8020150715502474e-07, 
    6.5893754960114129e-07, 6.3832187423799808e-07, 6.1833438107893507e-07, 
    5.989565025361424e-07, 5.8017149407570146e-07, 5.6196454774286697e-07, 
    5.4432270954759179e-07, 5.2723460752003723e-07, 5.1069002225054499e-07, 
    4.9467935259982338e-07, 4.7919304162579055e-07, 4.6422103068641156e-07, 
    4.4975230230153568e-07, 4.3577455742874595e-07, 4.2227405242313416e-07, 
    4.092355997288439e-07, 3.9664271674475508e-07, 3.8447789296555714e-07, 
    3.7272293686054802e-07, 3.6135936215305072e-07, 3.5036877620652404e-07, 
    3.3973324032083055e-07, 3.294355799545241e-07, 3.1945963137454279e-07, 
    3.0979041779979217e-07, 3.0041425328477592e-07, 2.9131877544637529e-07, 
    2.824929105621376e-07, 2.7392677613790885e-07, 2.6561152860314224e-07, 
    2.57539166593536e-07, 2.4970230411679723e-07, 2.4209393110635572e-07, 
    2.3470718163446707e-07, 2.2753513039307115e-07, 2.2057063650949813e-07, 
    2.1380624903717305e-07, 2.0723418219784248e-07, 2.0084636048665905e-07, 
    1.9463452628372205e-07, 1.8859039607024977e-07, 1.8270584755560072e-07, 
    1.7697311855865159e-07, 1.7138500028120885e-07, 1.6593501092334161e-07, 
    1.6061754051580965e-07, 1.5542796203094204e-07, 1.503627074617241e-07, 
    1.4541930889801781e-07, 1.4059640471524177e-07, 1.358937092258785e-07, 
    1.313119424492459e-07, 1.2685271512473246e-07, 1.2251836457870327e-07, 
    1.1831173920581136e-07, 1.142359341561727e-07, 1.1029398684623599e-07, 
    1.0648854810215699e-07, 1.0282155080298152e-07, 9.9293902592899721e-08, 
    9.5905230375672186e-08, 9.2653702434883068e-08, 8.9535948045210607e-08, 
    8.6547085995215662e-08, 8.368086265925364e-08, 8.0929889433118709e-08, 
    7.8285959142911836e-08, 7.5740413633626018e-08, 7.3284530114936839e-08, 
    7.0909893439369622e-08, 6.8608724202168163e-08, 6.6374138847561542e-08, 
    6.4200325800230135e-08, 6.2082631000387093e-08, 6.0017554920402159e-08, 
    5.8002671172864626e-08, 5.6036482552172997e-08, 5.4118234256544413e-08, 
    5.2247705197472835e-08, 5.0424997762727181e-08, 4.8650343611624739e-08, 
    4.6923939560374731e-08, 4.524582276765701e-08, 4.3615789887995613e-08, 
    4.2033359956890317e-08, 4.049777695073722e-08, 3.9008044475609015e-08, 
    3.7562983160658143e-08, 3.6161300119686349e-08, 3.4801660400692781e-08, 
    3.3482751475337836e-08, 3.2203334341602493e-08, 3.0962277366397312e-08, 
    2.9758572113041524e-08, 2.859133276793631e-08, 2.7459782857136934e-08, 
    2.6363233751942647e-08, 2.5301059699876082e-08, 2.4272673109094062e-08, 
    2.3277502726255418e-08, 2.2314975600146944e-08, 2.1384502662183788e-08, 
    2.0485466623171659e-08, 1.9617210958860249e-08, 1.8779028829631312e-08, 
    1.7970151876838455e-08, 1.7189739609659388e-08, 1.6436871261744869e-08, 
    1.5710542324161855e-08, 1.500966825809711e-08, 1.4333097149638736e-08, 
    1.3679632312703978e-08, 1.3048064277556053e-08, 1.2437210416986326e-08, 
    1.1845958920038976e-08, 1.1273313136222421e-08, 1.0718431596237897e-08, 
    1.0180659363000842e-08, 9.6595468302295798e-09, 9.1548534782385353e-09, 
    8.666535403994202e-09, 8.1947173615689398e-09, 7.7396515019123373e-09, 
    7.3016666318308548e-09, 6.8811125621795256e-09, 6.4783047736204498e-09, 
    6.0934741980329605e-09, 5.7267262998259854e-09, 5.3780122130440253e-09, 
    5.047113327837891e-09, 4.7336389490301236e-09, 4.4370355337439249e-09, 
    4.1566048045769196e-09, 3.8915278808934359e-09, 3.6408923787930083e-09, 
    3.4037202230491929e-09, 3.178994429771429e-09, 2.9656841545215761e-09, 
    2.762767713468264e-09, 2.5692538565743926e-09, 2.3842013268011598e-09, 
    2.2067366606200655e-09, 2.0360694997791786e-09, 1.8715044330643386e-09, 
    1.712447931758554e-09, 1.5584091783359577e-09, 1.408993820317075e-09, 
    1.2638905862956555e-09, 1.1228514258510265e-09, 9.8566694979279914e-10, 
    8.5213951111327241e-10, 7.220569156862068e-10, 5.9516963111725324e-10, 
    4.7117423619358407e-10, 3.4970500367219051e-10, 2.3033488243474763e-10, 
    1.1258598202494553e-10, -4.0510603349386289e-12, -1.2009045264395615e-10, 
    -2.3601942644774004e-10, -3.5226397951171562e-10, 
    -4.6915501142625517e-10, -5.8689799684480402e-10, 
    -7.0554901121673744e-10, -8.2499983639954538e-10, 
    -9.4497409821581356e-10, -1.0650358236888976e-09, 
    -1.1846105961343934e-09, -1.3030185774898191e-09, 
    -1.4195172914466926e-09, -1.5333512110739798e-09, 
    -1.6438041443723368e-09, -1.7502501622124051e-09, 
    -1.8521985398064501e-09, -1.9493288092747386e-09, 
    -2.0415126690354326e-09, -2.1288208372650366e-09, 
    -2.2115140993492566e-09, -2.2900194188766683e-09, -2.364893049513733e-09, 
    -2.4367738915434192e-09, -2.5063308642660311e-09, 
    -2.5742086880538203e-09, -2.6409762926967465e-09, 
    -2.7070819941778243e-09, -2.7728187442561219e-09, 
    -2.8383021593060398e-09, -2.9034628515794872e-09, -2.968053624330144e-09, 
    -3.0316708289952091e-09, -3.0937882197115529e-09, 
    -3.1538005046741757e-09, -3.2110731450197688e-09, 
    -3.2649942928851781e-09, -3.315024696184322e-09, -3.3607413957581357e-09, 
    -3.4018717461089322e-09, -3.4383149706576689e-09, 
    -3.4701497614475485e-09, -3.4976274745379544e-09, 
    -3.5211520049643267e-09, -3.5412483270535096e-09, 
    -3.5585228510359593e-09, -3.5736191430749536e-09, -3.587172948214174e-09, 
    -3.5997701371366188e-09, -3.6119108629819136e-09, 
    -3.6239822615876825e-09, -3.6362413014386493e-09, 
    -3.6488082045145067e-09, -3.6616701277673946e-09, 
    -3.6746937988580472e-09, -3.6876453953692646e-09, 
    -3.7002153857671069e-09, -3.7120461090023532e-09, 
    -3.7227597330036048e-09, -3.7319847091876415e-09, 
    -3.7393789993450265e-09, -3.7446490271893891e-09, 
    -3.7475636201559784e-09, -3.7479628655467641e-09, 
    -3.7457620124286909e-09, -3.7409510747424275e-09, 
    -3.7335907910708053e-09, -3.7238058692032863e-09, 
    -3.7117762124015217e-09, -3.6977269354358397e-09, 
    -3.6819176256308387e-09, -3.6646313782210016e-09, -3.646163813844544e-09, 
    -3.6268124512593963e-09, -3.6068666253405152e-09, 
    -3.5865983776577147e-09, -3.566254634929005e-09, -3.5460512102877261e-09, 
    -3.5261689629353413e-09, -3.5067525086565023e-09, 
    -3.4879115406279385e-09, -3.4697247054808232e-09, 
    -3.4522455516051847e-09, -3.4355099614793473e-09, -3.419544136128084e-09, 
    -3.4043722718894537e-09, -3.3900229219497834e-09, 
    -3.3765333868073171e-09, -3.3639515115326913e-09, 
    -3.3523347822888145e-09, -3.341746718386436e-09, -3.3322510585804395e-09, 
    -3.3239042850344074e-09, -3.3167473800194831e-09, 
    -3.3107975984791183e-09, -3.3060412394081151e-09, 
    -3.3024281172707925e-09, -3.299868479048157e-09, -3.2982327259857339e-09, 
    -3.297354222532443e-09, -3.2970350477975101e-09, -3.297054420494011e-09, 
    -3.2971791239679083e-09, -3.2971752191277573e-09, 
    -3.2968200226085379e-09, -3.2959134824851817e-09, -3.294287950654079e-09, 
    -3.2918156975907527e-09, -3.2884135611014964e-09, 
    -3.2840445824408225e-09, -3.2787165900358595e-09, 
    -3.2724781219277735e-09, -3.265412119903768e-09, -3.2576280934244566e-09, 
    -3.2492533576788942e-09, -3.2404240744092312e-09, 
    -3.2312765458297327e-09, -3.2219393017897417e-09, 
    -3.2125262137581112e-09, -3.2031309212371022e-09, 
    -3.1938226299369696e-09, -3.1846434274149878e-09, -3.175607070834597e-09, 
    -3.1666993408149567e-09, -3.15787983157634e-09, -3.1490851903413102e-09, 
    -3.1402335743978058e-09, -3.1312302042014003e-09, 
    -3.1219736258767445e-09, -3.1123624318345407e-09, 
    -3.1023019542427174e-09, -3.0917106107744506e-09, 
    -3.0805254258315338e-09, -3.0687064866627114e-09, 
    -3.0562399481018721e-09, -3.0431395005553953e-09, 
    -3.0294461290981854e-09, -3.0152262349571459e-09, 
    -3.0005681528610841e-09, -2.9855773213948362e-09, -2.970370300023255e-09, 
    -2.9550680676746006e-09, -2.9397888990624043e-09, -2.924641351612517e-09, 
    -2.9097177327345596e-09, -2.8950885498691178e-09, 
    -2.8807982756206684e-09, -2.8668627975339767e-09, 
    -2.8532687086692826e-09, -2.8399745912490055e-09, 
    -2.8269141823187069e-09, -2.8140013200592374e-09, 
    -2.8011362924461723e-09, -2.7882132559226368e-09, 
    -2.7751281629536554e-09, -2.7617867237711835e-09, 
    -2.7481117758665351e-09, -2.7340495977143221e-09, 
    -2.7195746066347919e-09, -2.7046921348311371e-09, 
    -2.6894389447672768e-09, -2.6738814646970568e-09, 
    -2.6581117472197878e-09, -2.6422414721198343e-09, 
    -2.6263943631893347e-09, -2.6106976583606749e-09, 
    -2.5952732331693686e-09, -2.5802291718571252e-09, 
    -2.5656523922484475e-09, -2.5516030187737816e-09, 
    -2.5381108632562603e-09, -2.5251743552877492e-09, 
    -2.5127619065795279e-09, -2.5008155901768897e-09, 
    -2.4892567331536503e-09, -2.4779929479213904e-09, -2.466925942155394e-09, 
    -2.4559595105954178e-09, -2.4450069892522755e-09, -2.433997681803492e-09, 
    -2.422881703960793e-09, -2.4116329930178859e-09, -2.4002502441058955e-09, 
    -2.3887558206193336e-09, -2.377192739961426e-09, -2.3656200998884493e-09, 
    -2.3541072955846793e-09, -2.3427276065803991e-09, 
    -2.3315516470202142e-09, -2.3206412950234026e-09, -2.310044525431073e-09, 
    -2.2997916208110404e-09, -2.2898929458448629e-09, -2.280338485819153e-09, 
    -2.2710990014814873e-09, -2.2621287004488931e-09, 
    -2.2533690394936806e-09, -2.2447533566433141e-09, 
    -2.2362118438618391e-09, -2.2276765452103579e-09, 
    -2.2190859695827524e-09, -2.2103890884564993e-09, -2.201548463635201e-09, 
    -2.1925424462708464e-09, -2.1833662980012286e-09, 
    -2.1740323039456351e-09, -2.1645688354171298e-09, 
    -2.1550184914128298e-09, -2.1454353578305757e-09, 
    -2.1358815747334646e-09, -2.1264233252518873e-09, 
    -2.1171265308077755e-09, -2.1080524173487885e-09, 
    -2.0992533098276385e-09, -2.0907688512321685e-09, 
    -2.0826229851628449e-09, -2.0748218579904967e-09, 
    -2.0673528732302041e-09, -2.0601849151871917e-09, 
    -2.0532698317538456e-09, -2.0465449920708739e-09, 
    -2.0399368419272194e-09, -2.0333651410305163e-09, 
    -2.0267476605581804e-09, -2.0200049518064338e-09, 
    -2.0130649252971489e-09, -2.0058668638909094e-09, 
    -1.9983646706889823e-09, -1.9905290735873065e-09, 
    -1.9823487182450221e-09, -1.9738300432008632e-09, 
    -1.9649960507305259e-09, -1.955884030236874e-09, -1.9465425024738769e-09, 
    -1.9370275933567586e-09, -1.9273991834527109e-09, 
    -1.9177170664068546e-09, -1.9080374587470813e-09, 
    -1.8984100320138578e-09, -1.8888756780146548e-09, 
    -1.8794650549621556e-09, -1.8701979915105385e-09, 
    -1.8610836137026024e-09, -1.8521211505545582e-09, 
    -1.8433012201219139e-09, -1.834607478118682e-09, -1.8260184112021205e-09, 
    -1.8175091893130304e-09, -1.8090534175825086e-09, 
    -1.8006247690371099e-09, -1.7921984130696547e-09, 
    -1.7837522699250444e-09, -1.7752680646687733e-09, 
    -1.7667322377057699e-09, -1.7581366744590366e-09, 
    -1.7494792837456446e-09, -1.7407643787018188e-09, 
    -1.7320028545796022e-09, -1.7232120659261773e-09, 
    -1.7144154164996618e-09, -1.7056415538747063e-09, 
    -1.6969232169903867e-09, -1.6882956783631351e-09, 
    -1.6797948849860721e-09, -1.6714553314533022e-09, 
    -1.6633078279935127e-09, -1.6553772818785369e-09, -1.647680689942877e-09, 
    -1.6402254956941482e-09, -1.6330085217251368e-09, 
    -1.6260155506431376e-09, -1.6192217114704547e-09, 
    -1.6125926435056509e-09, -1.606086448649117e-09, -1.5996562632033757e-09, 
    -1.5932533358108365e-09, -1.58683031046412e-09, -1.580344511088081e-09, 
    -1.573760907204124e-09, -1.5670545570565226e-09, -1.5602122729568594e-09, 
    -1.5532334081519084e-09, -1.5461296644744605e-09, 
    -1.5389239900000241e-09, -1.5316486186512758e-09, 
    -1.5243424693450338e-09, -1.5170480896656948e-09, 
    -1.5098084387188377e-09, -1.502663718322721e-09, -1.4956485370822201e-09, 
    -1.4887895728724537e-09, -1.4821039198164502e-09, 
    -1.4755981898710584e-09, -1.4692684204465382e-09, 
    -1.4631007454176182e-09, -1.4570727881579534e-09, 
    -1.4511555936326615e-09, -1.4453160225700706e-09, 
    -1.4395193523914286e-09, -1.4337319468903662e-09, 
    -1.4279237813867775e-09, -1.422070663812861e-09, -1.4161559728154747e-09, 
    -1.4101718338098285e-09, -1.4041196067849287e-09, 
    -1.3980097101774916e-09, -1.3918607512945584e-09, -1.385698079918344e-09, 
    -1.3795518496040446e-09, -1.3734547723557423e-09, 
    -1.3674397160510166e-09, -1.3615373671243805e-09, 
    -1.3557740991732223e-09, -1.3501702505276492e-09, 
    -1.3447388831139148e-09, -1.3394851352453443e-09, 
    -1.3344061425572896e-09, -1.3294915449381528e-09, 
    -1.3247244572141917e-09, -1.3200828159142257e-09, 
    -1.3155409657117706e-09, -1.3110713645885571e-09, -1.306646249904846e-09, 
    -1.3022392004960131e-09, -1.2978264550458991e-09, 
    -1.2933879800089599e-09, -1.288908201022068e-09, -1.2843764278691365e-09, 
    -1.2797869311250431e-09, -1.2751387221417136e-09, 
    -1.2704350364046823e-09, -1.2656825798477529e-09, 
    -1.2608905697669016e-09, -1.2560696585204046e-09, 
    -1.2512307881133566e-09, -1.2463840871208136e-09, 
    -1.2415378728618175e-09, -1.2366978760501377e-09, 
    -1.2318667269116804e-09, -1.2270437825534975e-09, 
    -1.2222252935371264e-09, -1.21740492172956e-09, -1.2125745320092085e-09, 
    -1.2077252075056849e-09, -1.2028483612536846e-09, 
    -1.1979368465692977e-09, -1.1929859385582312e-09, 
    -1.1879941007283942e-09, -1.1829634373974284e-09, 
    -1.1778998161142261e-09, -1.1728126107785315e-09, 
    -1.1677141548790471e-09, -1.1626188853056856e-09, 
    -1.1575423332627485e-09, -1.1525000110077868e-09, 
    -1.1475063216027921e-09, -1.1425735783994257e-09, -1.137711235400069e-09, 
    -1.1329253533931512e-09, -1.128218383441796e-09, -1.1235892209544187e-09, 
    -1.1190335648146804e-09, -1.1145444820568442e-09, -1.110113159514245e-09, 
    -1.1057297404652954e-09, -1.1013841911564467e-09, 
    -1.0970671062234891e-09, -1.0927704110048417e-09, 
    -1.0884879001179795e-09, -1.0842155903024394e-09, 
    -1.0799518625705583e-09, -1.0756974190408909e-09, 
    -1.0714550361479938e-09, -1.0672291743566638e-09, -1.063025454663472e-09, 
    -1.058850062405321e-09, -1.0547091040580115e-09, -1.0506079959884172e-09, 
    -1.0465508942383367e-09, -1.042540251167289e-09, -1.0385765023178135e-09, 
    -1.0346579400595497e-09, -1.0307807640704449e-09, 
    -1.0269393308290038e-09, -1.0231265500554293e-09, 
    -1.0193344275894746e-09, -1.0155546633738426e-09, 
    -1.0117792774955284e-09, -1.0080011813257349e-09, 
    -1.0042146520270847e-09, -1.0004156645831677e-09, 
    -9.9660207080135042e-10, -9.9277361214762332e-10, 
    -9.8893182101618875e-10, -9.8507981606944959e-10, 
    -9.8122207810880167e-10, -9.7736423181334291e-10, 
    -9.7351289415287653e-10, -9.696755954469526e-10, -9.6586078616559912e-10, 
    -9.6207788763749148e-10, -9.5833736229487266e-10, 
    -9.5465071301331419e-10, -9.5103037076444989e-10, 
    -9.4748939472576967e-10, -9.4404097233888271e-10, 
    -9.4069767871599139e-10, -9.3747056511019122e-10, 
    -9.3436809454205466e-10, -9.3139505918593167e-10, 
    -9.2855155494337242e-10, -9.2583217824662007e-10, 
    -9.2322551377800236e-10, -9.2071405896295758e-10, 
    -9.1827460369763237e-10, -9.1587912003511853e-10, 
    -9.1349611628148812e-10, -9.1109238464936691e-10, 
    -9.0863502097051842e-10, -9.060935752224931e-10, -9.034421386688944e-10, 
    -9.0066121326910265e-10, -8.9773917828427191e-10, 
    -8.9467323543769777e-10, -8.9146972214048929e-10, 
    -8.8814377281321525e-10, -8.8471832191197854e-10, 
    -8.8122255254889943e-10, -8.7768988267048662e-10, -8.741556852263643e-10, 
    -8.7065489846392591e-10, -8.6721974891844052e-10, -8.638777252920472e-10, 
    -8.6065001162218169e-10, -8.5755042223094448e-10, 
    -8.5458495270112891e-10, -8.5175190946385349e-10, 
    -8.4904260877878771e-10, -8.4644252021462285e-10, 
    -8.4393275222609187e-10, -8.4149172523439216e-10, 
    -8.3909688426743428e-10, -8.3672629067203274e-10, -8.343600079985557e-10, 
    -8.3198113505620759e-10, -8.2957648587720374e-10, -8.271368563456978e-10, 
    -8.2465693802444727e-10, -8.2213490347327984e-10, 
    -8.1957177203204292e-10, -8.1697062871063712e-10, 
    -8.1433581249692404e-10, -8.116721449395244e-10, -8.0898428737225049e-10, 
    -8.0627625925995254e-10, -8.0355115801520957e-10, 
    -8.0081104847404148e-10, -7.9805703153642702e-10, 
    -7.9528941544218566e-10, -7.9250796971563044e-10, 
    -7.8971218306677765e-10, -7.8690152803855607e-10, 
    -7.8407565388106857e-10, -7.8123453121833935e-10, 
    -7.7837852946111015e-10, -7.7550845778256815e-10, 
    -7.7262557638606869e-10, -7.697316206067142e-10, -7.6682884484032152e-10, 
    -7.6392012588987183e-10, -7.6100909697469161e-10, 
    -7.5810034417083548e-10, -7.5519960166424243e-10, 
    -7.5231394273482913e-10, -7.4945190620523673e-10, -7.466235261309314e-10, 
    -7.4384022474078802e-10, -7.4111453913840557e-10, 
    -7.3845967625733102e-10, -7.3588890269700056e-10, 
    -7.3341479338706575e-10, -7.3104840769160818e-10, 
    -7.2879842515812552e-10, -7.2667035420959332e-10, 
    -7.2466584656445387e-10, -7.2278222690114399e-10, 
    -7.2101226312913814e-10, -7.1934423725359895e-10, 
    -7.1776230078739593e-10, -7.1624713738109734e-10, -7.147768486713152e-10, 
    -7.1332802840932855e-10, -7.1187692454763806e-10, 
    -7.1040061608542061e-10, -7.0887808640401903e-10, 
    -7.0729113921803066e-10, -7.0562505676987407e-10, 
    -7.0386899861645384e-10, -7.0201607745733358e-10, 
    -7.0006317541625904e-10, -6.9801050391215175e-10, 
    -6.9586099925160423e-10, -6.9361961095991451e-10, 
    -6.9129259281862296e-10, -6.8888684596389857e-10, 
    -6.8640940785549029e-10, -6.8386709431500535e-10, 
    -6.8126635727238401e-10, -6.7861328707589707e-10, 
    -6.7591377674420168e-10, -6.7317374124607043e-10, 
    -6.7039937955798726e-10, -6.6759735379683908e-10, 
    -6.6477488796700227e-10, -6.6193970531551038e-10, 
    -6.5909982589296885e-10, -6.5626321100498401e-10, 
    -6.5343733292965439e-10, -6.5062867360887427e-10, 
    -6.4784227041947548e-10, -6.450813417124207e-10, -6.4234706244419535e-10, 
    -6.396385259804938e-10, -6.3695291456105352e-10, -6.3428584551166786e-10, 
    -6.3163190933576409e-10, -6.2898529261804652e-10, 
    -6.2634047976576747e-10, -6.2369291681651789e-10, 
    -6.2103963818355874e-10, -6.1837974567853552e-10, 
    -6.1571475678671873e-10, -6.1304876419611501e-10, 
    -6.1038843379580624e-10, -6.0774282216484422e-10, 
    -6.0512305458855885e-10, -6.0254186216789716e-10, 
    -6.0001303608192242e-10, -5.9755077339963383e-10, 
    -5.9516900543187838e-10, -5.928806595036338e-10, -5.9069695028866277e-10, 
    -5.8862666589883492e-10, -5.866755459034084e-10, -5.8484572512487169e-10, 
    -5.8313533680173784e-10, -5.8153827265737095e-10, 
    -5.8004417874239368e-10, -5.7863867182677611e-10, 
    -5.7730383024015334e-10, -5.7601892516381496e-10, 
    -5.7476140172689754e-10, -5.7350802297581502e-10, 
    -5.7223616160402732e-10, -5.709250883124295e-10, -5.695572345018758e-10, 
    -5.6811924967301733e-10, -5.6660281810847858e-10, 
    -5.6500510916426182e-10, -5.6332884637980114e-10, 
    -5.6158192807772154e-10, -5.5977667255178514e-10, 
    -5.5792868484055307e-10, -5.5605550343032209e-10, 
    -5.5417508325401784e-10, -5.5230432085630146e-10, 
    -5.5045768628420483e-10, -5.4864615734815358e-10, 
    -5.4687648866193853e-10, -5.4515091643499548e-10, 
    -5.4346727067024907e-10, -5.4181950528217598e-10, 
    -5.4019850905112337e-10, -5.3859315729081828e-10, 
    -5.3699142840730383e-10, -5.3538150029353655e-10, 
    -5.3375269253831066e-10, -5.3209620403825086e-10, -5.304055684175568e-10, 
    -5.2867685059635711e-10, -5.2690857556493691e-10, 
    -5.2510149626956023e-10, -5.2325819780637322e-10, 
    -5.2138268954981243e-10, -5.1947997267033436e-10, 
    -5.1755570240664507e-10, -5.1561589614045535e-10, 
    -5.1366675961496158e-10, -5.1171453770244127e-10, 
    -5.0976542097584281e-10, -5.0782541267216294e-10, 
    -5.0590018529696578e-10, -5.0399484117298521e-10, 
    -5.0211366016888785e-10, -5.0025978230880041e-10, 
    -4.9843492485146589e-10, -4.9663914029208104e-10, 
    -4.9487071063596543e-10, -4.9312615780153838e-10, 
    -4.9140046381267113e-10, -4.8968741085842388e-10, 
    -4.8798010658341586e-10, -4.8627154755393531e-10, 
    -4.8455524066757159e-10, -4.8282573774662769e-10, 
    -4.8107909311278801e-10, -4.7931311985916e-10, -4.7752750410770596e-10, 
    -4.7572370129744564e-10, -4.7390471588682592e-10, 
    -4.7207474683397331e-10, -4.7023882211561971e-10, 
    -4.6840241713398687e-10, -4.6657116924890482e-10, 
    -4.6475066239908611e-10, -4.6294635256322335e-10, 
    -4.6116356803087403e-10, -4.5940761990492336e-10, 
    -4.5768391363114532e-10, -4.559981027805138e-10, -4.5435615160362169e-10, 
    -4.5276437546945012e-10, -4.5122934465450597e-10, 
    -4.4975774925902915e-10, -4.4835614161174991e-10, -4.470306669440963e-10, 
    -4.4578673711334048e-10, -4.4462874014760342e-10, 
    -4.4355974513668241e-10, -4.4258129319481678e-10, 
    -4.4169320341064324e-10, -4.4089347177784798e-10, 
    -4.4017818463168708e-10, -4.3954151207246713e-10, 
    -4.3897569611820743e-10, -4.3847110619636853e-10, 
    -4.3801629219318272e-10, -4.3759810879707738e-10, 
    -4.3720185463286503e-10, -4.3681153105669765e-10, 
    -4.3641014316264442e-10, -4.3598014174950455e-10, 
    -4.3550394218387135e-10, -4.349645819915888e-10, -4.3434642389428824e-10, 
    -4.3363594808047989e-10, -4.3282250588262245e-10, 
    -4.3189904807739923e-10, -4.3086270183466011e-10, 
    -4.2971519470796506e-10, -4.2846301597128419e-10, 
    -4.2711732973839231e-10, -4.2569357934199429e-10, 
    -4.2421083960019517e-10, -4.2269089278368827e-10, 
    -4.2115715326982619e-10, -4.1963343634107595e-10, 
    -4.1814273790270126e-10, -4.1670603460943485e-10, 
    -4.1534125893884707e-10, -4.1406244983743696e-10, 
    -4.1287920693486587e-10, -4.1179639879642119e-10, 
    -4.1081419398629174e-10, -4.0992833939734086e-10, 
    -4.0913069908054132e-10, -4.0840993070507359e-10, 
    -4.0775230140635663e-10, -4.0714250687345784e-10, 
    -4.0656448567840082e-10, -4.0600212286684115e-10, 
    -4.0543987108835156e-10, -4.0486319898436632e-10, 
    -4.0425893694072574e-10, -4.0361546645606293e-10, 
    -4.0292287216315806e-10, -4.0217298347021303e-10, 
    -4.0135943437640582e-10, -4.0047768806759343e-10, 
    -3.9952511091987307e-10, -3.9850102099664222e-10, 
    -3.9740677748891898e-10, -3.9624580507212785e-10, 
    -3.9502360748743558e-10, -3.937476638798544e-10, -3.9242725411175529e-10, 
    -3.9107313671954567e-10, -3.896971577932663e-10, -3.8831172546371932e-10, 
    -3.8692926703449012e-10, -3.8556163739933322e-10, 
    -3.8421959785030056e-10, -3.8291234045418291e-10, 
    -3.8164717120212952e-10, -3.8042930293361153e-10, 
    -3.7926183078222358e-10, -3.7814581376642442e-10, -3.77080524843216e-10, 
    -3.7606372738842104e-10, -3.7509203884713903e-10, 
    -3.7416125328414326e-10, -3.7326668466544056e-10, 
    -3.7240340967694742e-10, -3.7156648965191466e-10, 
    -3.7075110346200111e-10, -3.6995268276756703e-10, 
    -3.6916697147611143e-10, -3.6839012774625147e-10, 
    -3.6761879146616379e-10, -3.6685019708420415e-10, 
    -3.6608225698653701e-10, -3.6531368200458604e-10, 
    -3.6454403250470566e-10, -3.6377376240456495e-10, 
    -3.6300415828807156e-10, -3.6223724115384193e-10, 
    -3.6147553776623899e-10, -3.6072182128513966e-10, 
    -3.5997874102667089e-10, -3.5924846820186282e-10, 
    -3.5853229756334927e-10, -3.5783032781145512e-10, 
    -3.5714117522693636e-10, -3.5646184604234836e-10, -3.557876961430071e-10, 
    -3.5511257903661696e-10, -3.5442911113081147e-10, -3.537291192606704e-10, 
    -3.5300416851985375e-10, -3.5224620985742009e-10, 
    -3.5144823614426258e-10, -3.5060496603586665e-10, -3.4971342118109e-10, 
    -3.4877343487956925e-10, -3.4778795015283999e-10, 
    -3.4676315130719892e-10, -3.4570832780936574e-10, 
    -3.4463553804264313e-10, -3.4355899659159928e-10, 
    -3.4249430131713918e-10, -3.4145745918816073e-10, 
    -3.4046386071054201e-10, -3.3952719432358637e-10, 
    -3.3865846539160734e-10, -3.3786512074363772e-10, -3.371504460167659e-10, 
    -3.3651320418769816e-10, -3.3594764891376693e-10, 
    -3.3544384852175708e-10, -3.3498839942943806e-10, 
    -3.3456539210401842e-10, -3.3415764351875182e-10, -3.337480394280877e-10, 
    -3.3332091818806822e-10, -3.3286332136665248e-10, 
    -3.3236606929871377e-10, -3.3182446316710066e-10, 
    -3.3123861407499672e-10, -3.3061329219416795e-10, 
    -3.2995736381429606e-10, -3.2928278318379941e-10, 
    -3.2860330003380847e-10, -3.2793293583145162e-10, 
    -3.2728444679084875e-10, -3.2666784839844992e-10, 
    -3.2608923219078045e-10, -3.2554991233967927e-10, 
    -3.2504607205659491e-10, -3.2456887356474315e-10, 
    -3.2410508981170136e-10, -3.236381238734968e-10, -3.231494121807457e-10, 
    -3.2261997321177718e-10, -3.2203204884129611e-10, 
    -3.2137061974245263e-10, -3.206247291566828e-10, -3.1978843835468158e-10, 
    -3.1886142140601818e-10, -3.1784908977562656e-10, 
    -3.1676231065871055e-10, -3.1561670691080484e-10, 
    -3.1443167162572962e-10, -3.1322909310696213e-10, -3.120319755987332e-10, 
    -3.1086297387158938e-10, -3.0974302576762406e-10, 
    -3.0869008305793829e-10, -3.0771809060562641e-10, 
    -3.0683621010480923e-10, -3.0604840148341019e-10, 
    -3.0535329719835969e-10, -3.0474445082952939e-10, 
    -3.0421085496422445e-10, -3.0373776730676276e-10, 
    -3.0330769341109779e-10, -3.0290153270406392e-10, 
    -3.0249973758029609e-10, -3.0208345298080078e-10, 
    -3.0163551327374182e-10, -3.0114129101994964e-10, 
    -3.0058927844982961e-10, -2.9997145660465312e-10, 
    -2.9928337408341121e-10, -2.9852401932898368e-10, 
    -2.9769546644734664e-10, -2.9680239642776509e-10, 
    -2.9585148693482923e-10, -2.9485081209328369e-10, 
    -2.9380921345317666e-10, -2.9273577817723445e-10, 
    -2.9163937417458293e-10, -2.9052835183144903e-10, 
    -2.8941032898592802e-10, -2.8829212088959085e-10, 
    -2.8717973111206112e-10, -2.860784376255495e-10, -2.8499286572438192e-10, 
    -2.8392708541225354e-10, -2.8288464689339333e-10, 
    -2.8186858594360099e-10, -2.8088135711813493e-10, 
    -2.7992474543412284e-10, -2.7899973047404589e-10, 
    -2.7810639128955899e-10, -2.7724381264584238e-10, 
    -2.7641008606145248e-10, -2.7560236455118343e-10, 
    -2.7481703160808139e-10, -2.7404992176071794e-10, -2.732966346175659e-10, 
    -2.72552854572461e-10, -2.7181470043949741e-10, -2.7107901234551891e-10, 
    -2.703436192349903e-10, -2.6960748048874091e-10, -2.6887075384858229e-10, 
    -2.6813473029895761e-10, -2.6740169495536469e-10, 
    -2.6667465861965362e-10, -2.6595704108969845e-10, 
    -2.6525228332822738e-10, -2.6456345759905168e-10, 
    -2.6389285995582801e-10, -2.6324168225424476e-10, -2.626097198517126e-10, 
    -2.6199519485678022e-10, -2.6139467539465563e-10, 
    -2.6080313993826322e-10, -2.60214126757383e-10, -2.5962002635833209e-10, 
    -2.590124331156408e-10, -2.5838258874314486e-10, -2.5772183237758834e-10, 
    -2.5702209472008604e-10, -2.5627634084724605e-10, 
    -2.5547899852810838e-10, -2.5462630735149644e-10, 
    -2.5371661714843191e-10, -2.5275057681334328e-10, 
    -2.5173126237443735e-10, -2.5066417317989973e-10, 
    -2.4955714551895261e-10, -2.4842012933778657e-10, 
    -2.4726486698881944e-10, -2.461044310297513e-10, -2.4495269078117035e-10, 
    -2.4382366173524383e-10, -2.427308294172578e-10, -2.4168644900248457e-10, 
    -2.407009147377642e-10, -2.3978220013799394e-10, -2.3893547158718215e-10, 
    -2.381628658303154e-10, -2.3746348725274475e-10, -2.3683359088628237e-10, 
    -2.3626696175941493e-10, -2.3575539845169874e-10, 
    -2.3528930245454561e-10, -2.348582527975341e-10, -2.3445154158980654e-10, 
    -2.3405859558381809e-10, -2.3366930163536152e-10, 
    -2.3327415350657712e-10, -2.3286431155526838e-10, -2.324315471789967e-10, 
    -2.3196817086528062e-10, -2.3146693265706336e-10, 
    -2.3092099620899214e-10, -2.303239706255126e-10, -2.2967004643669786e-10, 
    -2.2895420618273201e-10, -2.2817251819823685e-10, 
    -2.2732244829135205e-10, -2.264031894921107e-10, -2.2541592933453883e-10, 
    -2.2436407999414484e-10, -2.2325338516961355e-10, 
    -2.2209195063939532e-10, -2.2089014724107022e-10, -2.196604423009089e-10, 
    -2.1841711936060254e-10, -2.1717594202724269e-10, 
    -2.1595374162432984e-10, -2.1476795936774402e-10, 
    -2.1363613290937824e-10, -2.1257536104851431e-10, 
    -2.1160172291997895e-10, -2.1072971381120847e-10, 
    -2.0997166886854068e-10, -2.0933724753836346e-10, 
    -2.0883296934400378e-10, -2.0846187991443641e-10, 
    -2.0822332693024856e-10, -2.0811291787664388e-10, 
    -2.0812264550040885e-10, -2.0824119777041693e-10, 
    -2.0845443724609283e-10, -2.0874605693007741e-10, 
    -2.0909833031863668e-10, -2.0949296229901241e-10, 
    -2.0991195156210156e-10, -2.1033845244353795e-10, 
    -2.1075753185913543e-10, -2.1115681289246842e-10, -2.115269290347377e-10, 
    -2.118617785669244e-10, -2.1215854154565812e-10, -2.1241746516100704e-10, 
    -2.1264143061816899e-10, -2.1283534062186046e-10, 
    -2.1300537101863844e-10, -2.1315816057017323e-10, -2.132999995595515e-10, 
    -2.1343610751337855e-10, -2.1357004234969017e-10, 
    -2.1370331176765166e-10, -2.1383520067437146e-10, 
    -2.1396284239619036e-10, -2.1408148970583642e-10, 
    -2.1418497195980805e-10, -2.1426626696914179e-10, 
    -2.1431812869089268e-10, -2.1433370379865622e-10, 
    -2.1430709136314205e-10, -2.1423377370042575e-10, 
    -2.1411092373117092e-10, -2.1393754839974425e-10, -2.137145084669305e-10, 
    -2.134444034834872e-10, -2.1313138214446823e-10, -2.1278087897394325e-10, 
    -2.1239934046377294e-10, -2.1199392559107537e-10, 
    -2.1157222719397641e-10, -2.1114199966300059e-10, 
    -2.1071091108337717e-10, -2.1028629887982035e-10, 
    -2.0987495360919402e-10, -2.0948290272846187e-10, -2.091152414676482e-10, 
    -2.0877598425176597e-10, -2.0846797193922807e-10, -2.081928431350901e-10, 
    -2.0795108415810872e-10, -2.0774215345130715e-10, -2.075646696606071e-10, 
    -2.0741665623257439e-10, -2.0729580954320152e-10, 
    -2.0719974668474778e-10, -2.0712623247809753e-10, 
    -2.0707330746767985e-10, -2.0703933813253246e-10, 
    -2.0702295599103388e-10, -2.0702290405679902e-10, 
    -2.0703780558041217e-10, -2.0706590253384279e-10, 
    -2.0710479290468176e-10, -2.0715121549915236e-10, 
    -2.0720091706145957e-10, -2.0724866288781786e-10, 
    -2.0728834668836267e-10, -2.0731325481538027e-10, 
    -2.0731642703104872e-10, -2.0729109771425422e-10, 
    -2.0723116362965352e-10, -2.0713163780245274e-10, 
    -2.0698902816929051e-10, -2.0680162575429517e-10, 
    -2.0656964863988182e-10, -2.0629524747624552e-10, 
    -2.0598236247390708e-10, -2.0563646383917657e-10, 
    -2.0526418194958708e-10, -2.0487286919591414e-10, 
    -2.0447012909748438e-10, -2.0406335766520157e-10, 
    -2.0365930503237441e-10, -2.0326371035932099e-10, 
    -2.0288101340714229e-10, -2.0251417464136852e-10, 
    -2.0216459467301269e-10, -2.0183214779177984e-10, 
    -2.0151531556375185e-10, -2.012114193567358e-10, -2.0091691012306452e-10, 
    -2.0062772158028478e-10, -2.0033961909086036e-10, 
    -2.0004854369684966e-10, -1.9975090563471836e-10, 
    -1.9944379985017325e-10, -1.9912513995555825e-10, -1.987936995128027e-10, 
    -1.9844906542220461e-10, -1.9809152599784429e-10, -1.977219084685833e-10, 
    -1.9734141566774986e-10, -1.9695145371061304e-10, 
    -1.9655351057726304e-10, -1.9614906681735312e-10, -1.957395466810074e-10, 
    -1.9532631653654089e-10, -1.949107095690613e-10, -1.9449405160095371e-10, 
    -1.940776972187596e-10, -1.93663043138388e-10, -1.9325152798587269e-10, 
    -1.9284462214590173e-10, -1.9244380773616385e-10, 
    -1.9205056716861063e-10, -1.9166638289734775e-10, -1.912927579264785e-10, 
    -1.9093126193894505e-10, -1.9058358088756919e-10, 
    -1.9025158621114611e-10, -1.8993737763418585e-10, 
    -1.8964330011691241e-10, -1.89371912875712e-10, -1.8912590344784462e-10, 
    -1.8890793222864884e-10, -1.887204175701143e-10, -1.8856527271236392e-10, 
    -1.8844361193159973e-10, -1.8835545247023594e-10, 
    -1.8829943881313298e-10, -1.8827262220026944e-10, 
    -1.8827032109278465e-10, -1.8828608179009587e-10, -1.883117633145585e-10, 
    -1.8833773950227163e-10, -1.8835323099924208e-10, 
    -1.8834673701535146e-10, -1.8830656649919168e-10, 
    -1.8822141623796209e-10, -1.8808097084673102e-10, 
    -1.8787647559696207e-10, -1.8760125086903413e-10, 
    -1.8725108776809863e-10, -1.8682450416131467e-10, 
    -1.8632282980939065e-10, -1.8575012253018344e-10, 
    -1.8511290067189944e-10, -1.8441973483967084e-10, 
    -1.8368072721928123e-10, -1.8290693194277009e-10, 
    -1.8210976287866975e-10, -1.8130045363524331e-10, 
    -1.8048960148994103e-10, -1.7968683785437418e-10, 
    -1.7890063563409746e-10, -1.7813824736177061e-10, 
    -1.7740576290398395e-10, -1.7670825923046931e-10, 
    -1.7604998737087263e-10, -1.7543459204471648e-10, 
    -1.7486529215386186e-10, -1.7434503081735093e-10, 
    -1.7387655990564235e-10, -1.7346245617609009e-10, 
    -1.7310507610642696e-10, -1.7280646873717951e-10, 
    -1.7256823257287719e-10, -1.7239136624844433e-10, 
    -1.7227610449926414e-10, -1.7222175823043773e-10, 
    -1.7222657296020725e-10, -1.7228761786191175e-10, 
    -1.7240069451283988e-10, -1.7256030300427443e-10, 
    -1.7275962641657696e-10, -1.7299058775141449e-10, 
    -1.7324393613170485e-10, -1.7350939609864099e-10, 
    -1.7377586708957892e-10, -1.7403166629567254e-10, 
    -1.7426482507050191e-10, -1.7446341960726888e-10, 
    -1.7461593195920926e-10, -1.7471163919759595e-10, 
    -1.7474100056837921e-10, -1.7469604915821185e-10, 
    -1.7457075347189554e-10, -1.743613567581394e-10, -1.7406664830628226e-10, 
    -1.7368816656129652e-10, -1.7323030353626376e-10, 
    -1.7270030949278171e-10, -1.7210815160064406e-10, 
    -1.7146624738651006e-10, -1.7078904383102774e-10, 
    -1.7009246323729086e-10, -1.6939322714198426e-10, 
    -1.6870808386922681e-10, -1.6805298725112408e-10, 
    -1.6744227803856412e-10, -1.6688791804514489e-10, 
    -1.6639885719712068e-10, -1.6598056774563617e-10, 
    -1.6563482037923219e-10, -1.6535972253427564e-10, 
    -1.6515003077694464e-10, -1.6499772951232e-10, -1.6489284974417246e-10, 
    -1.6482443483242547e-10, -1.6478159296587997e-10, 
    -1.6475452376167084e-10, -1.6473542477152455e-10, 
    -1.6471916859364052e-10, -1.6470369325923033e-10, -1.646900467920102e-10, 
    -1.6468207247720311e-10, -1.6468577200022563e-10, 
    -1.6470842254603412e-10, -1.6475751084211699e-10, 
    -1.6483963311639115e-10, -1.6495945340386675e-10, 
    -1.6511884684568155e-10, -1.6531630471670073e-10, 
    -1.6554665860543144e-10, -1.6580114598264688e-10, 
    -1.6606780043381208e-10, -1.663321096903201e-10, -1.6657789460358668e-10, 
    -1.6678830185804959e-10, -1.6694684378824718e-10, 
    -1.6703841417751131e-10, -1.6705020247492258e-10, 
    -1.6697247687845772e-10, -1.6679922271669905e-10, 
    -1.6652858531961829e-10, -1.6616314638999438e-10, 
    -1.6571002035752961e-10, -1.6518077414284198e-10, 
    -1.6459116397503077e-10, -1.6396069004153051e-10, 
    -1.6331196586712929e-10, -1.6266990295898719e-10, 
    -1.6206070936312238e-10, -1.615107507472577e-10, -1.6104527196548722e-10, 
    -1.6068706959892782e-10, -1.6045516231653841e-10, 
    -1.6036354559009292e-10, -1.6042012642899536e-10, 
    -1.6062591404312529e-10, -1.6097455737485538e-10, 
    -1.6145228017277186e-10, -1.6203825271229695e-10, 
    -1.6270541044211659e-10, -1.6342167807833138e-10, 
    -1.6415156034306072e-10, -1.6485798743099643e-10, -1.655042993802486e-10, 
    -1.6605625384850439e-10, -1.6648391794415531e-10, 
    -1.6676329270447252e-10, -1.668775832229335e-10, -1.6681800636725857e-10, 
    -1.6658408169173615e-10, -1.6618338770076788e-10, 
    -1.6563080683317386e-10, -1.6494730502307301e-10, 
    -1.6415835237054779e-10, -1.6329208808567255e-10, 
    -1.6237739155516019e-10, -1.6144198321816442e-10, 
    -1.6051070849733512e-10, -1.5960413441886378e-10, 
    -1.5873755000534191e-10, -1.5792043650812656e-10, 
    -1.5715643865709889e-10, -1.5644380031010218e-10, 
    -1.5577622821473663e-10, -1.5514406747948749e-10, -1.545356863739449e-10, 
    -1.5393893941092394e-10, -1.5334257168358534e-10, 
    -1.5273745858007594e-10, -1.5211757690289244e-10, 
    -1.5148064402462187e-10, -1.5082840249330235e-10, 
    -1.5016653170375837e-10, -1.4950423586833243e-10, 
    -1.4885354808631585e-10, -1.4822844342703959e-10, 
    -1.4764382757948811e-10, -1.4711449025607461e-10, 
    -1.4665411675267369e-10, -1.4627441972499855e-10, 
    -1.4598444985058134e-10, -1.4579012956364026e-10, 
    -1.4569402328778647e-10, -1.4569534961161548e-10, 
    -1.4579021872221962e-10, -1.4597205080180167e-10, 
    -1.4623213632211647e-10, -1.465602835201071e-10, -1.4694548213149004e-10, 
    -1.4737653722806892e-10, -1.4784261892858513e-10, -1.483336790098897e-10, 
    -1.488407252949343e-10, -1.4935592924918279e-10, -1.4987258664183519e-10, 
    -1.5038493781160423e-10, -1.5088789337181668e-10, 
    -1.5137671373729749e-10, -1.5184666925117074e-10, 
    -1.5229275083373555e-10, -1.5270946839547537e-10, 
    -1.5309076592948733e-10, -1.5343009192167942e-10, 
    -1.5372062700352068e-10, -1.5395564684556339e-10, 
    -1.5412902333264058e-10, -1.5423578619812039e-10, 
    -1.5427270592180085e-10, -1.542388152121718e-10, -1.5413582424256008e-10, 
    -1.5396833513167099e-10, -1.5374382287133644e-10, 
    -1.5347236116020917e-10, -1.5316609840605242e-10, 
    -1.5283851121262071e-10, -1.5250349763590136e-10, 
    -1.5217440428908296e-10, -1.5186308825362185e-10, 
    -1.5157909721570621e-10, -1.5132907625596723e-10, 
    -1.5111645223152802e-10, -1.5094143603248261e-10, 
    -1.5080134344756785e-10, -1.5069119989407672e-10, 
    -1.5060455475118151e-10, -1.5053441814192183e-10, -1.504742201812778e-10, 
    -1.5041868163865017e-10, -1.5036450493528418e-10, 
    -1.5031081022717989e-10, -1.502592701708308e-10, -1.5021393087746394e-10, 
    -1.5018073352770987e-10, -1.5016679512628843e-10, 
    -1.5017952160616813e-10, -1.5022563765294147e-10, 
    -1.5031025395336984e-10, -1.5043605237026633e-10, 
    -1.5060268386767889e-10, -1.5080643945316207e-10, 
    -1.5104022057994954e-10, -1.5129381543563466e-10, 
    -1.5155444889603439e-10, -1.5180754893751379e-10, 
    -1.5203765046507571e-10, -1.5222935553054692e-10, 
    -1.5236826867896876e-10, -1.5244182845456763e-10, 
    -1.5243999169003773e-10, -1.5235572284433339e-10, 
    -1.5218529188546538e-10, -1.5192837878527683e-10, 
    -1.5158800604981268e-10, -1.5117033445627598e-10, 
    -1.5068434284614184e-10, -1.5014143512952875e-10, 
    -1.4955498478031015e-10, -1.4893984278947527e-10, 
    -1.4831181722996519e-10, -1.4768714064038272e-10, 
    -1.4708192830549843e-10, -1.4651163945850584e-10, 
    -1.4599056098227738e-10, -1.4553132768304109e-10, 
    -1.4514449853474378e-10, -1.4483822042934021e-10, 
    -1.4461798530398805e-10, -1.4448651497769018e-10, 
    -1.4444376463456194e-10, -1.4448706924406858e-10, 
    -1.4461140545823876e-10, -1.4480976603489539e-10, 
    -1.4507361025116491e-10, -1.4539337636270431e-10, 
    -1.4575899683289724e-10, -1.4616039180380215e-10, 
    -1.4658790261103609e-10, -1.4703263263324541e-10, 
    -1.4748666747488759e-10, -1.4794317038852843e-10, 
    -1.4839634432073624e-10, -1.4884128419395363e-10, 
    -1.4927373279259684e-10, -1.4968979321960537e-10, 
    -1.5008562483713498e-10, -1.5045718157799735e-10, 
    -1.5080002814633169e-10, -1.5110927380269257e-10, -1.513796283845538e-10, 
    -1.5160560983967174e-10, -1.5178185821414594e-10, 
    -1.5190354750996962e-10, -1.5196683128425483e-10, 
    -1.5196927975420599e-10, -1.5191023914254047e-10, 
    -1.5179108393446794e-10, -1.5161530158044539e-10, 
    -1.5138841316694703e-10, -1.5111771868973794e-10, 
    -1.5081189906721852e-10, -1.504805164546424e-10, -1.5013346006237356e-10, 
    -1.4978040077469502e-10, -1.4943030501063533e-10, 
    -1.4909104773099943e-10, -1.4876916773656591e-10, 
    -1.4846974776289236e-10, -1.4819644143845083e-10, 
    -1.4795160010731248e-10, -1.4773648620805833e-10, 
    -1.4755151629936638e-10, -1.4739652775132693e-10, 
    -1.4727100880934263e-10, -1.4717430600234763e-10, 
    -1.4710577254088121e-10, -1.4706488062634696e-10, -1.4705128947117703e-10 ;
}
